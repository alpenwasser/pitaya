`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mgBHxdGDKdFcNwl/Xx2WnyYZ7ba1BCdJcMSppx8JqLmJP1U5rviV9jaAKYu+vvTpty8wG5ySKIoS
ICgIgO6V5w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
igue1BkOrge2VpVQVRwbQ8pn3AwvEDZEEPivjx8QGiAj++94vrpWbiOuxNNKjjH1ls8/BaEytlI0
k+G45Qzlo4hEXwfSuLSzM8KYt7g93jXYIYktHgYGGNu3aOJWIi2cXvloY+pGimCQfcOaVGolYyH9
IhhuNsGI+eWWVc+rY1A=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gJvVWM2JGbFdLbLvMMWLTJj+1rqH54UUcXYKG5qFjk61PpU04kVJXA5qgHfKSfV47FFpOkWyN22u
u0uLrOs9ox304vJgx35pHrBVznc5vkixPUO5OgE9z6hg6DGVrR1ICyExjIUlE4PCmmXZSgHX425i
IFwgn4PSSI/h8v98oFI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t4ibrC3fv3Lns4KeFtgfU0Z9gO48OpMqyF8QTHX9pG9GXU6ON1Mwz9CGaY4RsDGBSh9SjdAjzOC7
DWGPrFvZZ60z4PHWFb/ltHG7ZyROVyTH8Viqlhp5P+JsNdL/PrlcBpWHVcuz+rDL86fTqg3qN4tx
v4r87ULAdYZgOZG+e9iHARRDB6b25+mXnOkUNhUVJS6cxT0RCQqXSCPbsLnYNHJjZavqWKw0KTal
tP9yKHaYnkC7UVygGE9noBkxODvffFE19n77vp9PheiDeUSy8Z47PUo2+siqo8e0gysEQHnxLlP/
fH8A43Gz3W+EXUPxtIzzfvSgQsbha1hgau3BGA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PAyVdC2D1HyXQ7ft0zBM7tk6aL5JONGo7BfiBFDG10oJ83HwdH56LT+Trixib8Kndb3P0tw1q4K8
EJpmbkhE3fG14gch0JwE/KtiyuIO9lgG2qguhfV4iePQPuZVaJ7xyqUie4W+bbBSVvas5rv6vVX8
z7W2qVRHYdfXNCetjqoY2ts6GYdW4uxn6oqwhrmhGAO4YoqS4fAycbuHV8FOP/q3flmo4ToG/B7T
bOSzfUIlSb0ea76VkzzwVtr6QJrrOqHBg6DD0qfmrUabDnqTnXyiGucIKAJwDo/cvtbYCZaEzNGR
0IBvCzC3/BXNiP2lgewJeUpK3r7ywO0EsZL61g==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eerX1NtxairFs8LyX2Rot1/JrHi6nVsYzT7q6CXGQY9k756B2QT2DwzPTG0l3px0LzPKCIrJleOv
BChpaRPWErPQGpaeonA8qUW64CRaVg1a7oKeczCYx3KJLZJr4vazqJ6KmIQJaJlb/nMqRDfBAMzZ
Hy9mUn6Zc3hOYohG+Ni3vbI2Ay3ZDCW5kiSquc4jbfTDLmWzKaAZLHg1r0vcGwUCEY9ZA1VG+ifo
iL2HO0b7txc9Cx4idh2fyH9tk2Ei2/s7hsfT9jfH62NP5jbwp1vrB6URWjZ8p39Bf7iMK8yzZBCH
MPph8zrM+5nJCLcrUf5zi2zCdvTE8t/M2h/tFw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 600848)
`protect data_block
GV5zZB1TdIcG4F0QnFDZKt2A6TGTV265tEPI2dP+u8m+2fQ4MRH7nId7KKBltEvc6wFyZ+E8Cf4O
+Wc0G2WLK4xgv/EuEX+prCARTv2Z2qO/YOoB3uWEQhKKFu6sXee00U1lRJnBmCezxCUuiaDaxVvo
qykfP6931Ke3RuLg7ovbLSJA3qWaA7HO9imPauUgrFwuIVBfsn3ggf17Z2sPEsv4gEIy480Xpl+E
Jou6auiU5sv/W6XN/Cs8CCobDqMiTtc+MgDSkkHyeYxKMMP4+h+Hrd3um9bUsU8ZXtWUNVXYBeIw
93jUPUXm8+xm3MefpyTkeRvKZYRWHwA4odqdmbIJ+fHy+iTx5sfgG27vxDbpBCaqic1WOw8FbGnJ
RuXptwMq96C4HEtVpKp3jUwGT8rC259F2CFI/xTkKoezLIUu45b1nLxAWt/QdoHD00Rc96oOwoQS
yk8WETxXshBwPb15iBYDBTnBXeI8LXFMxVSVH6ExXzxS8/NmoslpJJajKtbKTD/H5Qhr0uFj2MEV
cK1952ofTqw/DdkdWpmoRH6aPzzLIkYVWJAikF2LTTRUzwzoOexcLYFa/E+AuuYmwuEXA1g/IByP
63JsMHuiJZRFof1sSuE2+1QxT5HqqHWAIZx/0lnTAsIObhaIYWWJnpiG2KWH2hccC0hI2IvTJeFZ
t6sDMfDTO7USXK5ZscDeuGgs59j8a2Pdx7XmGPvH9m9Ab396R/gYdFUsQcsRiNlqIlircWv9LrtY
/tjIhR1frvqqAxjCom0Jp+LCv9fUI6I3xuxxtWRRhnhvqI7+plWefTVgK4sSrWw41P9/jAM3DaO6
5rHHRv15WeiGZvvhJOiyQBNFvoAKH7eZzlhmqUX+2dHycQIxmdCsyMP3OS7y5nR2dSNSd9Ye02uI
pYFcmXGdtUR5hiyBz+eG4fGkjFrsfuurFNZcytZIa5+it+I8tpH2zfwD/MD+yAQknMHqQjC+crMX
SgVihNMOvgk82bHUQxFuwq15yJcr68wFQFUgy9QszWYQfhjBgTMQheNoDqRBcCFqdsvrqKMqHQ9s
2Zj6MDI6MIGwhaVIp1EKeqcaK0tkZPEW/flbgWTnHDlO8S6jOvnyhxEh2//rTN75MoPCpvFzLnPw
bZBwbCawtLyResZrEqOFUnYVhIig/eKwqQ+lcnbl6nX4lU4hdZpWrYkoMFcbUl4oQFuVw4qY107i
J30UOiNN0pIgiSAK3frHoFLYLpJTafp7QcF5rcOZA0LpQVvm0WjPqbz5g29BX4anNaNXg7TmEse1
nMYGMZAQ1ylLYel70Its3gpyvv70hxReZtc4V8nkpBPBgg8/6VqPUZsZrd3fOjk1LZC6AJaU2eN/
G/9yQkXPTI7Jl1H0iremEcX0FeAasOhDHKg9uEj46QsX+1lf6cfzmzZWLGckfHu8Nzf6SpLSj80L
su2UG+hdcpV1IY7jU2mwDDsucuG/h7o4TslB8CxFJ4Q3nqfijXZYnvJjEP++rtuSg5XuYrRsaD1Q
M0X/V9S6W6QeRJh6+uKECDeFTL30ff8zC+8aO6OTjito+Dzk0kbtRFdY0MO84jRWEO4dqdffJYg2
U/Gignxqe/yGnnj1mVTIwShz9jdsk8RzkufwUeFjmQ9yb/hHwG2a/T/fmgawSc3/GHh8yhhlTdGt
KdvB6gpH0dMhLJa9sCzWqoA2T7z/2tvZ0AS9IumjbUOmzOMGdPpamRK6xJf/p9TOl6+yYoKLkKal
rnSvNduLxlvmRXDBfvYmfjdQkWEjpE6zZgT9PjIwWfGzs6obrzw8j6T4d3npAh5Z3BrQAvCFDCgg
UEPqxCMCK4cnXt0hOJRNY7aMaiw8b96iDa4+V+Qw3nNO6o1/h9wUsVFqmaMXhr5TgvKIgkmx6aRW
4/adK6pxhA7dJp1TnBigO0n4zY47xBZNI9ieO5hfZ+6FpicxTQrtAttm7W+m4IfX73HKipEstIo2
K27fBIQh04WrGktfFkZRPXyBgxMQPkceU4sP5GYx3pIZ68KtfXiauCNgcq0ELHdNT+/W16FjDlVD
IT0UeGf65ZVWTL2BuTUSSqs3GrmX7WlZL6Vhq1kWSx/cgH7g8QvO6upRzE98JZ0mL1iwgLR1OUqE
D6ype/KY4TtgSUvAAbI0pefbJ6bpDd34912zSj/ZzdRiEtpLVMKrf2GiN2Av+P/cqwkpPefpehoO
9SWdpyFuOhF7T8T59Zf9/DHZjcx3VHdPDG0iAO/CjP+4uxI7r3Uf0Gw4dqARci6df6WmBxFLdgNC
m56c1ktaBk8o6UQ3SmJlfqVnHgjsAkjCiht2LYNf8Gl9zOm/na5VdLcjXqvRjDACNhnrGCHlNQGM
u9Wk/AOj6Zefvighu7TqdStTWVoSGSM4LPON1h1KJUM95IbeHHLZ2MxMPY8qX9qQgILt1e6f417V
Qbn/+4wc1HpQRInI/EQHLal5FwUEhMvQYlDVrHUJ3P1PhY/abEs4KCZeheRDuH3T8BMc7aMXmLsD
5iNtx6uIzMCgYWJ4UHnECu7G2RtCBRMq2Yl92Z5IXOTP+43Hh77C6gzVXk3a2IW//W4d34Q+MY0S
OVXAMmrwnoGd/RUBlMeFx5JMnlJE5WVLIXr5BOoM7gxyRsatVXJWC5wzf51+X/SIORWymULDx7zr
PMZfmuHJijozN2jYLd2QuivjrYtj1OdVAB0XON7WCwlKKlWuKEQQPda6MApc+xxlMSJpLrgMoAF8
LY5+ppT6y4/k4aviA/Swe7pALpuG9lB6VLkFQp2qPyDBMf52BI5qHs2mcytZ6JQhir96UgS4hi5s
sHfUOHoss3pW7gjLn6VBkFGZ5BBe2Llfu+pGaFVSUooZDhCpvA8uFr+L2U4CjsYZoikVPmzPxBaj
+9gcef+QSRCSyNrkAVcu+ChqWsAd5ymqy9JNpcsZ8eng4F6Tg/fG4rDNx7KnDh4eDGzaXeY+Zrlz
UPjiG7Dc3v9AyaaunHsO6nM6Q2YGhTvH4HIo49/gZEI1QBT/bnCB4tUuJTzGXKAZ70Kkg2wh3RRT
ijEYk+2j5Ig2VaueVYXNQL+FKXd5NjISmgVtdNWkVta8T9AkCSM3H5Sqfdge/qIYdQa0u/ILhL/D
9OXocikL/UwIgpF8GESMC9FzfRvW5hc+bmT581ax+RiYmdC/Uj3Ba/qDpaOd1uk2W+JmdKN3XzKw
8LgwNj4h7lnRhaXXB2z6JIxTHzucvbY3GrK25h3WutXdfXUX7Vcu469fVmN8SMuQD8gA4AMFUHoi
rfk2+Dsso6QVkErQKVXTRoP7cQOJ31MZ5rFlwdRI1WAtjiL2KmMLkDRn4F49hvW2yXhxA/FkYp9n
SyRLFYHdZ1WVeDmx2u9nw0Hem1m/DajnlwsGttZ8bg8+cP3WfFzU9haniBbi0CfxgAZ8hvGtFY7x
AaQxFtShzl+0f1w1fIYeNHJ/4fth6M34XEiAYxS6ZTeQLC+Jn7Jz9MhA/e+YSBv0WC/KyV6JKRN2
vhV6TZsaHy2XpjKqKDMZA1+J6BKJGYcrzQKMuvCmvVetSIeDFX4cX7LxuP7h6m3IThNkQg42DTCd
WCC9P1tRAfByEqbfVMIwjxQ4xeDSB+YAeyhqGwA1AS1aKS3qhVYnmXTlHFIj5Fb22XGpPDqvyLu9
MLCZUkaG1i6Wex3gtKFG33JHOkGdJ3o8IRXf6E7RmoL335eA1iImvT5ZwPnGyt/HpotQEW21P2W7
FeozhyyYgA1QiuSx5+REyfMF/TvM1mSNhPJNl2Dk1jCDTRGERGAcvrveJa8q+uobUdVRpTHcayV5
fCv/Y6ilfRvDN4N1MbM2C8nDHOzE//RF6ZbwZJqG5mUI4qLduzahGB/aGe9bY9KS4onyeXJ5LXNi
Grik9bsexibxLkh6LTGEiyWyBZ6d8NZ9VbSdro9kOTTGLcvndKA1T8xcvTpoJBeSNUsN/OismDTY
hKXGoVPckLvZz0gZJqs1YWDilkWw2JEv/goncx2+4XvW8ljsuQCyold9ZRRIZ+rmYxD61A3bOPfK
9ZWEXqWkw90HY8PCgppNFqBxXrd5JtmaAhC1qg2TKA6U5qZJtdpq0QHUPiaT1KSoj4aeBs4OEYCD
EgwJkpWseL1v1TuBE0zQ7xFsou/WOZTwh+04W5inI9mcHvBiyK7aH9QVaF/SW3RqBKrEXUzLSHZJ
dyHPck0Qoqq3Bj2l5zdqiwN/tYdi4gs6pNcdfBzS7z11hvRxdZWpzhCsyx9QlLoVXtojEOGVyBpT
pMoU3i6JQXe29fU7hTVbcI0GXOapq5y4CwahVJhF1aCBWs8GHVtSNzSkxDrdK75p/zO6pqyG1dbB
4lxa9WuxL8duLBPG1XZRO6Gr8E/3XZsDng51WMAV0Y5GJQyOl7WBow6wiAHLxCOuJZJeA98TX0DL
L1ha135Vv74jVnMTdM1jx6YwZHl+iM27mAfSKBA8j4T9ovUqxXGVSqzV/7aojKtrfYT4dwkWrEoL
qeMpm2E/ffLCb/wC6SEvTEYtjVuIpk8QtsXj5r5jn80X/Kqb+Bb25LmTy43zG6I9bXeJCGeGqfka
tdtKEcMmuoMfy0ob2gkfP3qw6luCT2vrbJjxsPXcllNHl0cYgb8xBPotQxj33cRsn+QryDSsGpSN
EBedalkcCsz1YMBMEBD4j/tsOdyUnnlq2jmFF4Eeo68+ORJbUWHQ0R+EN/z+IIjI8lqoJz71RKeJ
1FHoKfC3E6rMPrhq5v6exde3BM6rlo0cCLC/A3sFLSxISr7jSXS1U4bHmePnzKtltmrK8b8ZRPNV
MoEk5fnSi/42cjAOauxgYgAGRmrHcyaP1frdQfHhW2hoT0CdCt6wZkfaacioZYq9wg+Y/zlTjPSP
A9D248zPIP8+ewgrBgxEmQt6PllX4axPJbXhB+IdJGZdc/2RCx3dwbHrcKsqJbkp0DSdBoxJjngk
7L/BUsPfOAlm4gJZ2nnV8ZA4+D9mWzvhUXDsbrUQ+CBgMKSZy5KvBQYP1f2C18Ipq3oB+paQOBzn
Mv5YwnLfzv0TKXo+IlnmrwT3H9VUCfSn+P3+JTew7YrnReB7AqO9EfIEU+B2WBAVSnFmpw4RWn4o
t/4+od6mcXHU9+Sq3XekraN/Q0E6J0Pm2JzlstUlFkWKMTrHW/zNBwW0Ak2aIKXgeSWrEZtqDl4Y
fXsyOd3cBC4GrjnplSdCxmRMvq0H8JhYiVy27cXoBG0lnZidEj9MLBUqRX6x2dTNSiENiUZSI+F4
ovs8lx+F54S9krFCUYKmLRBElA8/O8BJuw3R6xVobYfhtobsOzSFNRAUDvSbnW9bWONvufyS8YYU
ck8sG7UGiPavWw0T4RGySP8OpwZfllIM3ISger4ckumNMYZ0O+N/Ti5ntt7FYT0iCfRF818XJyQh
Fuyw53u4EAEuW+v4K1MvwYdDVrL/c6MhGvVuei0xtPALIvuhX3mhynScSPEI+00df3lFmRAmyKOW
B0YxOr2og0Kqw1cvth1WZYO+uftlLKvaprxwTmQhyEpn8Rz64/UmdD8z8Z9PcCoGFGIzeCUMDxbW
ThES/KRW56vQ4+zGcR88jZdsznlHOQ/OYN6vWi8S56oCbtcmfXiGahLdUAfF3ptak0ySR+65y+GD
QcP0eUVKXMZHS6169hWTNotuc1jkpiY48i6nkFZbxHQ9Qkjao27swbnrUlz6sGC7Wqzm2+ScY1FN
c9ppayvD75/lqrmSF9Kao2KsEUijCDOfZug9uqo7wpdsi2BF0jfH3cjFjMZmFRO5qmQFjJmlD21A
LRoJuZV0uu1HXnneegQgNQ9K75bZBALdFHSgAKuz4eOfkPuk6JbWAVFYLS5fOfK0hBsrWPA5/jT0
xUq8J+SISW3xX3P6YTadn7xnzvgbTDaOxQj+6rsGo0ATVbM6oEvCZoxuUqVtGJPIOg38oCicqPYS
klppPiXcRfzSw5PqpQiXeEwd4pcRFQ2ZHkg0TItIQB7L3D6Gpy+xvr7APU/Yp6qRfDFwwLYoMn6R
wNERRmJUIg3e5RRG9JbTKQ98DucECSIRZhQnolJoL8gpwcHWtwZp1PvOHn19QW+1iZD84ZN6DGHU
I31rPvjRU00hJ4yjYlxFKdEC8Dyd6VzgoE8ts/mC1kTyFJ06OBs9xAZYC13GEmeDpcJlbfNtyDtI
EjVZagAJatLbWiFvuddKvqc4mSmIIpGZGA9W8pqi2e7EmYOZBbrLdNoNxlk64g5JnvzMRsGzj1TG
Dula0qDsU1UuRmuvSThPyZ0BS3HtvXW6HL63F8w9EiVq8rLy7V/AL4VkC2FyuORhBvumq05ntglP
N88qA9uOoG/sJJXrIXOjhhTybBz8Qbr25pv3XFkhGFev4AsQiv1qpmx5auYO0MZKkXC1CBWS23qQ
CJVkXCMDI2B8bRje2XyGzXLRr2nuOIclVpXOOl782EMv+2f5jsM6yWu1LEmvHtXHpKa2GJZ1Txob
slNEPvZYxxdDFjDi5q5JOket5JD+GtCRVFR3tXsKQyjCtkZzfwwCtsob1pg6729BTckNi3dR2p77
VKVJ0muvQj066SQzWz2edVMh5dbSosefNQcUKfUM6lQdmHsRClWaI30oYGTmpnRtTGOis8whVHi3
eSmJqd9V/vxxJvKpZ0eji60OWs6X/lBuQrOJqtqTOyVFQLhYFD/vOii6Dj9mZ8LAbTOF3ke4MHs3
NZN4uMglFU3JYYNhX8QWrdhOTuyCFpV2KGOPf/RBkJvlDVqZBqw1noTVH3P1wiGCnz5dfz6y5CMl
Kt2edAj9KmNpuD5WG/TI+Rr5vZYKn+bJ3GFOfuGvs2HzSosEysJSJio28lTVCYOKC6DEsomO3Std
rG+hNBognT88whPdxAbagseqPHQH7Q/fc5WE7niYbLhfJxEDVcjuTo3eXW+UnRp3oemgJS9OTwUn
BTb1bnOK/36hx4A/MEsh1Geva18bGZnw7uJnpJeRq4JBfVOp/GKrfRXXWcbI3yU2Y9UkLX8rTD2f
2VimBAcxT9ZiJdLW82FZBa0v4RL25d88AMR7JF9pAXPgs53TKQXcx8vtVq7NQRka9YSnGvHkycVP
vETSWkBZFB9RXGIqNrbPYy2OMWjxDvBhQq5TtzLZ+Sc+2HlfF1eLxcP+Msyh411or+E1Gqx4SIsM
vD9f06LQy30snQFsnibGpmbBJl+kHsKb/f9poY38rAIkB+zEy7fSpdLqY87i48rRN0Z6nURFdw0n
axVYkBO47rGQuGQaFYoGYZNwckKrD9WmciLFPRa/mlJ+K+UgJmbFMLIDx/I9q8oTlYK/UkibEDVl
zJVJ1/GLgXwB7U9lgi6hk6RgRPz9AEQH6n4S9pfICtVOh19OJhm7+l7/4EKKrXw/4d57zd1AbJDD
K8oyU1lolPuIhhuRDf8MSQiTeBfTmWOWy7Ea6xYNqOPlAXQ+O/IDabUIBuLX16+qI6KIO2lIXaMY
slj4tCd0f8Fa14espYziobTb9tBirazffK5FSNh+YTY3yr68gCdgt3riADQcLtrLwCdgWpqN0une
3OMTYJHUwXYg0omXBs2/cN866tOSaFOSbMIQ/uxjg0zfTbufXke4gcWl3vAFbI0YqIolv6XG8n41
0KotxXBa3QvXznMZdfyX/ymYCoz0tTxC6lU7DfJ1YDqyLCHb2TyowMr6Lq5NrcO814EgcBU6T+54
5w2IJ+kN3gsGVA/IqMjD4zHPloZvzCRkqNaSitSRm/AG988gHZWuyGBi6MSvmDn6z2fPQedJiKwJ
az68HDVSUrrKHOJJWsdaMr3x+1M01RCalD2ckr8RksZif1U9Bt0omRXuCFmaIY6SBqiQGoXm26f2
L73dCfo4EjWr9Gq06haHNjdqPDLKgbIKh78FS6vp2mj1xTfKCtWHnaRQs8UmlFLTZDeBZvIf08aH
+ZGyxk1hng+0dyyxHw5ip5+eO5B+mChYQ7AOwp48GQz5Tl2zwWkUkPkvTiwMXxugrhxfFsI+/T+Y
ABOOgyo9KxH0PrOoiMd8RczJDHbdkTtyZxJLWXv9n+Ggus4Fn1W3+L0ZCxHpv4hyH62sfe8T8jSq
r/ixAptqKzTUIqyXi8BHbIwPu1UxrW0IUoRM18z3IssHX+4IqhS5WPOLX9/Y0fnTmhFIaFIZqvWB
iIdU/U1NJY4f2TlhUf/VpiuEfERsq6ZJZRpvS0S+GZ4NUn9WBx9J4q0KzI78IUWpoMD1/Buu9x5Q
FIIN2IzpaOnpDANgMkhhW4JzIWoPn3+Ac4AuYQkyPLM/giMzTyhLqx5a/uHnBGxvAoDWrPnPRsRH
PRUjARw2nQ6Sn5XNyZuVpEbej77UNg0Zd6Yag1jcrxFoyi7qQNmYaqA8g1ZhlsGkVqGdkKpbH441
xRcEjNVWdbRyVg/BwKyF8OsLXNy9TD7CHg6Sw29ZFPjBszv9QZ+OjYVt7UUwVKCV8xF+c2uuTmZh
bM0txNkTDRJ84XGulLDabN9x0u/JzayG+mWQSn+lidJB6u7LRMX6K7BZPBMPfBffor2h3CQu9eim
c3Dmpyk4pk1IgUDkzIKPNAoG+sPoMyBHnrgnATBB+U7vGHXijjc7u0lfgy43eK23ACd1W8NDcFIt
L35VJiTFh5I8kgH8gFYEF+Y6lWDYBv2IY5DCraYvECeC6xt+Y5LlVzMZtZTqHUn4n5Qxy+9KkmrC
48wc5yttwFtmSj2WVaRd/jUlxbkSqBFi2hcQl+hv8xIqQZUKTe0CoimL7+PK9mhuRYyVyAOarvPT
nST/GHMT7Cx3vsUONTAMzGHXikWMiAS/ms40wthz1FTqdBrseG4HsahxO4eJpn6v2qsYkbafAn1J
cQ7aQodJtERprlFX0vIjEWmBmQ6evtm2xkekwC+y8leFLLmU5oTUZBJMHmhtesRqg97h7+ekRw9H
DtM3mRG8Z8lggAVnuyf7boBFgOjQPxlXaOwa2Jpe7ZqSfvGRoCWQshGOVBTrjG6AF5uJJ+anHG/7
WNeN55cwLqX50tIdrKnHGdLcor5uAce0msbuVqSHnSfTeRLyvI2SeUTJd/Q/KtosRMef6BhFVbG3
zxAOyix1PFjw3Byhz2Y8zv00/lrQZhvfopjrW9I75BK86+5CWOia09dAKudcFzQj0tIRCwsd4K1Y
5eqcmXG82BfoJb1Tj3fOnDcucJk9jV4mDVGucnWNWhSqbYyBzzviKWGf0TFDAuFYd0N1e0PmuxcH
9GR7TH3n0vsV/dCd9xnehFZs3f0Z5tBGmvqU8fI96vW9Njh6ea/bBj282ziYCKkLwzg8K0p+bcLP
L2lNS2SD8EfEwxu1GYNjdafY8wUWdDGBgJi9dajuE+LTPFWzoyPMyoF3gGSMBYTQKxhZxaP3R0x3
mKleEV35eaMnRuPFcP8l5I7TWe40CRFAJGhTMLthwts6YJ0QgUHit+mQAwE6qp+POggfBUTgzQz4
n0i/eDcCo3CMzDtR7BuG3oRToC1EC5m/tRTJjgoGoBdDvbUVKUvzHm+2fiatO3RxaMrTiNb25C64
xLcMolhdjVozTnXBCspOA2OcaFeyd6M0uwMamN6GP/BCr7HDWVManQ6wNOoWgy5GxK+SG6QWkt8u
NjQm6n71b+bCMpmzyh7TmxiqG8mITWcwiaAX9WRmvkPW7WsKfj+BnfaIFPlvTB+TQyv1waiiv9kE
liYUEPap3pw3rjn03d/66gJlgD7YU9q+1QvEOpMwUje2nul/ueJlTq1rehAtNpJYp/HswZ+CBSWf
CtRTpn9lwX0cqB60OwRED1rXDQ+dzEW1gbWx0viUi0Z9mPawmSOaPy1m/ZLu6F7k9BxVyRWmAbCW
nATwmvP5sr/n75GYZtqKlG1CoHY8ixDzL7PQzKJUshglhyQHZckz15VWxY3b1xA6CxtByPc5YiJB
pWcyF79kEEWbX9VbQzDXFWYC1zxTULJVlu3J1ikcubrXtqUkJa2FeheyLtIHxiLamM+PzpwUcDLV
Fdo8CCF2crfD/2g6JABufSulfP2NvaWhZJ5eqBUrn5a8stZPPDaOPV55NZKOnDLLJcVBkEn0ZQ29
YmRSEe+sV5ltXl6I3RpxXjcPgc43VWjCojeHw7HmnLEVYJ0LmxAwXhdTLr5d4zno9IzKez06NhpP
K/en1zQQeVb3xGHFkp9kxcAm1kzau3cYbZHkqT4nmIfVGxjfcM/Yl3M5T+k97e6TPoBrf2BoV4d+
0rAN7gaWVmYvJkST3Xqi8tVTlXk7ki9JODpAzq+jVBGS48mEbCDWuDLypjPH71fwbEnAdXPGglDh
n0vWpi/wpHIblcFxfwhhUcyCDKJIQpVyH3HeLF1LN8mMVvEp6wPlI5sxMTUp64XPEaNMTtGjGxm2
LHDprEmm5C4YU0ykIJIi27vP+xFMHYIk+FiGLnTScr/T5BATpX4OIuxHSfhWhmgAWA+W2QmBfrcG
luw+IzX+5yOwo8uI0y0yhZs5MQ+M0gGvGESD3OIX03CaT42t+MCRB/n5VVtWKJZBHgGcFmfNmrE4
bFVh6tc80grN7+7FvibbG+ftTSUvC2QWMdIg0AJGZwugzD57Ba2v9eUFB2PHxU64g+rsjazPaJrk
w+HO1wmHnyYfVt1f2JLu65p33rJDrmauMuV6+v1SCyScjT+1tBloKoQs0QUwZHLK713CzVbphibg
R9iqW/zbJw+maoAdHi/NqdUlikA6vB3ZOEguKC93XtqN2FmJsKo2oQHdOXWEc8HU4nQKbcUhzHHu
lc0Xs356NsdNqS5Jcl0uaQjY1DCJyep9V17w/QBjiNxA0qvqDRF0RujmnJLYqyxxOz7HkhZfEkuT
TlMHn/qhYxyOMNZFhdsJUXVCU5W/aE7JTdlrah3PtP5PlbvAJGmOl/KWY7InyOKQZ/j0EfWdZFiw
MqvJs6BG0PotLFzfqGVKVAa2Uq3bNaR8+mYDoMQ6ezcbUcGhHdOPsH+KxIHF//+0cepuq/ejq+7v
16AAreCaXvzSdwyUvretpiWZUwRxf0NnehRx4EwQCRvvjdcVW/aOCXWiRTK4y7lxyvth5jhR5/3v
6jaX6/YX0vM40M1xpKCwIjOzR228fgYekPuSaDPs/WnGPGIo89th5nJbWGUMmxXycBwIjskhuReh
bB7/uyYhahH0nqDyGwv+871ehTtae1gzuw2mQHwZCSqhRmasWnogwGoZh7zP76EjtoOvmMLkDgIA
odN8LYqDLMNNZK/sZCbZtc7enfIGeUo6d7swqjP+INSg3CAGPDVIE73S/PW/mn2v06r2/y1gUlrb
wNBWTy8h5orEapToYLJfDnssi2c0w9s+jPdoA1P9K+TmZIR5YpNqPpqDKXo/62QXHitxmd5lfFSA
m+ZzvQ/THTKqXPltYiSLB1z2wpdh/ol4+ezRQbw+KlZZKeRfzoLPJj/gLwn6cJ7JTdV/gkAvr/TO
MQhrGOCzsymbG43Z6d3YOXs2JZZRTsyeblqxQe4D0rM8PWtN80KXQmRTQCPfqnk2+CxPkBPQm3uM
DgMbdSjxtozXNPrVlRA44C+1XK8054xXQMr2UnwEQiTUf5gfDMEvZJYFicyPalMisOv/ZRPufko+
GGN31nj7GVPnAFtdqSUfdcFTXMwxzxherypxd2RVcMHih862b4D44FGsXXi7OrEFhbAg5cXCP288
bhYWaxgNv7qpWuPKWbZ6cokqWu1/a3NnPPNxuNio7tShLpx6W5a5eOHvqVLydk8S3U5CeNfgtaLe
zRh+mBOQoWtpMAvPD5it2EiIZ+TbPj71/N0Tlh+4fjEjHilmN8GkYD3d68nZotQkm0M7DdOLpLkd
vm8mfuKSUDp207YODICXZjQZ3pQ99BsENQJttthBaFQYjtP3xw1evwUhd8RKFQUA6EwgWqCKIgTz
cTDyk/e4ROw5AHBmWkIHIwCAVGAJHLbUDVFQR4PhYbwi+QYPVAvYfyR44ZGkn4Qg6ZVFmwdjVUTJ
ulX2DMnPsUlQ4Fk5ExVqfzLc57GOKPjfcn2sJR3CBZ+l25c3uXQ1Xc670Lo11L6FRzo/wNIWb2IT
46JLWZgllFt63VxXd2nFQi9SN7rl6pf8E86rjmvsCs7JAlOkcZGzv76RsFJKO0LoRC8TfPqzuNk3
qD1mfnWd41dAVF1XFFRbHevhB4klB0TAhxsBXW4dSbBWCcVoFHGeTcAvx7izEqDs5QRj5sFzp8Ms
VWQywHa2gth5l8OL+og5ppu6KAnFN3bmMuOVBi2LWdmC67KA7IkpcBBgO/RxpYej/KJX+hYyKR+g
pHzVU56fZ+/wrRFWx/NL4F8EsXo09N6r06KxJTqVlx6sl9eyvRY65PEp9P2EKxQaCwxahPCBhnHL
369TmcJwqiIr/5H/uEocvp3tNAihhNxxV53vBe2uniLnWcxl1Mg+lGKrYJpK22oSEhekwIKEsqRM
tP08iUDLSAkByMLXDfvISfPARuwW4Kmq5sA0DSvB6NBqljwtyDeu+uCfvpGsWS31SjMMu2iTgJAQ
UOYiaYdahiQL8Z0/o9blAAvU6k4npZQHLHQzPje0h/WM8vh9QdHmstTZRPb5Wvaf3xK5sVnl6BuX
TF3fAlhNnJLYD1dG4gOs8t39ypFZO3XG+NW7wWPR/gsxVm5PkiyKHeICo3gvH5wPIRdBn4RwFses
oL5HQbPM0kGsm3rVL3MPi4Lxc7fZEV4JfhcWxeLulnWE20ZHFksRhBA0gUaAYgsK9EzCWRjTHaM3
A05KgSrlXqJFfAY0wR+Ug0yXiIsArORHgH20iiG41+Ij2sWvpiAvytKJcgrqCbCqNqYojJn9KMVI
/qZlZQsp1a94JlsgADK1gTwa/u8ZVpS3TkWOIs/JXiTaN/FwVDvEIVUbuqDH8xp2mfDokJofdH7r
6DZYPTJFjD9bxHR3GZVLQWpRSONoj26DthbMWIHabRHB804z7Y+Jr0YoYFOyexUrJxCdPQxfDXzB
wEKX4JPtM/a2W90PWxs3GrdTjj9npi9RZJfRwmHbdGpWOProb3uHLzvj4PLrTxdjEh0isJfYfEQe
e8XM8bxRNBNRaV6xTjmGQq8XCEXIfZLgeFojGJT+xkE1vkFtunhTk/NMF5qaA7j05vXZiyvxvbl9
9qWuckbMh3bTmfxtCb6OeB9l1L5H8+N+xJGQ8t1T7D4YSYaQ3i45alK1C011OtvdiRNWAt0KT/kA
p3UrRMBuOLHfG9uEhbhWKUHBA73oqBYB6JC1rmGVGRSrrrBYR6KieMuVIEWNkpvNeQ+xEKnbt8Wu
1FI/EaujltPPKNhuAJLbVp1hd7ubqL5yJ+iyEgbTao0+Hw11PKxsNZX8RjnHwnVW4QXZ1oA57igq
YrXKM7a+xWZ7Ny7shmZOzEFnaEVBcWcSvTLak1F367dFwspZnDoj4n6A2Z6yHUoqOOdpD74BX0iU
evu6uWeKEeu9JwlsdS6Flnfl5BAZY9W0o9QX9RGD+SXDBJIOmqUHYoCFxsUSYlBYk3m/ToTZQwUZ
qbdmZcobH81YsLolkot0WLoDLt0HREdBnsgmw0tN9S6Vy7FXmrHNsEIBADzrMJNyXV1FzXJROIzt
8G5qk6j1H16WKMbHWC/wi5+FZTyyxzUgoz1Fd8/sxH8O2/izFrasWGKQsbvpS1wWaw9r3CCDttFF
iIO1NQbJLtE+0hk1EcAThbSjppXDAde6b96Df3ROnSC4KPDQYVb1TKr85ECQwf5+FyYEuVI4gmTl
rfIg2WkrzpocMTr7JBNFMT/hLARIigNw7GCaIlUudYwhR7eGQ1xe1F+BGhdhmczqH0zdTA+RAi8p
QPrJAEG1xX6gMfeHz00cYDoo8mzGtmRHvAXh62DTHj86KXu8a2g/Be6n1WAwyBkIjHRLp/LYitNw
n9WYwv9LEihjtfdIl00vPo4Kx6zG1TFLdOHcEUmFMlIGH1sBFDZ5XOS0WTkdslHQ5ycTw9Ruvk5W
MTTqR4wPlw3w6/LUpkyzB4KQku7Eyv0Zu/U6NdEgqhbwbsAwBm8D7iOpjiqN/dXJaGJcYoCPMhd4
KdsqBXuLrlk/UyTqBU3gg3NdVpOuVrQp1es+BqGgzdWNT4kihb2od/TjPDIhm+56XlC+nXpd2fsQ
QHQ7PYbdCD+sLDuhoLKsnTOdGhyJ8vC/PiESNhF6isty9xNJvSCFUycZRLYAljvAqSLQ+P7PmTwW
T3rgoncf3afHTYrjMKMaWMh8NI59WO/9zwaDfrzzE+UhfyQiSpfbvCqzJafomqDiH8gLt0rCxsf3
kSVs9w1eLw7yTQQzM8sRyJ867rr97a4L4ZGWERg1s4T+qW1MGce10QsEYOAaz8R5uDjuU5zfEmBK
zQbdTnfMw02+vC5+OlPN15nZ6YcgISiDjUW1YUcLIt3/rz3Y+2YdORv5LefYMOr9p3NErImiKSgE
DalFaClNc3BGJ1NSowTvwuQbQ4e25gidtZya4Mou61aCjZRrNFqHqHQFb2Ziio+MnUJWiq0izGUp
569jhpdtzyr7NiTDtLkfJgTU0S9MI5kqhIHdcmexdrWmm3N1PnVQcsWSkuN9D5kr3eAG7dxjriAE
4FLKZitbhST+NCmK/BiSIeFtZk6RvqktNeEog7G2ggXgFgSCDQF8dliTF52u3MjuuRBEDFy8eEme
3Ylp15DPuebGReH5BGvsnjKKxiEDSISq9GS1JPk/bxLChN6WyCcEe/5k+2KBIAMV9MozLZqc4vzL
getWujsxKJTIj/p4cu91435T+aUbOqbAxEkkF81AFlauisrQCJcK+WFTJcSAHFXEGPgwtsB4iVJ+
aT0pTGIAgOYKkKo9O006fnp/UZmWc2rZCX8NoFrEJB7twB3se2kvYvlP1IhZJiQhe5RYMsoQjp90
kIO62FVsB0vHyrHBRNGHVLjP5bdMmEwSe+C8KMCC4/mISekGx9EpbKBjWOVlJL2pn7NXIiFmF9Xl
OY3LxCFZhSX25AaryJUYpyKUEqfGFJpOMJNjbsxkq7xCwi+cEH8sN0MTnJaN/LQ0vqvNxd2q6/43
ZP2OTebtUIZzLH6r0b5Sb5icLBygHt8HpF3Fdgz1dG3ENFkGnybbJyO2FfqndOQbhIK5k7sbhY2Z
ZZl8BWKQfTuW/4uEea1n6xUMHAQ/7xUTLxY36+j/15qQQTKGBcpVFKSIwx8iFV6yxyP0sE5MgEAd
E6BDJAcEoTn6hD8SvBQKZEeYHpb2DfBNnIxtenFQ1DpCU30qQMn2qE/A3mXq2ddIb3ttqopALW1M
M+V+wBiy5RV/5C6Xuik3Rs6rTgmy0D8hwPM2jEYPGRmPK5MZ7zYhAKuuTwNsiWFXtKRW4eiOdOyL
WfPPNzoQCz4m0ptJaUhTAdaoNPfWrdn8DQNejMK+1mj51D3NAAjYvCdn6lEfHPmQjXvPFVilaVG4
Ke3uTtxrJiBsTXRJ/x7QnwTdWkny2nKQ2GOrHW7WJAdw6340kMVqRWmy6RqwYhYgZPS2pQZKe6g6
v9sB6EppgixclQ8SS97lbVAk3GvQYDQxxkUxICc5+kS6lNQzNqE7OS2Wkoqk5dXrEzF6XALw0sqb
v31vOuTQpQ/tJmEbgCuRHGUPimQQEMVFXRc8I2bNNzQLYLLEV/3x51q4N5JY6GWBxzl4RzkYkvsq
PwEUdjFEHKBm7PXnf3J4lL3CHhZdswQL+hEPiM4vQv4bc23N3eMrPXUq/p19po9q7UXXRGSwlAQi
e0rO+S4AXdwm3Hd0psilOWM4VBpMHDyl7qUfgexXqolIreDXu2LKX/UA0ihFbQaKUMdTqi2D0zXY
bXQJkilAJKpST2BIJzknUVN2VXERhomA9TDaGP/S9E/1frPYakAXJL/iSKvOSPBw86zEfffMf/a1
kVZRBHAzw9CrRE5Zmm/3R0MFRTO1eW8jeWFot4vdNk+xuK2mDkcYPPIsft8eRjcOMrlrTOTkW166
mjL351cLMZvA0IKRrhM9PjiKCBpdKRtQ+ctY068Evs4FpQsgvXOLEGgoatEQ09bzyacPHRr2YdH6
/DGLndhwn0SIAMNiUPigtrUVHFZlpjRx7FW/8oZTcJF8NFM3ZcAw6t2QiSfWziwdoPTHfbQWb0TR
XSxA/QgwJzGo9WXPvsPCXJv1V4IjwRB6O8e8fL1CLk052tpcJBWGLpWAacQ3aCFynzUOpJyBqNDi
Rc1YZvGr7DsUUj8uK7GxJ9VOK7gF2bozf1kgNlcEQt+1Hp00w18b0jPBX/vzSEiiRuisp9DBDbmS
UyI6RTP9azbWAHHFwh6JPDhxnuSlfFQ05tgb5fm0WxrK/Xz59R/HmJ4OGQMptNhJYV62kbWkicOl
Zd6smEu/Xj6cWyp2neNvXsMhdSf6SbdT6hI6gYcIONOYVYa5DwVowH5BHBOyVCINRumBgGd8U41E
sCNIVLjtkr0ok+esyGAbn+yMq9oF6I5KdRVB2ewusjjDhENgIxyb5mwYnijSS89WmORV8ADBfHOj
VXlYmW1YYA20T6s7/8hovPZuqmpGFbkNDPQ0FYvbxBYv1uocArqLuoxDumOQMCALHhMtq2rvWees
vQ5DBy8kd7Q4WICQh0rl3UEO1TyBMBV0RNNuVGIRd/WL7NjhPydBKiruAYhnn5myVWxxYU1VPbpi
6X62urQxTGGKMhuMX2GTgvIBGpLPSfn42KSnwN1jR0OIGL+1rrfFgnYQU/4TiVvHwBDwFGJXdVXJ
UySe+7YJNwV/j5xF9J3aSQuY57nfzh/ZvYMZ2DHkBJ5geipkWD6IalVEBEToqOFVDJvD6OXLGMJt
FUaY4u4q5UXIUOBy4X/rNK/ril6SpY1X+F3DCQTIYMpzc8/19sK4xEd3rYuz9axZSOTXj+SLpch7
3Q0o+pm76H9bBilQdJ+wTc8vImaEAMkxeIaIVIK+HHyxydNSZXrAHpipBDxQL4LaJqfChVwpHwmU
G8H/s+IBvB4E/pFJzfpTzEVOiOSn+yTy8px6aMZ7dWECnmIJtgDgTayKWV3px/7gBmASwGMmlle2
nv0Rt0Se+pk/SnlGgO8YHEv3aDZAN0Nsq5MCkAe5ZWn9AaFsbo2W29QRg6AWtZ0UUgRwCeHUB6D6
czuiaI3MMF6DoRq6gb6E2/sDEmDRAgbSGh4twQjzYY5siAR3gOphW37Hm0gid9WHzas92KJTKMUc
Q2/FYn5+lBlXTJifbz04k/vXKGIedC412aduQqLy1XFLHQcFZ9bHrOLd5qw/0H9osgO55/7+V5v2
uqumz20cC+0T1JDOoHSlHaLQOcSQSu9tpG+N4FTYVFNcinFdJNgaWEo6mHRaJm5HnBuwAH4sTtUf
DHd8xY7d6T8/swrL4vaQ+e1F4Q3SUI4oB6/1GeNgJLBW32Fe7MUj1AhJ6Q7ri4MnmQHHAaQGGnaK
3NDRgQmkbB8y1JEMA4pSnZ2czUoxA82WqOS96mZNAOBmSFnzWUEkPCjk0NS0mPyC46Y9ofdju8pQ
LUiYEeXS6FFOZOWHr4E3HAc+ZvB8Y7//sZN9uwzWJUCDynsqu/plcOpLmtSxuSf5VlDUpzrjW7ad
Mgcbtz/dn89otB3L31uXmbdRE5KNnl25KJZ3zqBt3Si1DCzoNlVstIP+urKCf/4048a76lYJxAKP
/rn1Cws+32t1HT8rWTWSaqcqryKBCpylPNTinWP6V+TgmGGj0QFipcIEGBlnXMBBmVzeBDtO/kcD
FpMN9YPeuIGHWfIihoRD5VVH+SQpR+MZpiK80iZEooGsQKaYePTj0rV/c9n8juJ7lbHvF5iXjAD4
n1Q2S7w7Qfwxu5oqmWvaLvHC+dotdapmWV3oa1Y3SVYmzW37otdeIJcQQofcLS8A/WVzTeeCCRzN
LcVdMFRZQHinagN1Rz6Acq1mRg4YT/J0h1pmHWQbgZbYUto6rWNeDoQ9KO5/pohvZRvGru9lIypF
ofhkGLMBHOawfzvWHOEkBo6yrvkXyyMO9SMtE2G2taeW/lFNC/iPfR2Za9PhEtRTGWbx9vO8+dBf
pQrsarjmnc1rBVI8Vxofao/VUb6eZ0g7t4tPdEDYGt+pcUGbqyYHuOdvt4rl0AQeTM+8KaDzRSeP
4lCsgR6kMmnVG6fy5OASkvbS8AmSFHMNr84yRg4NUj1vUNm43W66GZkVOm8h8z1Rsl/c9t4V2x29
dOCU/EegyVuwSQsJoChYnNinRdJw7cKPWwtVbdufoS0BGBSf27xUPyQLvOt7iK4oazespsBszFyx
n8NkPhECuTortZiL0pnGwIxg4TZqayNUa2CcPTglYC06feZnbc195xOmWNSgK2ARCUkN02+ix4Hz
/9UnSslStznAoKisqJwxfkKRckq1xfIryF8hrANehkuDba475/w+KlsE+98tLJS7gsdTqw/62bOQ
pSEmKlF0xXu1x7Ku+A3eVpGRNBvJUUdlSvqLGsyMTfUBdZlx1XgRPQWUMGodmoG85uHfZBKE8Bks
KcVtIYbZtLrFiCjh9E1ztZlmQvW/ghv97jdlwZ271UafqJ0WeEM+Pp3HYeopUZhj7nYPZqWEKQoa
IdJ+r+MmbAU6Do5YwyFRM3Re+tG1E1Eg8QQYjCUckNR+5a+06Cw9BKP7qOZpa4qWZ1R0irkTA9Ai
5WwKsY5DRdQ3uD3dGaFIo6aCaNmWvYE73jdwg1q4hTbvLuey1jeQq+46/3PtjSKRCmv3KPDSL54o
Y2/umQ/Gsm2a3PrRQQxvQaZz/K9griBSgaMUQ8/vPR9ZKQxfUb+WLWGawWRAWNQglrmqeBhpVo6H
8GLAb7LUTy5gIggM3Louwue61yY96L1BNWcuhHsbjeHapqmnK+Ljj9q+Ft3Wi9/awJky2kduU/9u
A08L1YHRSGawokCZ+BdWbpogjcWMblHBG3gXcs2FjikvdI0VCasbpY6QsC3LOLwbEcRpCuTm790S
njFsQyMGPYHN4spQS9XtrfeYNIaACjgPYWYXySYuOTPL+1w07JUWYTfGVh0Y0INmlFmjtDqfNi2N
YjEbzWsXlPHAex2DetJbKdcgxlaUBDSgXabVCH7jf/lJEEcUMvBz5KG8fn5wpn1DRlmcd56syDS9
Tb6PgZ/FC0r0XPsG+/KG+SqTm0AeBnPTVPUbaCaqNJWaJ+UwDjkfWrrkhTkiOCP3bMsnGGosMOQL
coDwb32E96pjvnz5vkZysM4Hxw/D4j+r5o3s87un4lLT/ri2Ow7j7TGHWSdfRsJsHRdvk8mnfgDk
dbfGuMH/CaUsbSBrGe66FaJMMSGB/vD5prEfC3rpFSwTNJdeFqQu/bmvOBerI/oUelarSBEFPi+g
b7h3MjkG0S7j5gLo4BQT7VCTCh0gRWt/LVq7yvgvQrsTecMzQVdbCtn8U/rwvlJTXbcGxyZ8JrvU
UvgK15mfKqZllVO6zd4KXDqSyDG4JR42GQ2wVStnSm12BCpK2VzjNHf2Yn+zy9iW9+Xs3yKgG/S4
9oaHtqW6kcSDKcbtZjzISDGYSxfjXNjsyPKgIke+KISKekvWQYZeaWWIHXoDnJSGc2vgCqyarXzX
rWEleeVdwAOmpG6avPoKYQ4fem2Yac+pgAT3mOmuFErI5b99J5nyjZZvwvV120KOQGjD72mLtK6X
vVNuh4yMaYvBn6WBQLwveJjV+JYtkNM6lsXzrvjbPRLWWb7zrbqi9fhofWUweg5O+agIp+b82ZCO
M+BTn2LTpGFProO2fMx99fhHSJW0Omkknhwe1lX57/hx+5luZjMNucqa1EUjHjGVqO1Skf8RZaPI
2maT9pvRGBUmnvqvygkyA6/jXY6foHIyFNs62EDKWEIg6v4nAAj3P3OtweFMGMYkjmo46jMGpRhV
vGlwkrwmEepEp3dkzZhI7UFeF7C9XdYyEM3cLySS0dz3/2Hn3EUvQ6q13Tkgcg71J8tUWFzUYJiU
uWJDF4cX9oukOk1PWlBYgSd4T5nZp7kXLBhssF393KeecuPX6WzEz6pzUk9SFYV904lpQEhfz+rF
fHBn02l0flEotPIMXAh5eGF41KbuLM1tlV0GuCkfUjkj3f+F3g3ALv7i52hEOvI5r6Pa5nAI9yfT
3XYeNvsIToM/4aOwLJ36UAbGItV6yDmXW9+d08KOkpxBkpDBPjb2VxVs1Zl4YXLLl6iQVFfRPqh+
ZnlqmEdXKFJgIXu9rlgRIp+lDp3IJtIh0waJMwi2r6dj4lqc9H33s54LicSYZ8bez5u4iGRhZvq7
vPopCJltJsnXsot7gOR6f7MD6pYPFOD4Oxeb0jPO5codoQNj4fTsdb54yFDz08skNYUSU6TsoAxb
5NGdFX5wt/YjwflAKzm3SxesijeBRrFkqfmKs0wRAhFrlVwYVSIylKWA16284xUPDQTRwpQGrmcH
GNOGJRGqD5SfuP65rGVICRU4z9n2crt5bTjq3QdayKWW5ZzTWwP0rt8b7WmoWuWF9DFyllxeG2EQ
qD2XWcPrHNMRQSBez+wZNZwjI8U+TscoM4PTkvJZu74ARDyYBf8SU7NhXzxj9Is6Zmmzd/8dBpS/
H+E6CMY4KvVkTaFKQujwBg/5T8lQMYYMkqWFCC8aUC+zGaDd2bqpqhKqwSV4iHnWAdnKeImX65x7
wZ3XE4QkF5cwuIw4wvQB/Z8dwDTbFX5Es6SgzBgKHyzIeZXOC41xqzqZXIt3Rnsu4d4EhH+0VycN
ZEfcE/qSc9F4HhXUb1FsSr3cuO2qj8yjLcLE2AuZEmkfL+bnMjUTCjRu0liTGULy+dTDWEal8vjU
RFZUU4/a4F1ipEiYCD1vtBj0mb2F5F9WH6ZAfxlhu8NRrd/kJr+S1nX6nnV08hVD7vU6sFANZ56R
SlnfqIJwQhXzWfSQPwGERMHGqrdCIOgywrXvQLyYnkvL6WSR1XJFonYiEAsKehTRrhBlVmahDObV
2ztv9KFBTeGgzvv+GS6OftjYx2+UP51IOmQyAAke7EAd/hnIWbJbt1uP7E+63+Eu3ZewkThqPrhk
3LZF+Vo624sflDbHlvPiN/l3A1IW8Q3gNJOrf3t+DiVbQz+Yasjh6Ni8BPfK0UZsIRAXdZfLgD4e
VeAlJ2HtRiBlBn6vuiz0sKYbWyjh24M4n8dWvf90R8AUJ5PXrXhi3PQoVUd28jPUNUp8cF2sFsbN
4bAbC57yO45C47Ofgra7vg+kKIPkWEWxtGjIt74eZBF4g2KWkbUINbZHbFonOl+i4SlmWBrl6JkM
4lYuNy7ApH298v/8b4Pv4fR3om4ObZ8IKqpiHhm/k/mDTiF+WjEfaSD+BdoZ2Seordh8wVIUSB6D
SrC97A0KiJm/SVfT5UiR00zpH0z76+3VXqCOoLMPM5bYeKDGTw+7/EBe9HpsM5K8VGMxKxUjC3/C
QGjwe4CuwdyKKW82l570ozjsvQiWNia8XVd9ca33e/FF3pBCYqS93iho2jCg6yerByqTEVjdTb6Z
oL01+uNibeL6GpqY8rG6W6+H1iXJ1KqfSjywbFPQ57jU1nOqW5/YHbJswv41JvqTp9UueWxam0tD
QM27GH7dRsmrBwGfKSYlgB9PXIJh1QoQSu52sXu1+4vDfP8/fq/fNjyqbWnnNDItAsBG4ZCz12Sx
1AHSvLy5udn9UP0RFdQgrsUy4f3WpGgIOJb1XV5aiu6xWKO6HhT1xKrnH06onHaj1/QYd1OGXJS5
26WOS6YlGmrCb5oSi6epaokcKaMq9/BcRC9fogqg5BptS6O0iuJl+l5WFUrBZp1H6P0DOt9Y2h/p
HgiGme546pHtTpzJ0mjFqlyyCluPUqQhgtH+EQQfYk4MwG6WFA5ya53uN6W13K+hCCQHHkBM2xfU
z1BrnlrNgdYwp34mslQhl/Sky9tqFRvTkoBJ9w3s2v/0OlMw3No3q4fYu7yESwSKIED4PJr9Gd2Y
zFRbTEVUpLHSdErueUuaQ5X2c1QITQEXND6eEB0d1Xemp74qemUnNwnF4648d+pGkSaHIFlWHRWH
gOr/GBbYwBgQe+QDRnjlfCCwBTb3jHqM3YnNdGEIEe4kDShZFsUTbdiLc9FRU5v6prmfW+AAfSQN
izr2yaM3nTWumtlKeQAR8nFr8+rmLoIH/FLwV1aej3suL1b4D7EJOQofeA+ZeYbNB1ozPiJM+7rV
m10zkyVaMFkWu/NhZxafRP2MRSR/wwFdqTbu7IWKfUSMlDtEFAreJtolHRd1vOmlU9DdD/0lyO/8
U4O9xGzR8XEJiiofrEDTSQUkgrVTay7w3XbTjZFKPLmLNGT7K4KOlSqln2JUBb9T+z74qA3dkVuA
wuluEs+QIiaEFMgj0iMAhtEUbu+qRfX+f0VnTuEj0gj42kbvNcs/RKLTIA9sSoSouMD0hFpAjhcr
O42ZXkEHuLhL5tTtFg4qAP1++692Vj+ViTK6X0SzU+v8qDicPFFdD3fkmZuQ04YlJc5WhkNio87m
9dnCjJm6HBgmpWw1EuBZrTIU/sIWOypJkiFbItSRuZQLC6YzFBKmg0hNajFNkLcqmWAmdT7OXttF
Xl1MfBppMwby+L3z4qDcftR7v5v3ZDKa5iydvaP5q3bpE3pne3yS842givTM3ttwUHSkvsar9S9k
+0litIBlApa9+nDqDQjS5zK1fSjkLY/6f+/FaZD6lZ4/NQMpVFFDF6KbvwpWpjuF9w0EEJuyePN8
IAETvSImjDhOnszB4gBd7XyyDs0b8A5z/tXz2z95PMEis6A4jNM6VzMvlfHYt1EmbaEhaZ2HTz2b
EAICFHQXVih92eaJqI310bCCMhu9U7/6f7oKF2XSdzjqwROS4ATgnzzZLcpAcrSPXRswsbpDqmfA
3PL0VW7AYAB1Ds7YPA3WK4gEFEul725O+gK1FbNSHpatG7shpB4wQZOBNvsj+2l+HIh2EA1j/KuP
iv9H/WI96GMnfkQZdWUtGiU89TKB7gVwpOydLXppT+rmwLj8RylNUkxzqzSKKQJ3Zf2Pc5VbDxcq
hr72mA5E5oCThYBUVclNgFEx3f4VgfcZWxrUnJZb2L5PHI5HRS6sQ7gXe2+s8R9qw2DZ5XocBDQ3
LrdxNLzLfXI6NWcp61277f672AVAl+91GK5GCfQV6tFXFn+9LANLfI+pri1jvrt9p9ZAckDlNMZn
6nrt3FOZKNViTnCJtRy/oppmyHqx23OTzeddA96q1HemQLamRirpqgvgsKvH0gAH266kvSbkUBrY
5lnwlQOzlOmtFc/8k7q8fUh1+jWjTHAAKocOcCsHyKmwovsmYNwncB3RmSu5dI0/AB3auvFkAvUp
oV+kGrTQVLw82YO9vRlf83Ckm4tJ+VxdniMgKeZYoGlHuFh0whYKPEPia28O4DAwS0qEovv5iFJ+
0FMC9zmC1I+XiNTzCR//1zUhigAMllZ00FV5f4NAnD2IEbjHBl8Yfw6h2pCZuc2I3bOOsEpGYCnt
4my5Dn8oP9cicZ5lUbe62zd66bzhlPbQC5uptn3tY6YgawbYrpNpQgHWPpdsC96Aj/TfEmF3xMVB
ohpOZX/EnYDGtGafUHwx62sqQpp8vLytXh6jZ47eHmIa/H98oG7WAoJSSYxi3rsueqxHoJdI4Jh9
kknebRIEHcrFXEDUnrgZ96G7HKPJTIHyXemH8COvpEEwF69uowzs6VjibPqO3p+ee4ROVnYqOv9t
Nj1u/6nqywFUmYExOK4jW4eLakNy/Z+9EWoLI5MjUNSduJZmh9iCObX9sZbfIbEwGC4/A8+FTInu
qsBdSyHxmSlV96bpTtvEsyaxLEg0yYSnX38JBB0FJwfFuTLjQdjWDFdQ4ld7V5IHedFNljaEwkJ0
m4d5XvW06Y/TxnTWp6mVsgrvmBuphsHx14Vl6LiT0jqCl47SdyIxqw8gEmabttX14u6Ro7ZCuVYu
DaA+O+YHczqCCHa9ABd0uqaqRKe81YAC1ErzpJ2hJjW1wvlOWq5IeIt7iIA0x17A5RSNIRqVnBy/
9HoeLwH542jfI0nsrnTU1KRCBEbSoDmWFjFkLsQ4LSB2fXsqcyTnZ2y8U1mNt1FcDVEUyRBhAALw
DRD9tTTT6GVqBdjhePBSSh1hXB47oegwZ1gWlxcsA+kS+Mgarnkzc4UJriIPyXxkJH910do67kPK
8lho+hifgTWbzG3Utb8yjfWggbsb6xDYL+F9kcYrs4koe2e/Ehjx77op4k1GNgd8UB3nwphqQeCC
LxI6feyotDxCRzfrRonWkMndP5HW+AI23rK98Dv27ezZuHcDA5NKh91AtUVTLM/EyJP56KPfDP3Y
7mdPevNy3o8tjjoRzxZGBmUwNqLDjDsu2FyEjRcfFlJKZNDWjH/ChdYZD7tGhd85jQKLsXF0CRm0
cCHO+60F8q+xvTNR1HEhnTuoTfRe9AZDIWWEZUoNMnJiOcEsGR83YaxvvmyL1+mKQzr4udeotiL0
KTT6ygMqM6MHD1uZrEgarOrGmtl6kvGdUzOdgjHjw1AHWrcJ8Sra0+Xgvzi3Mqpj10nV1X4dA9S9
0GacutfT7xpCbCt5ebojgvwB0KcwlsVwfSLe1TujBpOr4MWNVqKOT4wRMPLt0zvYiFHkfm0qYGRl
OTSx1apTj0w/s34btiomF7QRRUETJJuHvmPujCFuebw6zznaySqDxcLMxvg12aoeJCZL+sDjEqx1
KkMOK8qu1sdReJh7+08uvqOL3Ze+WdWZhgN/Y/c8V1mY+Lm05i0hgwFVfhhnOn4OYWqalpjOfN5O
EK0Y69EuRDZ3ymXlS3F1emwkwq8uobEBGxUtRKjXpPVKUZ5eEz7vacDEkTLGpIv/vTugPSJ4lvw/
SAItE0RDVZDVocgUHYP6v7x4eSyzLd3PdNEBSHmJbZztd1R0MsFI3V3uQMG8FsmftUXHp5iYETtg
eDU73sBt8dHFYuVOVmZo/e+GRId4+mn9A0TWTfKHelKdQWqkxCT2ZTXBFPYD2zLU51s40qsl1fKV
25OdepggRon+/92qT5qwN9SwjDuGOvLMb4RmRLSOg36v1XuvGj2j78tGR5Bvcy7c+uUXNmmJHkya
cQFUuWwjPm+F/m20vXmFSKJCcF+U+pj5wO4/UTrwMD5BR63H7etvyW0WsBeYkH0EiSLCTs6xyHmv
qm6KwqK7qO9YPWKOsAkZ7VDffsrvkSP6Lwe1toDI7dWhhefQ3PK4/9anx16wcVMJnVbrCKKIfNXO
i1E4QQ6E8bNSBKJjHGLrLDYXZ4fHofHcAriaMDDAkEg535yJ131wOXhEOdtHkdTzmlw5q8Irq/q1
pYz8s2wIZfLmofkKmS5GIu3WfmqBbmIq7Ai8NkriY3FDUJSyCScPTICNv1YSycxB/EU2RDRYIOvv
HhI6oXYr/NVsbwVf4bQpR1DXmGCSDnje6EW65l6iTyxo5O0HhmnJ9vpXRhjR0PcZH0/ynaksbwRy
awnU5t5+q+DEbINsUVFbpVLvTitiaLJtWiTxOM4e3bBxH4ThWtLh8hug3sfwpS8ckIq0urN1tvgf
Ekr3aRFPuErJoV1YxYH8iFjC/rHXliO3uLinTS5UJNZ3qU08PmQr6jHhefBwMRtW8BieYs0XkqgW
/5EgURE57ypJYZiJpZKszF5ajvZ47Nly2yfWymnY3YgacKMKhpshJjhOjlP87/AZIe0ptlwKGr/o
gkuhqshkkEHxM+LsRtSlhCARKy2XVIkaeSp0zw6Tbk2hr8DakZWxCHW4bcwnrdG96qJPoJeLwAYA
S3gnc2O31xXbyNYTAiHX645BXHecipo9GiP5GLisOE0jggb9yi6wSiuZOQCahOz5PMtHeYy8g3u7
2KUdB8I1S2V54xmzJBV9AqvxK5k0iBoNBVewMZkMlJPkywpmv4Mn3WQwK8wBBM3owd84gDJwT8+z
IlT7ARr1OADe+cK4jgWkHcQZJtx1CiOklG2n+WfftBTjTRBN9L+ELQEnj/VvKhb6QvvdTo9LIY3o
oLs1omDXhyEZ52CQngWMQyzbdyLd670b3Tj1p3RAQAkDlC6xBPSGIfRHU3cJN/8yapLjaz3d5K4e
PN4iP/37XjzllPjqf60ofGA4RWh/wYS5GhprBdC7s4RWy0TY1WqjoRHHufdgXNvp1+Vr89VBez/T
/9neO+Gn8z2kP46bieWhip5fNa2Arvf/vOlh2zEK3d7LJD3yv9aSlg4LGYQQgOq0qKyqEZq/0j00
B3C69TxCDZWar+7B9bxk7krsU2NsqrbVgw/f3I14dgyQuLegKMb0vA4iER5UqI7cCGPYBD9KDY7g
J9vtznKcViWCc7dwI8d5mQGEKnkVGRgAqW3BJ3EUf3pa+pYo0cowXtdHQQhbRRxgzdBjmgZV/yim
jQAFM/Rh6eD8SZNTTsISxTrdcod72gJJdK5DQ0dODzRSJGw6Ul6oIM+G7D0hjAkq2Rq0k4XcoCYZ
aTMh1BENAXm/nh5GG7kIwPF8XCQ/QJ/a+VpvxkjDoNvtAi4bDxlVLAWmzXpRzrASpdrKMaQhZQHS
g7FIyLo5DNRQUfukcjb2iMKUSIXSOOUwamzFHAI2U9TDCljo/b24J4iguO5LR+7mVdL9FRUViyl8
0XiXO8KLyLkDeUiZPiSdF8a5dZhiEYzHWb9JKdFjwoLCrkClRRVda8kVS8ijxG5lxVhQ9XMBaNvO
u64QuJkOakFyic4nhWULBimQfqAAv1s3iL1BkgIm3vfy6JGCv590VhdZOELacEhKqMG+c/oVLv8I
JTqLYFT1zBBcuBP4Q380Ec6VLU1nYPPZWDQiSyLf4sv9ZCxSNu4yDfG0ZGtEKYMdVEphR/CcuTb2
DMvfjj4rpLCW75X6CMxAuk1rwAYW7OJ5Fbi1X+01NcaQphttWhEeomdZL8zMn1p27gRCWmnHLmaq
PyzxpRmBZl5LsgHGQZ3HtNR8TMu25slx87vBtebHScaN+LITcq8AFWSU4UYfxTpdMpLhISBBagky
27EK6Ak/Fni4Z/OTiU90hvWU4AzFzxhw5W7ANdIgAjSbYIIREPpZjdDmt+JcfGeUHB2MSA4VNp1d
bZWhLdoceNkzlT6lNGXt1RLHSgFLw9pUhn/4+iRb18quRwsKxbAGrGzhfrm8oknUMsaxh+WPEdGZ
fcm4LLTCi7JaJz6EE6ojG/BCiD6vGTkTInDy7WgGCIreJwu2o+kLnJ1IoRHM648aHZiZDkqg7t1J
ZZcCYxugD7+icbFtYnKFq6mBLIHXZowSuISiR1ebaart40J33XdLNN+nGQe8RO5F9V3oXVTxSQGZ
UjVIKULmFQheU7Swnc6cEIbCskf6BA544/416g3QC1YRSanSORhVBoBqvS8Fed+OxPzvBvJDeoMm
WIWTjRf/g9AaLVZqgku5V0hnUekPO1H1hvnRcK055Hg2yEGtofvSbU8oeJz9Z/Gc9LDs/7zE4new
c6MQlGcHmsSzROfUl5iqvc1eKqKPg/muPlxaZsO7WBoY1Zv2uB8dhBltmIiNqQdaUZ3wjmvciyvF
9QdQxXJ4TYLIsLygNqKhrIWQJgwEZExzgeQAiZooflq8lItsHBLJZDyYzt8CRVYCP1Yyc+Xsx81W
GVZ481+IvNokPYHMf3WTWyR4THajLYllkALYnFYETqNrMf6uvZiXrD03n9+cqcoFRdUI1DenxMle
6lwLkOcXWTkTiPQ1PYf7Inx6wVc99G7VwB/QEKSONC0DaFi5EK4ZhcRTMCSuQy3SNR6QBJyZ2vcI
tUFeZzj2PC8fcz2TOj+wGoFQnHKUK2cSzOwHjWoUK0kY4dDUQucj7GcHp6MnxFvGDyPa7HZNT7AL
ZqwyADvv/HHWCFLnNo4plA6/zc1OBkDtrhwSICQfZrSTm4hED5vLudbIEBRPiRN89gLrccOA5jfe
27JjYPQjDStI6t+7jr6cLlvTNzxFudyvzI58W4tw/J9Qw+FbuLCzWGbqB8FffzAPjBpT2qusFp0v
C8Io+EMnKsguW/pOmFOuLxcztnb2qJHqIf+0escJbpyjcZvREtKd8tVgxtxJT3oMj9GhfTPqmwWB
OtwA+Rbk0/bROA7wWyPs2KW+r1HpZPDnViQig1FZOgjFGgOkNeKn6VQF44agA9t2nLg43zlSA28w
Z0Dus72ruEjlkWSybXTY9il9d7SbTrBbY7P4NC0FHt2vrQW0kTk0d67YCPScfZiTyim1Cb6rg6ZJ
A0mHhACtmYCe5pHorp6Nfwj+EVNpMgO3dUoVMHRLHfVrsXgFix236SSgcP+/s/gWFSWKEq/FGF6T
AfzHulD/c5MFx+/RG3/wSvYx+md/HTQq6+11ntlxJ78bFXFAQ9nVkubXX/1xaChNUxcpe/ZzP4ov
5UTeiG/xyXZSN4qR3YhnvxSDWrnHtxcfrjgxrYvbLlPS1XBnEb03fmEu2NrKTbk4ZjVzEWdZ682A
xXbdMBwlQrreazaaAXP79PA9mxrQTbc7aRIpAKtWM/nUxex/sEttRnfJQCfe1qDIEHLD8CgI2eug
3ptJnkzi6JObpuF8XCtmx8RML6CgDGHsNgK8uyAEjg0NSQSIG+XaI1pqK6eEETs2C68XiyMGpwwA
F9m57kXAi4vVkq8a3Hqb6//okueA1+HUEqpvzhuSHNryBxLQWzvTIIfM2244eqbsptfBkhD4pdJu
Aj69xzCmru3oEBZCwWo4FwZ3e20SSYIMdlW4ApTU5VZgoB3xbUE36mYW0n8v01GDTQ+tSiv5gCQ5
3c2/fext+Li5hGfaLdUs/G5+aSkU0Chjfzs+SYshWTvwbcHcs1dS0WLjCpclH+x+bcSP0eoqHnF0
Knr5SmPh8HJOxaFsnW7iNorUqavv2xRTAxu2eKcKGBZRUf5g5+zcxifFbvJ7gcs/MpWzNRzHzn4b
WoghJVIloTrKNI4lAJ+qYXgK/vWkZAmHFtmyx+vRy4rNaEtoKqxqZkNt7DT2UEhP4mC60cIDJPPa
RhdE4zpOiHyKUNayyuJAAqOa41RweIdqiC/1Sy9Rk/lsIhpYwTG8RT/8EusIgE6JlvSNZI7hoQXq
3/cPFRImJhHwzennKqgKxLWv4rwHIeKlDrQMQPHhFAm7DDQPzseCMbhec3+RBrk6SpFczXYOq75G
3KBla3CtbtqtTe20S7Ly695P/XV4rFy7bCMMJTkhfyYu5iAxK8uTHpOUg3QcPnzhXrghV9TWV7Qj
XbVJTkvD/0FgM7a/BoVh308u/7OMYyenip5jgZV86ppXpu6xX59U//CcDkELv0pfPNLhbZxhevBg
N5ebkCcmAxZ9JJLKuUyH/44bk5RnQ673VSVocCdLsPFUQ9mx91Ct4lnQ8fMHFqnq7sJQLo324bc3
9V/P426yrkeR/eDX/hnECOBE6c4ia2mqDvjgLwWOPCChKdLBV0QiGgbpXq5a+R3N9I1ZHpkL1+2B
cNX6yGn7Um5AcQfDCmwfX5xGN0M2Ow/swXIj5myiUpKnhewPmFVhvKTwPm1qR6MuKFoR/RpbDMwj
7sXAcA9SQPznSu+BqDP4tmsLOjU+2ceS7E59S4wptt2k4v33I7R4uy+2ej4t4ayZkNqfu7CanoYA
CX9Dab3J7ll9BpfBmyxP5rRSozV66JFRZnQ5hbJMS0ey2okROK6CAB1u8qcULGL9Dq/AAY9aUQ1I
1c8oP3VBSuZg2XKe4VEGNYUzfheVX1AhsdEsppfLjA6jetnTkTLkz1gBWLMGTyV/m2Kk/hCYehDy
K8CgKj56dGrAQiYM5Dy5uLp/Or0Pq3f728lnR9SAYnqOC8JdOimdqys6SHKwUlJMLTJXUCdFySGc
BXvd1LzSxgYiYDMSe1A4yhMcOwMTmQKDdm8CFwllVKP9uZGdadtV4OpOjka5X+DM7F9EDFRLvmsN
bi21kgM5CSAFDyq6tdhWkVXSIU1oxtdN2fB9Dx7yy4NV2LwkWo+RfBi4YpF70SG9c+ZjAvHPei1l
X0vI2rKGRtkyES6j04fbpn0mHMSIwUa3uqUFMiEJ8rlNkDGhAG2qtu1sYgqH1c3n6VqBqXhQCbcl
5gX3LC9FvIrfyEDHZnPkxmlmr1/ruelm9I3lEWY4wk+B/CpNzweWKxWhrbL1j2yyA3YIAVqP96Ac
1YKmpv6tkXRRjfFc4C/JDXwNSm5gprIPpznPFL5+v7d+4D9zJ/teY3z18ToWACRhZM1J3EyantSB
izJ3nUCtB2LNOBoPf3wIvjVrYlPA+SU7GXOdm0eRFfssPCAta8AFI/hYNw6sQNJffr5Fa5FHdEBr
V61tYTOP/wGgHojdJITVWl8MtGJFmiDrl7q2QjPWe0ia8/yOSXzWp+1GWXZSkFjAhBAWEaS3Vhgn
VU4d81KyQ52yjSfTR8exOCtA7M+27fQJh4dMWwwuiaCjlu52f0gqICAGxPWL1gSbsdPcsfPmRt1r
vWf9MgElcNXepycTq1CpYtigQF6sQvp5hBoaYEjvD7ZsqrzYTzuqpjOHOzY/KjCkbtSG22sPKLLn
Wgsvhj+W9XfAt45ZD+lHNsuc2inX2wJkxg0UQ+h/A8WgvsJbwt41fj+bXqBtFvwBo6t6BBOXzKzk
dE1gruamam0rkRKUyREsciGwQqnFSv+QV/ingRKFOnjbHgsx57NBQpU1oYv6ZRWscY4M2GgOewo7
WG7CUAYK0mc+wmpTvWRUjaOG2jTkW1upA49rAoCgLNZ80BMRl+30M7l5ZnAQSYtF1k3/6OvimtTN
ZXVgx9+IaTt6uwXjP767rbPKbTEOs56MSOR71ucMLokSTLf3BHLQInq5gdKC7/ck42nhCa2Q6KxZ
LAWqRSZIX8ZV7O/iARfDkGfYognzrsM8bnun15Uj7b8rHEQmhY2rV74EI7kr8oosIESxOs81CcF9
m2RFh0MXN/UTYaFztwdF6cu2Wqo2eYpZdMS54U3NqE12ZDe/k6C36wPHDzCidv7ZxCcxnHFGizA7
UcTi58nsnI8n7xm3nqSXOwdd6iGT+YCm5/PTeHY4505RRQ5O7uJQHa2zh6H0kaEA+uGr3zaQdFJy
40Qs/IWlDYNfpe0PBnM/YDY1I41iRljn1K1dVa/kbNrYvZw8In6BVbzB1L20iWfZnu6Xv7nl5lBK
+N4V9tM558RD5YQ1B2L6UWcpC0/+Y5bxFv0mJJw+ElqC1N0xhzyTeNp+bizivGWOELrecAc8dFEK
mWvo6NK98UdEEz3cGzOhK1XcBKLp6TrDmXB/7Ef9Ca6CctNCvbwltXmg7zU5iqMqDy2alUZdbNUH
KvLBWQuaUMmj4Yx3SdHnlBp7mCH1Oban8sdjoHDwzKDIq1wm3iXfMrmMkpQtfehXhE40Wu4iwUgZ
ZpW90OHrX11B7b8zaLdrQLX4RCC3mx1Juow9Zq7J8yJJsAffRh21iPoksAAbfEhkOU0jBorAjLnX
QdPMvzle1d9zAwqPzXcqYUjY7Vu0HS2zIgiO5eU7c6C++84WTtuK0jKoSwCj3gX0mOfpEM1Br+yJ
JI4REOGSRPwuEF3+FYJ9iQsWkSqThgQOyJqXO66ATQvFqAQi+k6PKC0Yn5ICBkuB5/MjxgG/xSpW
aD2O0XbVM4IlTGRCvz0hKKLpGoHonZi6UlriDppgzG8o1cJ/z8nNhGD7Xn4l8Eg3+Q0+TtDq9viM
9Zp0ftQvFD/qOuKW1jN++vGvBFCW4U2Ns+lGT3P3Hgo0H5jRjq1MghUiUxbQH1kpt0dLytF12M8l
U2duDL4it6fKsxaeDdtOu265PwdJihkze/EC1quUq2Vp73+X1h1aKbI48nqiNdLvRf2XZJXd+qEV
LXylOoyP7h4s40rYQh6mFvSWP1vCSLbc8lW4Y+3wQJ45srZE3nnlm7X9sLepi12zxdomZOFjkNqZ
ymcSXhyNWG55akLtxdShfIWS32pKoOqBzAnYEiH+fKXlwjy5DPVMpKGaOjbmSxaWI18npq/NX14M
PrzTLNFyl5wLmeF8pprgDgGwbnpayYLNJ4D+D6vJG4ka6S/L+16M3PPb/Y/mvGQauQJNyTo/FYkx
okxiw6fm61fr4HqvZ+tZkPyJrHrJ/so8L2e2J4K0H+E6m/2jh1vRwrnJ505S33WVOKSqs7WrIJNE
dxOQjrBaJ8ZNQ2EjLM/MuUarlgfjfcVXLu/4GpqQSMOHUkR1H8d24SNEu2E2xcTDc8QDngaJpkLZ
KnrrJYSITQzS1ezsbRFZwFdb/f+ksHx3BVAk+ugSquUv1XKEF5iD/KKdksxSBqKzsrWbZRteRYyX
zw8lQFlyibGThoBfPaVYt7zEUoIhwpLy28PiY0iz+X/AvWEUYXI77G15IkG6+G/kkK5itQ5cBxNw
glcAgP1NEHf/6lhrQh61IPZPAT4sGyGo3LU3oekLOMxxudTVONbJvH5/WEM0JUUzzGtXjkU8Vg6i
57VrAsbkWXC0j01/YrSywNO/r59h+LxpBIrLqfPHR2mhVURZBMli7E4BzdYf3vege2aYVLwkBzsI
dBw1y4vOvoihzXbtxpiqE3MnNQayf+u7nqiPZPmVJGt1wtx7KXBOT2FUxLVZOYwgxqmWinBpFy7z
GfDPmFWXV6/pLP/+57u2oCpDOxyb11vkSma0DCfjBXFN7zYns0hKEzPvpCsFNLSQc/qpxXi+7dAu
Xe/qoZLE3k5rwTko36qn46J3m5bONPEBp+myuxSk8jWAWMr6uuM5J7DtxM7EpVfJgw4kBMPQQsOb
mgS5T23FcddICzn8MjfBWfen60BWsHF4xSSnrQXsjfU1TAJhCgtWILcBtN6ctNF4p/MSB2HkMs6v
AOjNEZ+pdENJ53ANV5k+AGH+ZMn9/eQ8qXsjzPC/g/ZJnzZQn7RyKb2qNj2WJAgkB5ju3Nz5Aiui
zWmug3AyimkDetpdcfAUGFrb6K+9Qo7mozxj39YGjHGrnlzm3GIuqR4ku7x6bxPs0YSMWV/cjAqV
GUjlIgSFOxymlImPXfr8WvCI7q+jcZ7RR+yee6j2NqK/xY6DbPG42saKWAadh8gPaUilIo5erOMw
ePz+aW06BVIjArJh25EhXQkOiHL2tRPjiSUkskA8VJmYBGxBvz2vZL6yHXMBcAh99h1jzAbNV+SU
wnSOHXrLqq2wBZ3L0orHST5OJQMSC1rHfc2B/iv0o7TWUc7J7nC9qIhTqaQnEGbxps7isaatYCtk
Lw2Bsnvj67nvdVLJ0WG//lnt99/SgX868+wnKaEMYWkCMenCvwZna9n6VnhxvAOlJUniyo0QOZTM
mig0DSDbsjgln5MWOJ2TBlyu9Kx8EVAbfarEPK+SuiieA6SRM4kJZUMvFBg3zBsUWtD62AWogYKk
YcMD3uurkJlO0E0xp+AjZRN6Z9QQEZtvqWXaUAcM0UtYjM0AUNkGSeqcSgivOF5O5ouur82Db2hT
hGXg/S9S0s9I91Nvf+SqDb/Zf1btF7LOvKPXRQfdIIEcrIgV0N2jXnbSE3QIfiw40Of10D/O56Q3
l1VCT3xbKVw/VHjR0Bd/9FSN6wcN00lhEIrLWHqM33oTaCNMi13QQSE7rb47JNPaFsxdb4Uoajek
yzzAgx4mOG6MB6VyVIUL0tlrHw2pbIg6VJLVRHsx8XTgMHs+2OnilX9x+s5xN7nyy45RusQ8R8eP
FyRm2mhhoo/+LHnjw2pvgVQEHnlf7NBkWNhWspd+rMebE24MnnA5xDbJUAiGvdWTZ4OzT7+yS8Nh
ip9OP+YswYqase2wE601/YFFarP9HuJhkOiRdOZnbwFooL9HSrf/Px2QJRYNlMNybgbNuV5vKUsN
AHPZi/NAz2LuBxf0XEILgxBShKFzefWMIEhS93KiMVpmN3V4RylLE6Mmdn06xdeNQsccTCxMUgs5
fGBX24kmml4wTTVG47kUYkmjLq6ahNr2eku3UqdI9pTcvOLp9C4kMAnx9ADaTt2v+3/on47t5ZP2
ECXS9iolWERGuckDeWmgfpJid5G84EA1wNNaWpeMtIU40AXI61yJe5y5mLtFXZY72bTtWCFwjtaw
d2dQ1u3CkK7xOZI8XG0m+4rrHeEJUqZTs4w9YbGPuFttvEo3s6Uo8PUQ+GoJkOwJSZjOtwMj5od/
+UTX7jvYGpx/TjsOVtDks/aLUpAEyiEUkUO3FpJpvwfyR5J7Qw+ZvVwjH0ebkZfrZDkxk688S9jB
SCPUHsVUQvuDR8FC6X388HQvK+LKae8gWeGKvVEbYbfs3noRbJwMsPot/uBXPQdoogY2RcGWTDxk
RPKhu+y/3+brNbOCulXLZK5aSMo9/ZtzAHumPO3qYyQ/5f26STZllwoIypuAP5lwy22GhOVkMhKF
gwq/oidVS3egnC/waHLDEYDkjK9VG6PhAIILOerhBlOIMGpGY34VRd8wOD44X35wGuZBN7y+OccG
6TpqdJPac2nGUPOO5r3QTqRne83uLrYAMkrsQFGlyyolYa96qtXb+spfpgaXj0HIi8+GXCa5TFEf
x7zxXOTm/WnjBsNOpAvL34HpW6e3xF6p5jpJ7/sTAPVd/sgW7gzyG3+oMGXJ4zNUjLhJ8OJ4llLA
rrYU6AE2uWpNKrd997zsbNSdPQpYWpjAROOOtNkjFNgkWSM6jw4QV8vahl1aYAfvqOjcMiRezJo3
XyTT5rQFWEgetxI8RRAVx4Kw90kBTuZ4aXG3A8CTZn0Wc4IMYPdfAihHO0UmaODBOGSG9eoYjtRF
rf9TOFSItE7izAfXxVQMtakiTpZ7qFLeTy0Jj4DGAR2m2iNnW+pHrLnl/Jpm2t749E3tBs97ZNnD
vhXwZMJCXehNDZbjxNHxSJoET6jrPUCmTz6aO2MnKfm+1gFnNGqWGeX/g0Tad+vGcEq/JOm+NGpV
hYatt6HShf4lACm7ZTopq7USniBuw8dr8OXprixKZ/trn1SiaLtjrY3NuiZPUdZ9XH07Y+XrGRgB
cF2UPpR3bmQ+mkR+tK7oDjCHCyqSIfDF3szq3s7wqoimRP/15dHlAMPS6eU2lptI/10mUFzrho3N
BNfTVBRuPdZgtuIrgGhYYgLH0UleJUbzBHqvvJelIGl3BRCQDWMT67ZXs06M/WG2+DE0oMYKt20Y
u4zkYZEJDbASQYpgSdnoVEocCaZWeQQB/jKioOVV/m/PUJtZbb1uIC7acp9UygV7Y+8ax/K/+GuF
HD1YNYmfM2Qj/RWFajXcQ0JHSsZlsRiYQE0ddAzduRqmEZzBb1S0KA7ipLyOlKQveYyBebJWQ2vW
RjXNNEZQ+yo8HWdPilxjWzP+tAhRbWB0AuEj83RiOZZP5pp4Q8hmR9+ika+UspuG9YIZtkHSTXVD
zhavTtCFzKQID2cHhCf+XmPiyE4OfNuY59NjkLp/Dk0TOXM/XeikdLlpvDqrFIQQ+Gf7JglsdRQ/
K4cnrSNjqeyaLDy4+BuM1usTvCSnJOkdFiBzfx9+2MOUWGFDyAD8YleLUGYQKlQekCj+3LnZERqk
PCcS1Sy2Pv/CgRvi8WNCkcMnZvWzDuDVV+4Lj+CtCh2xNSbMska/0w18LjkGBEuZdgBzmSmc22TQ
+JMxwjtANZV14Cca7Uns83gEqgnqcXtIkolpkZtAQnfarD9wJmIWpvwrziU3nLpAI7uALB2ZL1hG
KEZrczooZOGFLv7o22EA1I2/ki8D8deL57HIKY6fcv2m1M+zYOG/lmRRv7f0xy8TgKmuyRCJAJg2
iGOWkvSEYb+X6F10yZXCVYaKEeYJJj+ECnmuSO4zYoHuXMqTRMTuxKDJgqLEx3L9s3DPPPgqXmai
dDSkc3L3riTkWtgDwGw5X4HC1qN//WTbUH3BfrPC8vl1hTP1d+DGjzJFn8niinG0IIUsw+iJq4wf
qvyih/VDo9u22Mt0adJDXEQuc/d1d4VNhKngDkdVwg0/4V2d7s8QmNe2fxY2ENq4bsx8nR3RvyqN
wtgHWovgVzm0Bg2Z7DgDBG4lgkQmwjgznPtmK7yx4sDH7K3jAVVyNSOMGQJ6WGkuVv6YizTsrzmu
EFcZmpr6mUurr0nmwzv0oGjTd6HLZ5AHyJj8rIxhCqCnktcxIdNR+ub+9LDW1Ykfhl+RPfWsVRFK
Owldt6iunVfwh2FWD//8i7DplQhkpHi9d/5deNpeLRRKqg+Y9hbH4OFALqb3nvEcYOsKYn2t1DUR
0Xz/m/Lh/EggdZvUFyil1rG95ah9IxrlIQUv+JL5pi7X/ILe6UwwUTabPuuskgn0u8U20RTe/+Eh
qpyEzpaA+loJPSS+rG5mogj3c2Bl4FoxMhzdVoFnPWx0+gDcsZkKyPI3TYBgddJgg7dBZ+PO2IrF
ndK45AaNJxWtvlirR3t59hLluKjOmf5UXGjHWBRpSbE2zuMrT2MjS67HwVKBKa+y3Of2RSv1sZoZ
7HMtfzaStzEbpvFeUFYd8WXeU8QJTHOmyhxzBF7JmjrVEnXqdfd+jJ3CWWHxYUeoX99KJDvRxX5z
AO6CTDSh1FKNKejIr3QmApXG5mNby1pchCv31okHMnTBf2hYeMjkwGbGMlecj5iuG3va/Dyupwbs
BJen0k4NFX24UtcQiVwH3pb2s4yw0wuMcLcm9DOb6T+mn2F8Msys6gf45xTF/y4vD/afaM+rwF/H
dmgr0Hr5sJVF6KoKYm2gACIJ7G8hhJA5pcUvqlWn1Amu9ZQ3WgMirMumI27UuLl6eslg7G0eBos7
OU+1j+bXCc1B5Fh2HB1rofCFxX75OLi+fyMOjyc8Hlzyx4qRfD7R1WvDokh438zgFsHIzeMulgBF
j/JRWjNmp1MJZbUts529X/Gv6HUeolN43xidfZhP4sbizD1JSyu9ZqQlX8SPlre3G8obGJzl7UTv
bTHgtX3oF86Ux07lNDX+mSqsLuhr9zStJoBexJZJCt0LOaTQdbaDOulwcbWP7B/kVxlVQYewLhi2
dIANlTTGzJD20elo/wUWkqGYtnAGDNqXqKo+lyInyXSV5eRMvaKSRnJjZ2lK9bIaF59SSFHZG8ix
XZB2rYkbjI//ZnmA45SSzsaU+MWu0BHabO6PJbvmhVvda/zOCYNBkFecelKhpCjwA24gKRW3SwGO
6V7LDbhdL6Tz/jRUNBq9LLFFu1yhEB7u6hIhhGO8876terf+IQlFxzQPFSKriAAagOJONTpGOwIr
cpOZvhc5FULGUGl9oiQk4tXQUPcMKGWsYC0nAirTaoMm7I3WthLWEbKs0ZAEc1DQwIFpGP3LeWMi
8H5Vu5qIdMieYSPV2nYF3mc5eNM9aiqEfXDnNHYar73VPGHKs5JB6MPD6UrTR12bn7+IM+rMfXgM
RdHpe2ytLPGQLohvIPKB7H55kmW4MLz+cFI+kj6cS4yALM5f6CQUx2S2K/Lnf7L79k+uSUo5lRbl
p7i4f7JqTN9hgtS+Vq5SVScxVV4ictXzxLmWGNj5rY17mUEulHSDka44RvfTD45Z2H+IGoDmxuXM
v/Bq5x5TbQzYdV0wdmJo2O0qr7O1Vnb8t6/GyC+S/dcwciw/cWiL+a+uqn9OkMpHjv58eaNJg2SU
xiO/s5+iodHaaslPG1WPqACf2Eg6JQkHvgweZ++QaMOaD40704lBuzzCZABnlT4MbTwL72YjWGgL
3W/k7Fjezwo9wZtDwgxEMU+5B6VfdDhm5pMRYpVpAFD534XEswMLqmrtnNg/YzA1+TlTao2XM2nB
iycLX7fA9v2UvDZM97LLoMjvaItWxuzeJfh3hLEiEYs9SQ8d9n2kf6v1My1O8I61lhkuDEHMhBrJ
7nbLJFkKdxHi+ihlnRq3mr/iQqLfPuE+MRErZoUEImGScAkfK8ZgRuRW1wuFOfu0DGq3Qnpl8Q+J
fNbNY6CIXxDwvVyLR9NHlfHlQN2y3RZfjNcY//KIFQGtcbHd8UfhIIqhpNyCiVY6u5UrNWpYSMqn
r8YmG5kstOEyVG1wmy9foiscCcRJWQtvk9TgsWnYREIK6sq9GMP0khZQuf6apXVIjAWBqJq1n4X2
tKTb7Cba8lsGnmRQH0oIT0O2CLO34b0YhWGvcRilZfXUflBvy8HsQTHLoKy7XvasMShfnloTp1pa
mf8Ns2FHh0DdQYEgChyrjmrSUgdVAFEPGdIEl3lE/op01K588LBOg0nr1tuSm6vd+RKF40PL/2bi
VeruT1tIfxfteLvDuKSfpORHeEPjQDU0nx7B2FxhT6WAneCrTsgOamo0Uic8y5jo9Op9c0EG1g/P
XuC2WZcNkHcnehkxLfcOzd9sk+MIFHPIjrSLMvvx/+DIK2lHvXoQkPUlJT5N/njgj6/RlWhnwJLq
AuS3FdueaL7cpUzal69x6eebzW5B1AcGvBxVTvOBIPth1eYwAOWUb5++yDZ/lo3HDWShMDXIGhas
MSWUpxb9Guptp9nBESDKveMUsNcHvF2njAQZwK/1RHjg1OHk1Wi4WJzxS5J3jYguhemYOBQ64GAN
JQ0fM8qIKE+dt0GF7UqDvGIC3DZ+zk9oLe2ypnwT4qPh5qhmNsZtAjOyrCReV2lF5ZXt/xl+4hoo
4oEvQfW8Y4WwHhOK1MG6lxRL8OO/nGirIFKS9OrsOqin6/ctoP1p2R1Tm+wuekTR4c/qLIbjhs6o
UfBS9YgkX/UxGU6mpHZ49VkqTl94U3rawigOsgZmLDQXBriGBsG+xCSuz3PTVlQJ0FcGQYkFWiAZ
zaUY8vWTYkCU7r1pmxd9auJwTyTakHi60VE+Sy8pri7jkQxVRBYlFgg91o3ahcVuADQs7Gf78VEb
LnBP9UYcjuxhoEw5HTudyx3vnxrUn6GxHqLvt8tEtqF6FveCGKVSwu5xcLOGiizmJMCRUxa96yzT
/kFYpoyPwWbWpIkfud9L9VLNaHkiAlXu+YsGwd0AZa10YoCXt9G5d5UbaXk7k/WDUpKCCHJ5fDBx
0lKrH5dKvRQeVcqr/TOPcBj8KSKzfes4fjy7IVti2A30IJgLb90qsejI/Sob6Tu/FoYhXcCWCEkk
qipAkUc2YW/uTJAzZR7HKbfn97XYvNtoDojO0paVXQudvqm1qcBiIHrZ1ggQ47zUqDO5dbEAHDAg
UrThRcufjUGDtclil4yQeqrinjutDGovndM0kVtG3i98Eeklt5SbszpdOiev52QiRW0P+9gAayDu
1hOQLQG2rW5kIFa55Ur9ZvFLSgvZXATk1x3Vm1JBBxSdz1DgOpE6ZNZyYS/fbvADIEjl1T5XRmi/
RCKtBZqvj/+8Z+6rwiz5Ph1j4AbpBjpK0J0SsDUUgi+luhUqt44LWiXNsW7hpNoUacyc93SK15e2
CIIanESosFAa7XJAJ6ZhHcFx0opL9AVU8+mlXa31UB5vNwD1nAnyf8uQvCxt3H5e8d6SEkQacXBK
6xfuaIcb8b5ticLdNL+KSNt9+Q/uEOqRFtEyKYjQ6EKBYPafyHN9CiCsP3+mWHepCe4aV9+cAbkC
Yd9Jwm/TEUZ1kykEcPazlTTmyKPqIcJo6fjEWxRS8zmh/MjMA7o3VCsu1k0aIqLGu6knbt7t4/f/
7Dickh6pcUvc/xYzQpK5W1YCsT5A2a5Nj5fKWJWA39PdQi0gvsaChRHiIFNmQb29Ic7qDcOsYsKg
ujGraPE4XT/mExT6Mejhz6lC9ay83v5NONNuQMxuxVN4RXHlmwIuHW/U+YNp36LlYINcbl8w4HMn
UkClEv5H/UfxOppaeQlYOER+LXOWyyJ2JEOxKScC1iWkNRDABYDRH2cEhYh5L3tVpWM+E6WLdGXO
Q3Rgt4QpcEFqOKTd7uEQG4ij15X/GBwJQs/EJOXHBK2C7JvorJCYFofI32f14xS7abk60Ql8nt8Y
8a8ZqrHimw/IXC626bj9Vjl1JRKgvv6CG5evtZoTpb67NGuaXUbER/rqS1ktKjF2e27br8DljzYo
+/LNqxyXDDqfw2uTp+o87ylq9ZuNpdICGhqRo3D7U4V3AqAgImN4ILuj7i+szprmG425mpiA/lMA
lP1UKVX3JbJqqSnBBOhjTmw8R9Y9EOLF4IGiOSGZ1Ju1S5+r529iOWVc6+G3cTM+LMsS+JDrJeSS
hCtulSmnN3Ub/voJgZnaYzvQn59iEaFIo9UfIlyJ4wLU4x/RKvsmQChnIGYm13cXLLTZDNOlC1HW
2aGfD25bkjcfgaISfUpD0Q7JqG9jdP7rOhOAv1p15VcP/ZQ/L5dar+gpbkyNfanfsIL9iRA1dVTW
mwEhm6RAswwImRiyVYuh0LeLAb7qKpGXKA6bo3yuKWbPUIy9H3fZkv6N1vl0zGbJzViTEf3B9WfY
mnMLrWSot5scAeLJmKgXwIri7wjuQEzP4j1cyR/DtFw/JjhzmfuVn9fW+DwTlyjSU6bBT06RKvSz
yqyLAS8uMoYxjAnHkthUYR2UhJzJ0qFBKY8B1z6FAessvjvQphSjeEdNwYRn8Ajuq57JYo4M28ru
mggvNK87p54tZqWqU0SYMbrASxf1WRbViexRlpAync7XP5jJxykeU4OtL95lIzEhKawnND8PUkC4
u2RB9FR5WS3w2BaSngZsMe6Pbtm8ARtk0ZlOJY/yRVHwUxCWACrAAMgeViY78MHJZQFW6FmKdt5d
tbzCzW2CRVm+T0V9DpMrRb+CJYNabPatkUwRFwsMcZVIkoq1Q0Hp6LFwaUaUMJ+wg52hyW/kyPuq
XHinbGwKifP+XK+/y4OM3uL+w4Bc5RnfKmX/yvOkwhWV9IhfcmjS5f8Ir672gRYmn7Nm6Ij1O3V8
pRHjIdjqENvXBdDlrB3oYUInky3nhZJIf35VYjo3bmYN5wssRhY7Y1dA4bNDJgTQ1B+1z/r0oWqM
ooWuTKf31aAyRTLOap2A8KfY7WafKvfzCK4SgPFDJD9UlIU0h8hjteXYpyGsz6nZXEVW1RduEDv6
juAezrIxFoQVTNxTsrrK+x330Ml1vG708OzoTgWqI5o+1/zrSSAujmKoeenP1XoQ++A0PHFDIoZb
v+8PbUvG6ILdjmiSUuoJ1wRUIu1YiRHdq8DB5XR/7/YMpKTM5mf0BsIKwtrVVsfIfl7X2O5SRb6T
NgWKmYXDKtaqv361UpgR8sCQXeyCMny6KcJN2mxs7Z0eYvakINyT33+icKJF13kqB1D0d8kmjS+X
2hmSKmvT9Hz8bfLZIJsXh7W26vQGaDjVv/d1LX3uX9HvdzwYNEAm6v4s3U8HJ0PJm3Z+v+QrJYbb
bu9AvuuSOoxrFZteCeQR6YOwTv7ggii1PL44/MZ9WCD2lPGlBwJShFQpQln/0rpFhnKRsbvMEC4/
tT8SzYFc4mHXwrY5uiY2vEmjdWZDrzF9yrU9ztNMjAF62i9IRFza1yAVNabgVGrLAutLuZsA5XGx
YR6Z+9rrZN60ukPkSGCq5u4ORsCHFvCzOSz6x454rIg4EXLuT9frBKTWuVzpjdprWAxullUzRryB
/rNAcVgqKDs5M2GxczaUE2HgQI78SX41dv1/yVt5oiK637mh6ViklbY9BfAnPIl2QKIgs3SAbTFD
58ZDv1Q5jXYubkP6zr/D9p/Z7fDWMS9i113ESOVGCowc/qSipPbuW6z/JqJpbHz5LYEqipLm+CY2
Q1PrGn2hAf3J9P+aCCNH8ihqrbgZIa6Jhwx50cNbtwiSgB3Muc4eey+e7QQpZXHwzCuUVrbRaibX
EC9DFTE6+66jcPVrfr40/lWXrZgimOt3TvTCKWjIe+W9Wks7gYhoFgKWPvR9rtW66LZaXrALrFE/
FrufA5cKhMM0kT5s5jW+IZ/UZynpjH2zVdO4MEEdreULrxfhsqUrCE8q+BbXiiVsyi2F/zpjptrS
U+PYYkiO42P0FqCU5NIa/fmU7K8nsh0jmdJ3X0oyQ0yGE9chq6G+kkZal2x4qTcDNMXYfprRvbcY
lC/jp5pWOb9jKR7+a3G5OnhyssEGKzx5MutH7GYPHidkj0kvmmgkCBKVBFxlV2rbirxcdhrPs/mp
LzxWxCFsRiJHROYWjrVEc72PnGdYyLwzJQEW/Ac+HLL6vXDBqBB/G1KZRmCap5vavRRhkEDB8/nk
N4+Jni0sG5M5/z0bbcsb6SZjU1v4Q8yhTNCjuBmt12HNUB+YdtHMh0WF1PME6T/0jr4rpaG5AYlV
4v0O/8Q4MKCpek0SrQZzP6VyzU34E2td2JYHUU9ac+RLTDtCtmjA1t65WpUh8WGxUMslPiqZu1UU
lVUBeuMeJUZzl2XiMMNviueL+QBioUYeVYDwoVLCip84YDh6tGAbwm7pcgRp0eYyKRxIUwet3UDg
BtxTHch9jHXeLmg4WkjVncM/FTdS8+TcEC/V/0VJ25tyv4xFYIYArjCpdsvKiavTS34mtivJUS7e
bbciAwdXhSQ0hUWlkDZ20BTDe3cvCnZ/xJMbyyP/dHUv/DlnFOq+Qk54gJfvzwClX5j/696aSuh3
QXhIU18b2p2I5bdTj0c1GQR40+4yL6Q6HU1jVlF6vbl/Ntxr8OLIq68Xp3LCDtYaKr2qTxH20ynq
Jz1+be6JIXwopCZiHnksY3vP5aiUjyAFzX4jUuLS0yS0w89urBexpWaVZyS+71nES50x4q3ZETcF
E6P66sb5vJMeLp1MycmlwXA0d67l0sMLi5mV2HFgdSnH6W4KyEPKULXrHbI7V5tOP/Ag9+DfxwPQ
R8QHmbrn9956vNO9az0FmgztGfAqYZK0mCB6NFcTGnymJ0akqdFQ0tWGAnAzuk/81n9s3Wm53xFX
JoxGguGNs9q73id+nb50Q676lF/CO11X2tQTti7U/rxAUBeK5Ks+W3TdH+qVW9JUP1BX7MJUZA3U
g+AAhNEtZyPco/o/q3XCI6RonFPzzDJ35pbUsyzK0Vbj3k9rJb7NltUFiLdThXbFFUCgWXemgqKY
B3I5xE2XQgd8f9LSzSKc9J3Npk+kYuJ1guYoJHy13SYQPMD0PJJDtYeM53p4so+r8OHdsCJFqDDN
LXGdVdznDQ+9DdijFUuCwcduoJanp5BalsWXWYJzaYxrGlM9GCZ1H8HNV3UjMjXw9b4wteWBpg3a
NAutnQ8xa6V4O4cLyDe2/YNOxL7K1bZjJRaKeGPJAMsBSlASOeO1XdGzQLA1XpJ1gdYQBVxkzwpN
P6cDI3HQa9wi/E59osoOAH0KHcE5HO2QhSSVxPQHo2LunbGi7MChEJsHuGzI9dsdGsNOooJOAf5W
xr6skcZGB30kypfj9JkdebTOK+2ox1yive/afK/yT4KKE+4fYzdQwObk5WOuAUgCyc+vHAp4z4jL
ijgTyyhAK4FWdPWqbmjhoeM6NcI/XXQcDuqulT9cF33gfbbwuwQHJTer+antAYZT1QylrdQr3bNN
YlbEdQgrJkAA0Uc9doVjnqVAGz+KGdfH1SauJIMnJKQt3mMQrgDtNcZIZ79HKMb1AJYPHMAtQbFX
1y6DclUlpTnvfx0JG6qYeK2HV6PvPJMzcxjZa0tV/EilR22CyhZ5kRSCJxt7yOShgBTo+s4JdZ4a
0Beg1lkMh22K9CVvkH98Xuhgl0PClzPYPgRHIEjPbyMMYRr0tgYUFwgIhkX6Sw0mIfvAjQUFnkfd
2mRTvPR9uePmyXCe3T73/AEFDjw08DmAjr3JMoL0neZ1qbgIpkuB+ErtDzxUx+R20lL48Ci2Knz1
MUYYyvR/c/UBaw56ljyuN+dWaCBOvWQwutPwYedps/MV6L3yEaYSZUgDEh1ymdAAaom7KF7RAl41
1SXkfKqRToJh6IrSnMqU9Hui81hIUPTcbXXelD77eagCGUwUUvISdt6N5+FQzTXWMmSLEhyb879A
oPAdjAUTsnYRQV0Azhny6GNURRvS3y4PM8HbyqJiRKvPd8MpUPDEthCR5y8P2DtuIqK6gj8LOL1j
gRuFQwdjIRvkGMdQRdW7EWXRL9B3D5yBaBovitxaODL6rPa6/kQ4GB5d0Hs7UeyHVaP+jiRvBx+3
EQPtv1p/VRhH6IiZ926wFXk3xZcMaIL+IswYP27vfUxsNuSBNSVmxzsFtGEEPDSTm2J8dHbMdi6Y
8VzeVaFbICLrAsBPDTquVQK0VfkjKdx5aCKVDd6wqBOf0O7EiKWbW5wgDnn+5cIo0U878Cc+6eMA
gF7rIK6GeZvxH8TdEX2/4Dsb78sOv1RF4IY3wu6nQygo00fKa9rtT8rEScTWOq1h4XxIa53Zt5u8
UmBvnWGSZyeyenVrCm7DMBtnuD6GoGWnFEfETQyQkKOfZ4y7xUQSfB1lpTJnJwx9BrxNav8NQ2MI
Krm+uAj58Rlio5S4IqAd6TsuQzXLFvdNGeUW+GYNIL+94NV7RwC3jUGilRuu9aTi1RHljTtEq/j8
bEEl71Q0y24td/YeodZAfkpOHqd4/JTzfq6FW3Wms+huE+cJlXF3ZiwDlWzsU88UvJ4W21E3btfg
TNhFRE+ApchTJvEiCTtQCtTFlJoRvxnRRX0IorzS53n7wgy/XLd7POJaohW1AaxI5/53PcCxODwT
nVRCZvkvJIIyO/U0J76MAOQR9lhcqrtnJgpT8hB7ZLIPxJw7w0VKQmUaZF1klV6yZca1xTOmYOaU
OxHRDZ8rw1+jxTjy2ZavdF9McvN78ktC4Awn1TcYq9xCSZAIzyt55cujZOPHxxhoymDkPnAV6ViQ
J/p94r5gMl92Hqo9j6U7sCCPeZXLaj8xthoaMA0nJ51vx3bZu2VmedKthC/PxZ/eodDJDu+ZrkCJ
fBMEujf2XlkjlNIKn8lYAAzLgpe+XCAC9D/DXEO5t5p2iw38lTpkzc/gRR7bOk1LSTTMhvcOd8B+
qkBOJrylGnPMh5VyrV0phK/jMVlPyx/pBOWbMUXurA3L2yrEUHBLxP0HFZ6YbW+rLUf/ne3W1i6v
FWMBWwzw+fkSWU9NUHXSH5taFra/2EGtb7+mADSl3z7F8W4Oy5xYVtT0ypvM3R08Rhy41KFYs1/z
nKAFiQDe4P5nd1SIuon2BGqB8sEC8ta1QEjWtmudbmB/gTEC9mpsDTh1bceafilFkX5ijWTSA5TG
MAJqIgM7DQbJIb37tNN+0HHYCp9LizQdAOkQvTSwQQFue1Rz9pVZOMysvEpHXtTkc/FIk+12T2rZ
AqCmNMkdYY2mbEUIdjoFUurN8c6TJKblcGOMlgZZlufEdebbR2XAzTJIKKmYt+E6PHmc39dTGSXi
nbMOGmuxxmBdpKmRQxxjnSoMO7MVfBro2kZ2wipzo9AxHhALKOokuvsfAh2DenOOTJuqNvm7EGiq
5RMyMU//6oKqsIVasx/GjQzlA4sl3WsVbFb2IKQZVU1tCVx7cBZZRozpnvnPt4XFzRRCGPGNnXvN
bOOjHoY1hJM4xEhA+YJQBDXWrnBdeFDRkyKzg+Qx8c/wM2fK5Z+XxJTRi5CMkPNJCb79p/X4v4+o
7WOPy0QwlMPSkx+MNskQj4ow15YjQiz+yHi8DWW4+NiwmbEx8GwuUk5ogr9UXuOA3vAJkza0rsYI
6YeILmMFLviQ2CRUvVcoyDqvxc8/gn5VcKSH3EIujBg7s/kQlvnWovG22NBkpAVRu+pESHPujZVB
V8Pl39P1/HTJlZBzlnPoL5Vi+WdNBS9uLG/GfXLJXN7EY+Z4X/M3guchbb3NRWNzZBK5SqDKUfLR
JEcI75dNMxP9qxag+dXCnSt4+o+Gj3MEjlS1MEcRAJl21LAGaS9uJkVyDHlfZ8jDKkEYpSitgHPe
TN+7p0O2jNhqJP8d4/9od8CLP2WxcBfXfZgzldfcEe+4zWrvz8xsG8mI2R661TWqn7CV6mYtUIxk
J++qtESXVYjgPoa6uq+ey98ofJTvVANKMJ2xE7HKcnBqtTPwaZoUyi1M1flFxkHloxD0PLfMB+3M
HwaGlhGxpOCuGKl7XMfIQx4Fh11K3AZycUiCTfT4zzsPm5BE3S1mrX9tU26g8sbRxOWwGg4FzD19
x58ZoX2zhz+PS7Tn5BVTrJXRG3My4URMIGE4acYxK78MHPTXU0jqfMCMHWLkU2DZBjKyQA/xcdvH
q9S1egNQkYdL/M+d/4TCRnle7SwoWuuI5dtLFHyDticS83fsr05Gx7hKMgW4xHWtHkG1c6VzKfOA
YhzYjk6kf3cg/uKT07WnBQe6U0pTaiXi1lmWF53C+fxtbcLD5ftqTVkmB1NbWaotBHBjUZKlEFdO
XaSwCxucxWRNQWggG9nucg/UBdrJBX70ZPJ6SaKNXxoBVErt4veTrItiDA56+iucym5y16Dh3BeK
eNJ0ioIxLh1xy6b7iFXsLiTgMAThBFOVpUJSm+9BswgPXcRxNptElNb9h37skLCcXu+oy6Wt23Pn
Z2ppQQaBjC/rsASNuJYWoYltCpiCBAE92LvUvwUh1sGYlB9GVzRMxAGJTmxaKBY1dJdy9QZZ9P/n
AXM8eSnZ74iKBuhBiP75+9z9bjZSIjnOBvGtOSCFWdkMQGi4s1rLxfyY+REjmVoL2wCB3T4GzKBC
FrXnWzjwa68dtWkGz7PvI5ONEBZ/9qSSzup2DJuJQlUh3XRM9CfiuR/rsaCHjKLjfv6UoAK54waJ
IPATSS/Py/k1Gy60nUN0iCk9gNLDb6EYSNbh4ttCiKVGHp9GA3tFjwYoDGhjf8lu+Av2+zbusK9S
krulKoDLd7K7Ib6HDNoZ0YSUvrjglVdJEtRGsev9ibWjGgmg3bh1zMQM/18YEQfkmKD8lERXhXR7
fP9TQYxEzjBBm+xuY5r/00pKZulLV9hfdUDEpb7oq8q/s8yYZMwdnVlOnhuIh2DGr9jQb3TnKA29
GAhNcUPiD/02xm9t+cbh1q6mMXNCH3+QDd7H2zRqwlJQ1eCeBXHOmUkzj+E3LF4nc1kbI+ULifEs
r0lOz4SPMy6ZCNqnv0hWdmYbNny4AkPEvRGb9+Jh5sV96KEdOxRqrc7bua2fcQkL+dTIznBo8aiG
cMbRBXqiKNcGZZ72gofQv8X7nikqBb3lhA1cNPaO57b5Xwaj6/pKagjFDcBpXnd5U5t9tIA+qTc2
+d/2XsVs1cLQeMZDNu4VXnMkTRmsc2nLGHdf+o7FJjGFYPtvtcuCPdSvLWbNho5AIC7ul4CwFZdX
RhnDeBvha3H6sZu7Wg2bQY2KpXdRpU2/743m0fhzl6CWq15buJWdxxTINd2c2vzIU2Niaj7ANIFj
6Cfdh6H8o318HFAFBkuV9nxZBSKyRWFU8lI3RcqFaFUwyQkieq8qBIn290+YgLGYE1AgZra/t40v
Twf33BaVc/f8La+IhxXpwsOmdFfiCmeLSkJWV0EnQYMpTOmPmDWYaEFHzXwwTT+wDA24K3QoVbaX
284gAMWPFLLmBR3j/BDZ4RQvbVIj70tkcHikQA6afgbG+b2drW8d8z0fa4hd9D9FSeJjMkqB6uir
mO3epbEvrcMnnXbOH2eWMDauN7gYkCABE9yJQXs9V10TYA07yud0I3hZc4IHdRpENG9CX8DZpvZx
9vqEXt2ayS4HOtVCXqb4VTMWekSQvbneQuJ/TzxeFTFp57O+CIwpFdIZPMTFeQaEAKuXDTRIJeoE
81LADrwm56kb/qgDAFM0eyCAxjkm+k0M1z6jooUH7e5BgRZWit3ckjL8ZDrwANFzYDGWGe1RKBke
Di/CVSzBPzeocGxpu3SiTLsHdtddADiFO21EDMbThz3hiyMBARzHlzYJVsQ+QJurmOBrkM1K7yu6
u8W6+HN3nGBYCArNxgyDy0E/PgJLY60d12oIp40j683737H1kgg9o5s5hSH8DJkng3DVp4Y6552P
uaDvaLjbPnYRJpXvsysyCZqLA5tM6jb5rJF1xrkyXMP7YUAdW//H3CwmIaTd5lUDZsC6+FIGFbCf
ce/y23Ioc/6o7uNAZABDs/1A+ZqDuVnUmTbMjM8T4qPMTQdVfbeVL4OYbKxsaa2NZRHnphhZwLo1
0utxO+MBERKMCmGp8wykyPqBg+XqDBCU1xYCDc0kTrucL0zOf/Z4kj0In9tYXZM+lzK6FkTTAPL1
WSPtAT4awxYHh9btG9RutqwXpl7BJUvFgSOIk/816vPbPLX/Hfp9Lp5XcqCfdfQOhIg47Ao2A+2A
Rk9gXvJItILyWhZCh3SxZ0kvdEUVuWEhVEFA5MP1dS7R3H+BXjzzM53x8rBY1xNgwQOgDVySvVI1
k6J35UJ//12nTxFBNF7pDVNBz3Ft3mB7ic0aOBZXpmpcQEbR2P/cpNVHgBY9OnczG6Y6UqtRypsp
9pO2zZEOn2W24kb1uNXKnx7P4yt4rq9VRriMb0LJ7NcpNa53KYGOya6r/S299I5d3rWe01DTVsZN
i2hI15lsE05C06FzCAcYeG5s8uZ4pnyxja1oCJR2EtxjpMA50+tCNiUslzytukRX/7bsLeAguYk+
PaUMy8tsuYqbCgA7qKmdK4CLH5p+kxM49PbIabqtrpOv0+D3Db4ME44nq3DXcZ9cuunsGk+AoEMW
+JzTKaTWoB3hPVwB0BWcqmFzxNLl6/O8pa9rvcWR6qkBikkO7hD9anCgh+d30XlqsjsaHFJq20w6
A4B0BR5wrYF1oNI8RmGeMYt0iDBnQi2ff1/ou12qOVMBdc1rH7dPy6buQySTTYpyjXZmi6NGHfxK
SqvYBwimDKHenqQ1e/K8VeZB0O3IIf44LcXlC8pZjBwH1CpVG4vXbxm6c21m0pYEIHxbmXl+g47n
wraSRRcMx9WhmlcgmJmACBNkAxVDdS+JVXO0XSxfdxFi4nWkWq2jDSNYeB/yH8YQxPfe0k+DAJzh
llwx7cjuqN6DaZNxGX3FPGcbAYCe19dZaomm+YdG29QWI56ksHJkpz5N7Z0sDIliYECL3VnZLOfL
sD35B8vxHJfY8YPMM607JUIkKTY0UtDV8/EcDF2Y5i2RsPJc230l5viF8knelyI+iQnNdTnCCcSc
xlBCV8RaHf1Zgu6yTMWdjsRghsU0v1mqeG2LoQZJdZCbEBbpXxG4KklkesncLK8OfvbTfLjLCqLd
ttd9jgiUysiWCMyMpmnKkJJsvOvBwSGiK+x7SijfZHF+UcKvnIKK7qxc1dUegG4m3YHNW7kbBgMe
uCwAlx7xjfAZ6FreYfkf8nhYN/cQB7FioXRk4u5M/gxfZFe4Z423Mu/zThyDj44BKeXfnxjcv5j6
JFOhcUhXmLM356vS/aHuqXYhmWK+pjd3n/VCt70/bd0PscRhA3MqYPKD7w+Z28LVvYYB98/L2vT/
Q42SNkMPXxO9m8bLGOWDXfy84e7Xr4r5V3AV0oUgI66320A+H5T7yaLSgc7w86GjvgK07wbN9rX4
oYuFGlCRS6WRF3XHRlCFfSX0vNRXokUfUgjOs5z2tS+zCjTgSEB3znMavarQBJm51ZFgRf4URmBf
FpWrk3b6tIHCmmP04SaGZBLRJidJQWmXlTLO2qq2gVJVjlNLnxmxiAgfcP7twPbCI0+KSejxWr5E
jccSHVyYyyJJvsMX2FLCkMBHzdgFmeVuOTdLI6x6fNbL4z62dc1fO7yEZIWjl6M1XLkhxC6DkMPt
OYtMOKl/1e3pkIPIIjC4wu10sE7BCu5HC+3TWVBEPMS8ZqcuSZGI8FXt//y3vp/hFa+iI0Mfcbz5
pPvUMCqvDTAq8dDL7VBNPXCHN3MHu3U2eP4Njd/ZtJzIEEXvZ/pjWfGfxUKJxw5geOXAgka1NQqJ
CxNxpDnM44qiifyW+TMAQMNceHfDXX745O2AU4dmekaaE8eOfVy6rCFYXNhTUAq8Bsi0ayRDLE5B
c4o9TiakLQPP10ZlqCUYdyGurz8SxA0CZ41Ml549lpscJnblRcfOLNGBpCS4JRfM2ZCYV3zQ+33K
1uv9ltHldPT6oYirWRIhLhv/KfiHa0IoYg0Xve/YqfVv2JqNeKnGJ2dJNeX3HE4uHbDriFn5s9UH
Cfo37sNGhEc/gyd1qMK7CYCSDbm6I562B9Duco5/zzZYDig6FJazIcDhGEgib3x8x0yyYqXSR0Bd
Sa32qlqJUlfjgGYJC73jb4nwmC+uF1S8aPVetPVJHTmp2wzJciFyGE4aVYwU07OqMOdkAv0MdU0q
MV2y7DWGZf8Np4fq/3V6sYeKeBOTn2/zi8Rj/ZHRhDrfXRYAUuuT8WiXFDCsDSPZckDP05mNlLyB
5Tr63T2GIB34KQfJfGN5OpmwHFsxNisBwGvuMEO+b4WIzOgyPO/OE7ejpjNOa1V7oULtpHpY+ZgG
TDOgKOM4x3xz2C7mYO2ug7Dvy8E59htDd1N0gOetvprNl05JAF4vH5qGckI2bYPJD23N0UxwGe5d
n2oDkrZGu2uoTyGx6+K9k0BK6kzToRN1aYjWo9B+nCx1bX4CIeef+ftfEAISmEbgFHQPb9Y1fnb6
lSJ9ctdycKT6QnZ1wHxJ/X7TfMHVPokpN3GxE+3DqpaPYKuC/aSrTl+Dju0Dz90Q72uU6RzlOB1f
TddVazPN2FsspAsGgsUAmnh/6tC/fuQcZgqOjQg8/9iEq3VefDi2kj7xiJUX5TvFivwW8xsyffno
lY9Uy8qoroQ0hg3TUKGp/vIq3qUekEJf+7nElZfJlUU3uSXGZda+ivY/WIh8HNBuIC12B+6Fd49D
awzJzOStiF16n6H+HYRdB+2b7PYP//gCHFokfbOHtKfzbh5jihea7vEvkVsOP78lvxvKUSHwFMuk
Nv8gtk1QyNycnflciolpihXvL19MySd1vlZJPrEz25gKl8Phqq0sfHFfpUyIVx8uZPSsZ/ueShHF
4D/3oPTCW2F2fB3H59AsQJl3y//uS+e9QP7lkXU+xjoJjGwSOkRWD25iNDhLChvIwDuVK1WxM2ho
PiLJk9YkuUyjH0qLYme/PpwkARR/QusG/L+uc0iraRfeX9ay7HOiKt39bwmF4jHUeuVs7Ki9NP/z
dQmUJPmNn2WiXB0/C0bd1Gc+C5OAZ8zP+b6WDYOdFFyIttY4DyBHLyDjNvYFbaRFJiWUfeJLuJlM
ve+dmGwJkqpIk2o0qMR7wYuatCTk/h6ciHhEzmbUWANOAF9EJcrqfsGxCnpPzM+mNnEZAKKshCVf
fYMunu6doVdH35zrlKAJrBIcJT15+vyAg3yuJAueMBv0b+enyzJ3Zg/Ki+TvLFCseTXZAWq9z9UG
Itd3sue+wNKK0kR71dyhk30E9F6x2Ec/PsgNS9Eyb3x/IVZrLHAS4Y1EneHMd6rifm7EXO3wxNlU
uuLazix1lNEuWHen9MzL9TxlWeSinlIB/bpLgDHAVmlleKMtj2Vn70KpP5c3VbFgr68gfQnIjiPF
iVomUxb7IRHZWhgZIlT7uNUmpr0i0HJZb2O/Upmf6/ZgeVpmdcC2Y6VUrRkHxpFjjUAEwMmuX3TT
ahzNM9hxP7wMQGe/1VK4zm0Q36ppTME9ZnVJJmG2ZBlLz2QIroIGUqAA6BiqKr4G5oiLwwnjyCYa
ERbeB9RK26eAWDNB716GmE4kh4XuJpkGNXwMQ245iqHJ4D7vXrJVrCDIWE0/nronV+eMvICSqHhQ
iPv6Q5ykKW3gs/sbFMJM05nC0MWDe/oeAmW5V32kvXDRTlUgy049s86IkpHYGWGOXpkWt0jTvokN
i2TOzSif9jrZoi2VtQ/e+PImiml5wI/n3+1MqrwxSI0DN8Z5t6ciYQ3kF1DS2WRVBNr2Lb5QvhMl
CFRvEtgnHyx/GJEBapq6/7GHSVtEdFs08mui18FnHjsgWbkZcZsAeqiZY1xv1XQqZhQ1vnGGpheS
zepsyIobsrkb1a8IMmk9PQ1QV8xnSM8S0/OSvwtUyICGVrdlWTowkIXhS8aN5rbNCgvA43FB0znU
aFrKn2mQopSzp5uCoqDFiEh1cZcH0S6datAlDI3hDr7fgZOb49DtnP1R7i9N1cb136Xxhymb+GPO
3tjRab6RdQY2D9ytzYXc1nOmuQxmDOtxReKJXRfen8qz3TtKxoAyMi3jiwsjqh80YhIm+9GrlfSN
9FqrFqUzhxPMYIPudEegvGgSi18LKS9Rx8DEqSHDuVf4LAQe/nP6lel0iIu3hctU54B7Epl+cQEg
4LjSbavLOTeQs9h4Ee0gS2y/QafWvO6OgUoeoJxQo5JAx8V7GPRlcn1uCWH3ll8QOrLANP+jtCRw
eXuyLouGwIVkJqxV7eFA7xAXxTf497/Bf9QJUo5yli9+QZHfdiTTu8PcPvC0e2bCi+AqW8lc6LEJ
+1XOh1+ojY1wrpbeAl+2vOz13I4h8Y1ieKSrI3YQmZGQ56r24nqobr2hHLfEolTud3r7sC4u5u91
VdD0CmcnefGWBs04yTC9UiLxAx4PniEnUbA0bTVJbRhTZk4gg3wHbkBnmiPRj/Djie2+5nmL+2fQ
oaqAbSOeuwFhfu1tP7BwD1Czw21uLiK6fmoUG1LzJ4T4I0hTTRhrS4HxwHwkFkc07Y/KwVwYe72/
tP+tHsTpgAQLVIGLWfcNEZXMn2w1h/HnEa/43edczyANUdteOBsPuZfeY1zV9t7NpEyPsPyiOAjK
8mv66UGM5grnI325TDKJMdb4XzvzHPB8WUvtSUmBVr6uwoTHLLCD9F/o6qNsE+CEX5SaJ/kxstr1
s4oow6YMnp0A2YixY0UFrYwbqXzUFO9u5h6LwbFpWa7ULjYZCzvyPp8dDAmd/q7OBqCcE/5aF4FX
PF0lWRrxHcMojpP9zAPNAiSvDhbiYkiDW/vDUOrFfP96FIwAcAhStaNyVrNcehwEglOssOdES091
Sw44t5r2SDedh3MZTr788CBLw27J9fyZ/eK5adxjGcOYt38gc/QTTP7WjfrvJESb3zcmPAZFYkDA
tUYSKXnYfIlBpxYDVThyXWnAIDsV92Bmd487EdDHluLzbkppfSidHNYncGroxUqXnRL+IT3fTdKH
kT6837RLlunD2OODqbYaSdaAmh2UbuWexMMgKeqM+b3eJ9BndtGMSGTGtAHSx4d0MniC4wvEwHZP
G/iWNhmZ42QpJqLMKDAUe9bBGnKNLPPYXSfLB07R27eLsDwqQZ2h7yL/TyxrlWL2C9bMI8EaLH1S
4aW/Hu6g2BIRqMDKaOZ4+5Xce8SjS/HBBJ9aScOpBRzUjjuuRxX8qpFP9LOOksXqqZBAe5IGwazU
Ky6LC5PZnz9lbF5xh4Z1Py+bQWD41pbrI+lojF9xjEXOvsfHvDcHMDw9zKdeAJ763skcFa9VhifN
J8DHEado2IcmWZKvT097UWSwliZFGJrnsJLISsUbmvjGStdrz256gTHAgKvWVvm9IPGOPjjY0UAu
DJg7plwMLgmFcFVedJqwm25VAWulLXduJBOzHLoZKO4mSnjYmA4JzfC3Mbd8vojV46M/jcDdvMUN
46YXELcSfx7xCVY8m/d2oCvcC748F3tfDtM9iJi55IsH6vRi+4kf0i35080tzpe7z3bITA07f9Uv
KVJce7AphckALHhCvyqmJD+UqidOC1yGhUmBdjqLnavm1HVUjZAxKknFUGOiDtGgQ9Ti4vHB0dfJ
CijVSa1BeKshDm9LtO3EJkWxCcAkoKwWJ1dta1ZW9U5tTX8oWY6K5Tazeek+dO+iAydkuK4ys9f7
2yDms70fhDuGtN2KZhY+v1FSXJ+HruoVkg5HsNzeslr8LvLXQAZID9Jhw38ELv9+ICXuDKOUbQDx
EkZ0xgY2Yd5WYQGdfXBHxoFvBVRfuRoFg2j5nYG5kOP8/ThgaMMfyioo2PzEYkprvlX3h6L2AHg1
MT/LVd6U+KsgSOBgaULDi/r3vBB/P6CN6qZR1+fp490Y675gCjnDucUcX69qmr9SJQKWzYxOOKsm
oCurzhGK2se1SVw9ZEyW7/jQB/X8g2mdL3J69XkRDeVUWCcespTYKNUmAJi+NWyYCYTgJ+qTQdsw
HxCSbuHZVUN514eqHNPqaHpo0y6fvCVfnFPjs94zrUJoLcoXgQyU6WQl6ja7idVep7pCC3rYYa6+
ENnuGNobb/gGuAX3oe8aoXDx5KV1935ZSy4/F5xPPx561WMv5RABfUTfkqPqiT8fF+FxB0u+TBSW
XRaXMB3ggu3ryEwgPyF7RnC5dKT6XoupxrGfFJCwMGH3qlo+4XLPKzFfMS/I3Xyfvx62lM2UzxzZ
B4qvqvPSyWQ6UJuRqNxBjqKoyrpq0DNXRLZZTCPdXakzDibuO6HQP1jGdU85vRxe1EZfwFrxFT4y
PG5nfYGU2RTdqp5s+Ugm6ZtLa3YgTE5aVHkAMGDOsFu2NlM9k2ERJdhE+w/1hvwVFsThN/GHZXuV
Go2VEnbWHaVd16mVLp8SXVRrAhnLNHT2g6WaTflcnh66q1LahW6BUtZilZAc0YXsV0K32uC1l3Cs
vaSWCZtJIZ0yYF5ip7SjM71aVQu+ea9Ro+kfg4FsSME5awhVhu/nSj92hAhaKYeSqvOZeu1n8JVn
fSQP7J08KlE2ewoxNj8bCBHknk+fWntVgY8fRX059fPpTMEiYZyxQ52aZzExaFIhTi0eJpHatOaO
wxiATjYrTod46X/a5OmOQh+tfIACCdZD9Z6y/Bx7a/Ft61NOfBHi8PqU1p+kLm4AVCrEwgInjco+
nd/J9+ydGkAcgXBuPmDzjlMbS/0pkAbwoPMH5+O0gndzZYwqpnGzQocDA9BKDuoSW+zXd5ujK9xe
dyWyH3VTEfywgkQW+HtHyiNMuQqaUC+0lskWhtGxQoY+vwY5WNtdKmlMKsZfYk9R88lb1fz2pEnm
MzeQ+SWVyu7RTFryBBHwQ3tcOAFyWgexEwnfzLNdD/0Ze+x8Kn8wfcoKk7qp/Ujgh14eevHnRW/v
oHCalS05LjZle9qYa4AxPEnPVHU+2/rptXoxHwE+QLa7w3bXeaxYp8S0JVpbOyim4toa/E6MTaHQ
gs6goLb+7xwwzYqETNXABxWlsiuIkSLv9Fz50in8DT+XnLItFQj8bxKbwwPhXvq3rdNJRIXV4no8
EWI/4I11E13H9Hsm8a9fhwnWLoF9vDFVVKtUaNqOLuLy3nBMmCOPS67XiwIzgXy0lkhaoERO6zPz
hLhzsKgUeocmWQNGQCMwA7C6HTw6q/JkZ/EoytWEl2u1DhVnvvmwqZUfT9Di4c7aXbmhFMiEM8C+
S/aBRS+co6LgR2oquU8Or/plsZh50M1uzjbP8PkEIIxjegFjhS2sNP8Kr8KYElEYGcnt6HPEsnwQ
SpL/d5jZ2y9TzoNoRRK+MbAXjeprQI+aQZ7rl84INaTEm1WivGBjSkAjAVy88INnPxjzJKkXqhE5
VNI8PIOHhS167tQycwmqIA6byVUIS/rQNmKxUBLZIee86/MvnUpRB6pA4bhNUGdSDhmbD9t2SUAB
MIMWGY0OLADMEKOHoNvtQf4n7Qo2mzBzyhdmIsBNRwupto9TvgnmcEbr6SFAKDalpL9zswrc/VMS
nyiciewNXiNN1jdML8fomxG+5QB7wtsQOgKPvZqHwS9Mfvq/7GzEx0uaA0oCU+YGkn2Vh+werBUh
aKPz37p8jV7qHV3JRFiRxA7uPeL4ZVTu1L96tEKcUpD2MbFFQC3rZu3alBN3SGWQ/v5gDd6hq6O4
5zdIRq8U5wDQQ+K81YpDCba47IEPoLpDKIJbG0NNVSq+080KB6UWiENT0yqXX0AQGUWMpkLjmzwM
EKmkxwzXL4x7Kkzw0qJ8NItbqdj3RgOGCkVf1taDjr9IIeaQXqtK5iFq1dgOrLLEqMZlYcSPuj6z
KKCMzmSA7LUYbIhsMEfAdfblL68C9Vu1177EfCDhrHBrnGFEcxVYJxqu170ngDXihRWg3604fvQ7
Kny2KNOHAxJ7/OPBQBfFifd45jIvzjTiYw2yFTt2nVVx2G9dfGSLKzyeEWuahI8Eefzsb/ufiTLh
lh2dEInoYHcYWLLD6JL7Y1e22HljeaE1byJgkBboYBQQ8fyU5I6GOESmv7C04ycZVfWREmET7IHm
LqZCKexX88oXe0lUl5GIjboBjc/2GZQlte5mTmx6rJ6OnCaqE8mwHL+R1T1YxiAcyodv2c8Mb5r6
6pRfYK917mX7TceX5I8ugxkbb+CjY2k8amogJdB7Vtivd+8PPkFMIKaGThToJMzwuFoAZIPKAked
CFzS71pBHflKGrTR1vv+4SUbjuhO3TUJ0YibeC78N/Ruw/iBUMi9O/PeS5wGidCbXuEOpw76MPGq
/nZJhN1ghm/Zbh6cTJyQqZoc/bIpKalydd7oNxsEifkeN3hNp4FZLbmcf7e5W7fxwczhMyyxZI3u
uLEM+W6NueukdISrzlifha2RLZ5MkhXKHYmurIvsGqOrlG9cWFfrxwaPC3gLkDb2gJxUEp0YAMxN
AH1r2Nnr8YKL1QFmzyhBBkwQwKe7onahWQfg8E/0qD4kDEkVjkgRFzz9RxmemDlhso0FXkAOa8nz
cdByFAYZ1Kyc24jaCDEXjZQH6H4kvUKaYJ5GbOPlMegQ7/jLJ/4NOS9mzRoM0yF4GVVnv4YF2qfr
7yJ7LYDtziHJUtmfu4qZo+if/+tmCq7mFizpX/CQFV1YZ4iZ3VX0irDSOqLBXu4isIrJEBZmxGj0
q+CQs+27Z+zcdvFBrw8Qbh2URIFjW85LkAEkJMXHUEL3Eed/araAqY1gX3ddrZ4VjUwwNVsLHqMn
FCuPiVS/H5O0WKRChqJZ/OBhXOe3nUKDwMWbTT5P3/TD6hoQCMbhhEnvHVNmobGdP7Jm8ay2L/74
oXPG3H37ldCK0cLZWpxj0BckNRkmYLSNKL6Xsa8mAJBW52G+kvEwZu86+MP/oNSeucvcqmoeuxnr
jp+1r33Fyx+EUXkoy/0BKAsPHe1tBY5N4f0zYrzHF2175bxZ/oT8qktz49icvNv8hhu+Omgd/oI9
tnahWQNOwS6Z9/bWmn8i5AMAAYXwRZmX2PmhqMR1VUb05MDE+ALEBGIw2KtpQ68rx0LiH94bCwYW
3FC/1n4uJ4g4Nj9fIRoKc42AZezmQSamUenyhHmUJmrtVvNJkxMzHc/JjFldE5RKK5mYJxBarm0n
+Nmhl85RAZDS/vcgo+L4USZyJ+NkyRySURmfZhKJcFkAf/S40Pe+smeDPK1yCZYzUJ3FUphrKZPf
7lrtmncX7W2h14UhUZ0IigZNgEGZ4qkshXrQW5je/Dw8EgjT1I7TnS7OmU/SvhjtVzRnb45I4mMT
Rls2l5q7qQxt8chLDXs4R42kx6F6P9SR1GGjdLubHILiXnKo1usu6XpQ+aM3i5N+BXqTEVJSO9KD
Q/ZDlQ1atAVJZ54e0gV2pJbjlYH2h3aY9y1RLa2qzZ9GL/+DRrBnAvJHsmC/NP5IgcyFIrcl6kaJ
r/OSz63vfoypNEz1EfvzLTk3FF01nj+XXxFTssVCEyg8v5bY5jVffj9UOTZqBNOpNBScv5IuJDJV
PnOUdn/hP1WnpD3sZsvy5Ys7xncDnmD8eOzGJ8SUblhWxsNwUolbO2tBR3p3BQK1YExLQpx68DEX
hwI/QZhw81kcXvzxqiQ9SaEWhkDMG+LYjBLQXnn38AQ6LIZbaOCv9YKzmmF5s5UlDJiRu+bx+mOt
LY/Dmi4KpMVXLAYbQidcbtc8Y9QwoRDSbFHwEutaZM7dUKkVfWw9/rxVJlDr/W2aPKi/2Oz9m41j
W7lx7JjSxrZ2A1MAVh/Hs8b7ePDlYvl0AcOeJoRvMgc257E0WiH4K7EV9ESxcrYAsY8iaJw65PNp
mE5/cQ+Ipda3sBucADDneHzQfZW2y4pxi5vrq15L8346T+Ze8aEUMjxsgyUwmq2jkj97KTVTx8tj
vv7amd/Zwedfm2yDPW6A7x/pAI5ESf9S7kSm6Y8JUg6B9Jja1Znab3wVLwh+p4eO9l9wKXcCzoxr
WRqlzLvIHIpujNAqDznu4kh8LLROWWGwZuPgK+HXTBfkm/9rnlE+fPUQh0jsQskGOrNw4w2gYOGM
+kH7u/pL3nrz5D5udAdWL+Ka2joGKvX4b29WgpTYbs+/w1V2tWmy9nQgdC1KVW3tnyFMAoPwu/bj
arEO/G5UZ1Cst1r37YfsSKGlJzmL+QsE9DKQ3HAYTfL4WlZm0p1/N+oGlmcG3wyZiREj8Ftc5dqk
M80mrpGoh1WIiTCYYqTQbKTsewgWhlOOVsy2DV3ddcBDdY6mTFfHLS8/Vjmffp/9/FvdAr9gggRO
8KmW8Tu4iAgFLwQnSURxmWF5dvZtrYdDVCF5BB2WMiCMs8DaLRrGMfXuwf9t3GnKFETjiLbSoDt1
80K/1vieSI9U8okH6SSZIrS8vJd+kCNfzB4pVuH1IBX3g5ut2CR6FFLLcRx9A/6RjMs65fk/FSEC
e5LkapvCLVxVP4YnMzJpOhe2rrC/aOM4rio6rAEGFPQThCwtn7ymm5YF746ZllgCgvbssbV4zp5Y
rlJVz6B/q96C0UO71aobrF1mkCpKUd4Ndn5idub7sH5KHNvjCkAiQEYPYQDdZeMdnfQ4NYxQ3fcv
BeZL71NSv3bm5gwGk/6TL8dAl3uqoKxzttV6/mcmt7KfjCh0E7anZY3PnFDw3XMODqgjoosWc8S9
l6X65/9dcHGnXsNrgQGZfQbsjnqDNkJnKz0uVptXTbspLesjBM+Al0AhFvo13kMv0IFoNr/F364m
NvBmsXxgG1KmjrwZl37R3rHxRnJapTzepDh10HHR9cH5OLd3Cx858bgTITFwxYYv5iXezBDMKnYT
0Qsx6sHvCqu4jT2ik7avP+m2m+r1GHZweSaaLQvlUj6yp3WTPq0Mrd2ryoQuFgaTMVQRRBkyX8Qt
letxGQpTn+m9aQApkyK75dCgzalb76I+uwCMlJ18J6lFXztZs51xoA9dQIcx69QyC+KoP7g46nn8
7GJSCJ/MUNSjjJf+MwH6UJFYH3CazquNyM+MgDq2fzUI8xewfIdIAmN8BnjPYQ074QDU1MgTADID
1YYbs0pEWeWWnvHYUHGD8QdmUxnPiN2JO0thHgm9UVYdhXlktyLh9r2WP9E5OscC+T7J5RtsL/D/
TWT+ENAevqb+NW+nbenSiENaxvKGoRUWqUXdh+qRPgYOP2qdqmwRE7PCIGNo7Tpp8IPr45QVAt0Z
mIQjCtXsTkrN9+FSjsvZqK9le0Iyj6m22XD23poujak7ySheIHy6Iz9TSmZSRrcP+c2G6BcQI8uY
l/ZjlwL7v9iSQ1UGIsnxQozqGRND9lZ42bAy5M6QJcQNF1aiWLoMls+uOVx6OA6ej8iT6O2WWvvv
HksBvIW9jxHdbm7TUVzerPDWCD57VzpHuoMhE+Z5l3nwaC5VqMpS+t5V9FBqGNeKX8DzA46Rl4W5
bkQH2fWJRg/I27F8G4RiI0lE9fWBYRQna8m8bzNr+kR9haamWMaFv5vGOPpJC379Jc2qymQkEM7I
RTA2xbXq+GGNDPyTgWwgRasWkPPOxpOimE6e7Mpjq5p0tI4btPGIa4uRFBG54gKOHS4vhTEo+pWK
xj0X5Q9xQpH4F6YLgL9j4g2sODgpxSXf54K7vXaG/vQmlpDEViFGtnai+x3LE82QvCNJguPHKXcf
/UhmYMZ4B7lrvtmybFY7HgI+hxdCbwRwqvtos/GpawA0dONW6VBtzmpLmeQC7wKiUBwM+DkctduS
OHHU80tfupq6eRPs5hTNNWmBZTGRcfo+tZMzjZj94r5XCMZH3CsTiLfpsXxETgj37FQ4USaSm4Nk
E5MpZxznHjirGXq+JGtdU2P3bHEFUE7IFtytpbLa7n5iRaQf2TzMxwwfg6FS11OBQY6exR6RK7Qi
eHsiVGE9VbZVybz7Nlrpv0zI+QfNbcHGTrJjyNWUmLQhh90YJjooh8ulqaGMp7wzNcJItyvA6Mlm
sSYXFzwpfEtzAbhdfHW8PRq047XwrblRH0MtXCsEmZjXTboBAbUvzFzvxUn3OYFM3zQXtRW57tYx
gGNSfP5CpqvzhSBd+utUA/Pok4rIOmmtmL2zhehIb2oTjDDTLhtDn3WiqDu7O1PCRvWDvM4CSLne
6DLUPHhQrtT41stRc/EiD/0jR9CO9mSKvOzRwkKjzGDNIQ91jA1+PE+1I6m9r1L8spsdknmjcWkF
Xzy+vlTa1FHDk2LZADfZwBgtI7MOniozzGXbj3hhJ4h9Qd0cy7gBrCHd/vlhdNuhPCEW5gBkLTEo
D1ypruwGt8C6j8CQV5BojsO3N7IP4FucgQ3IJgSsStD9TrdgM2FrkcDF2QPLWBMU7EJ8/V6tzOa8
f04w1lcAO4YyHuHY/VO1RFoi3Q+nWciFGdx93+vzfGrjId2scbNf3qof+EcaLPUBRQ9RZ5Ff7TcP
+ONjfrb36xup0bgi58+3FV2JKfTZG0eH1wcYwsqN5rDudRLGT5eLVdvMr3S5o01etsPKdkjMeoPR
aPxYq2cHY5CyI10l57NijtdHmPt+0g9+6gi389V4YI+QCdTAhRW91bbLrB6H1yG+xKPWEWPiMz/U
1bRWf9mg+njthN7JIcaANX+38dn7IKlyG36pviXwvnbnvklrTyECW8cMbwWIuVdDEZ/QPcqEBvnQ
0ZD6DHpWzc2yV8xCjMMtwiXVMWYZ5zsDv23CLWo2WRU7YQHXkbODz+XpK84eu0lQJqZYJcnUIuJ5
CJMqafzTkEfrF2bpaQCVrd8NNmJgijB/re0EfJ5by/o8m/pA50G0f8T5rCvDsyrUil/+YJSijyNH
24a7Mz3w+PtT204LDN4K4sRvE1Rn+mDuQV1VmnZRUQH820aH0BuwC3gPShu4wQzcOG4AP8yeQ58l
GP7CjnNpqzSTzn8EVdohyzLZxwUSHgFfEERXqKCK4o04J1FP9EXckFeB3pgYRB44jid9eLYjfaj2
IbUPirYXw00NXTwEFOBBu560kpuKyj/yhiGQjYoSHM7fqCmu/cYo7HSiqVl0srC9ZLacJrgWd7qX
h6cpk6AzFEXfR6ZJy1ABYfg/dGv1C9O+mKnsRUZnXzJEcekelO3saX53yyG1OnqRqyxzZNbjKF13
ku+9oURllfz35KCGjwTK9rWhFO32lo5wpzejo0N730vZ2wusEMrwDaKDWiDOZIVbDNV5kshgRtgX
ToAebptC7U5Gr4/AwyWT+gF2vM6FY9d20VW3jzpFJAoXyD+KqXQDQcTBJpnuprQPGAZcEJasvvSr
/MUSXFftr2Qn42dIaBSC4ru+c4UOUMHHk0nHsnTiwvnia089S+Kbx9AzjV9BKnmIpIOWYYsPF9Us
ap0QxxfQfBsuWL4SK4dJXBaZWfQfQ41Z9Gcp8gE57RYx4OavFa0zq24edAp5PzT/Pc0cwJfuNoAL
zsRYQf0qye3H6ESSQHNTgleZXEeEGA21//bU9cUW6y0L+oxQFnukB4JuOLcoTRt9EY1STuiUgZ3g
jMcLu0Rs+taHkqpufC5DsuKvOY+7vcVOxYA77hcrTeGI4U2bpHizEkF+FqEc/KZ+bjOiQr8MRzWG
HWqY7/QW3K3r8zWWTIaVt4s93zeXy0KuaVtb+V4rJdqf7K9R74QPl4/+myfym8waDjz8zqxOhnho
HMe1mEZ6jfJg7wFZgykxKSt69CqA1OLizmqLc3MOGYs7i969eg+HkzlpOS2/NRRQ6NV+nHvQyi1n
3Dn1nmLeeY/5vSbrVXZHYy01yLqLBQQypDgHuuz3zmYXy4rTeuE+etKDqzmuwmeyCdXBF44Y8jGC
Nuns2/58eLrR3ZNSUViE/3ynSlNDwtJzOg6NCI2ohV8Jpjrvo8Glg/cPUbcmszGPROoxyvESAHom
2bndYl2ZL0Gm04JZmOkRdTR6Bd/K2czp2okHiJpTgQkmP9tzZkW7MBhkTN5e6ZtXGTdPTAitmTc3
3vNXgvsrcHn/xbeKYh5bt+yxQCiI0pvlyu6xkVuto0DODLPRnk9VYNpCDtUp+zFfWj6otMmgvS9m
oS5p2tPu1gnFRzfXTEZBbvu5AkdEvUDMrIvxZDughTwiHTUAWpPIB2hn0Rr3h/7RXtlFlEsYd75/
82Z/XiAJxeFk21qYnIf6r6WzezgDmRCKnNA9z/umjESzXAhb9IRxYarBxTseGDdkz81nc18Hurpw
NRtAHco+Tzt3GqBMmsNEX+Vpbwri1O5MBajc8nXM7IO3p7JQ0V2KllnSxdkDxnveVIlV3wiRK+Sz
37BBU9uvt4nqtdUkc5nk+YeMX2ANliVlBMYSk8nSLDfK0hsbeVmMe6jHcGlEQOT9pUx/5mWXCi3/
ltNgCPbFFFKdHjxZ06cfjLXevJveh16Wo4sBkdIar5OqekZMjbdfw//tJ59MkkeHB0gte6zZizH6
uGP50HrKepOGxek/ItbFyGr3geRPp5ko1pqwDQndo9p3jCkcuxp/KWXsym6frBgiFqgH53PlyK0a
CG35cr5ahB4TyTFwK4Mhi4uq53mbeZTtl7HL3V5zgBaD8YZhcier+oQ+GIFCww/LaZeCQOkLHqmS
fflVfNcEYcHX2pAaMKiV1IjLKZVZ0y3hJonJdjcisvmjrsQJ/Rj575Y/EFBRRSruoIYS8cSW04g1
PtlxHMN+jWHLSmlVN3fi5eL54cJ3B5x1bjKfbO3hEeBT5Tqr74KO8zLST6KCBAlvLrcUNLy4Ziea
cILG+jvaHwtNB9PoqnQT2BVPJrWVXuUcLusC83zy16x/hhKXKPuU5Lg1mwLPQM8ZsMJWFv8JSowe
aiXuKB0/NrJiGTNg78Ghs/5Deg9WTJJlcQ0vphtzU76TGrF0lnHO5gFHPIMm8aFH5poAgKYR/D1W
sR8YTqpGzCq+CdDUjDcsO9s3FkbVN2I2OzH1pzbapVJR49nKv2kIMQELqrqce1JmaMq+JrPnQ6oL
mO4JcblVzkStVrAM41B+VMcqS3rSqpowGKnV0DbJDHY0TdWgs5L0LjoKVUG6QFROzedmqhG3l8mn
XU+eE8pRCDC2+BUJgvCVA1buWJ+FYqBrIabUrJ2nGZtCiyGOtCj8BbnEmoGz3PeEqa5SKQQkZSYg
ysM6T65EbnkrZR6MgsLbPwds+j08wNa+FaKW6bPykFqaZdFxm1jvIn2EVe4jmhdIvt2lfVywKRI5
VuiMewR5hJrpNrqjksYlhPypj6Fcnl9vAJo1A64NuTt3VwKWPcHz01Etyn3J5pXq1Kpp7wQ1fcwB
9a5DJkddmRraWNsRO7kGueQ/CJ5RtLPjhP+zEtFwUXbPZI0sFtWr4wKwxjNFYgeuj/FWo6LK07Gl
4un9ayfNLEISLO5P1s9mZX74g6vAWuVXZG0NK0klD/fwFvdsl1MhbWWDFYbpR4dVKwLcgYwLgHMO
o/C9EXx/Dv2d+Q7ckTQloeF4O2V+i4+AJme920rNx8vB0DdYzckQlOfCinISXaB1ebQ5vpwGplsF
xx9m0GNTVV2AkSidhv9wDopZw3uHBQPPir06KVhs6NhE8M2iKena3acTqsaTrRgVuRMOQWviBtYl
N49g5IOue34N7dVVRQRujXt8NkyAv3MHN0rUpscyWENPWq18B8v0dTnzqt8SUzhvl4450lWzYqKb
bbxAvzWwDlXQ5nPZh44EZ3kMO++6op+tP5Y2xx7Dh7b7W497fdmsjrWZVccjMR0ztik9JpXzESs8
I0gg1rfCKFAJuiIQwpZ9/yyPnQdxigILWLwk0Ja1qHZi9HySFki4taWtnA5CRCI1CZPb7Zy6wRYh
A7zXWvlPPZG+Erc8ZzxudOLcYH1uYAjzRsgb0vnPlYO+gDSIBWZ0ql43Y+RYVWgv5lTjXRTsvULm
JDVzL4QCVriY2t3C5O3rk41Jq41vDO1nufiFzhGpP4nZ3/5CcXSmSNws9lVre/bZwwh46QnG2LmI
5g6UFmwNr/aRalHxfnxeaY1wSpLpfF4xVZ+jPhlkaWh3YOUcrT4fAJjf9p2CCEXog8OqFM0yWcmE
KhWvM75fYxlQgBRz4A8lXnEAOFV7zSxEs1BNIkc1vhTnQ2OYhffTrqqtqKQ4tUI936BYpRGJHTgC
ijfx6rFu3DUU2yzDsdxpfgEWW+FLHhRTwNIhkUQGVoZNQWVNL4i5raSShjeb7TI9LY+2BZbMdGyP
83sph8Tx7+M+7DwdCZIgjnvUIRBFTREJ2mKI5EOISN7DAGAu/kGFoO6fCQD+FrT2Ge/JSt1U0g5q
HXTU6uIfeKlyLQSIr30um8THg8JnGcZyIU9C6oRHILy2cQTHSiYGG5xjqvsUgTRdhj8oDi9PifEm
XgcCfb0sV3z/KeXiLUoYNW+DiyldzYIh8wZrNcSYpB1mrQ9Y54L5jjf55XnMy0L5KBupIWXEnGNE
EgK1TxAoL4eEe8bxO+bW26x8fWO4KQcSUK2cQ6G9tZ9YS3mwhXdsvd8brzsanpNbOdj3bgVWGmxh
S++7laLjFepV1obLtuJQxMjeex8D/oAlZUUxMmSIV7bdQdTgbcXfAhaz7gkZ5u9DuCkIYzgbYhRO
mdeWeZxErs8mwZbZYIRhiq5lmoZGZEnfOUf6CserR3pR3VyJMIUAjY5R9SdT5U2hqIUEwVPrNg1c
GgVPbuoxt5c8oQtOTn6nYmdy2+9C5Hq5ascxmDQJ/epnniv/VAxoWGZKRd4PSFcsBQfQWm2vp9yp
ZaOXzjWV/GxQ9YTbe55aQk86lWj80a+U8gJODGOH78EaDP9oL7MSEFnMR6vDgIdM+v0vePx21l/H
84MrD/xu/Mg9PgX2SBq5tVnvBu6PUXMWFtHjUTRhgzTGQxhTIruWnlRq1Nd0YQKyM9q9aKv9OJhP
GVGtNibdsMVmFw5sKM5w0qssMokLY4e/LdrQKAfKt6mG6fesem0lw+FQtiWgdTb8RKTseI0+QCRM
txT1GrChKErmXMhy1cNx33l7g14+3o5/CGa4stkDFMkaXq/UX9WC/Hbv5FmUaK09FUjl52HH7yme
Q32KD8W8t5gY/Sbet08HkvaimrxZ5BOAj2VXRm6p2lvMuSsV4y8lvA/ElVOgTdlChwylnx02s0Be
smRJV7TPhhvLsaVRYSYkZfRrARJz8mEo18GhXajhZ1xSwi66oosNZIXd/iTVup3oDdETq2hGOI7t
5ly9abLfi6P5iA9djxgmU+wFCSy+rSpa5g7bNrgDQMXGbKuwnMNhD6Zcxw4L33MmBtAwIn2d82ge
D/UoaIwNbo0hDy+Ci5xOeB6UILlWjLMo0RVqQz3N0zoHG+BdxEfHrU+UuiaRIjPZvSKAnzltkBBj
ALwgJL5U9D1HK+0nHfAH8ia9YaPjdC3fB5W4x/4ybvEro3sYwwcmcHNQsNx4SlMcpP14vJmLVZLO
k+iDiw9pEU8ifjhs696NehfeCXp3KAbcGBepaKpewbfsD905X4HvMYaVP7HH2+styuHAeCQkPhWk
P7gM3Pmt3alsFaTdQYvvBj87G4lE+H77uaG+bC4kZJz25BCunMTtgGvgxCtDTlBKWpm9P3cU/Elf
CJg9zz3ojMrVtvvWd5iVb49bL6ulRVsSo4ONUSFbnOfFH3TsLJ6AYXRiEkD9DgAmGkuo4U+r9zHX
m9B1HNmA1hq1L85PvmWd/H6dVyC/jk9zNpWH9xspZkQORxytqDhsq3wNTyfW5hUQ1mSiw5DyHKav
ol5SGpul2FpjsH3K5+rMI/GBhAtBzTXjvEuwMFHzdDuVpd4PWzJI3RtLvo/X+Nx9XONbgj1SAdwo
gCpSxAyDFUR/T72qvNu3MtFJ8ynCPyVqSYaWVPphMCuMiEAtKFh4h7jgBfBgAgKtl3uIfIqs5k/7
Q12sr9Ir1BPaunfGwNCzP8d1hRnjBASIf2g9M9uL0qPXhP8MaCyHkD2J5hBpfhH9GxsoFA0J274s
X4h6FD/ienmEUqSoifL1bItnYABbPphzHSyQg0Hd+j+2YsrX2uitf2F8kxoHGBgPp4WSJLDZDo5C
OryPm6W9Es3g+6t2Dsd5Cg9zec9XuiNj6kFOUcdyHmhY0mrDmDQB5SQdF0y5bLtcTNYf6xj4w5RS
+cxKwYsbuvfnd920iOhWmzQ28V4m6pJcU63yvxxeDl0b3QULounp7zzM1AmrDz/LPR8cUqDdOXFg
WxXOhkNS2c3SAuMECD20Dlpj9yztgC230qKSOK48VN/mlcTzdPnO5EkiGVfWeGPsGMOwMEtbgLTG
jv8MO8vvskLTHXDAV551T3O2ar2Jf0wTYHKJ7y/HmzVs4IpnEWaEp31pjmlPTJhkED+ZCJpd4tQX
i+qnkRAkmTTGhwSShVxDjcwtHU4/kiyyNYVQCh4VsZ725D+aX93OKd9PJUamG/C/sVD5a9t/SMDT
+qLHj3j3aaBpihsv+F0PsalYfB5l9B+Ic/9020OcEvX0t0HhsgbJc33wF1WI/Hn4P8tZ9YhXcy18
B9nbFpIKhVxiLWdbZmPf4GuwSWao0GHRExzyCYkBRjiyz4J3ttG1pSfppmJC3vRDssKco8X3+7MD
iKgyAkCAKzzCa90KDKRqh/3QZvOZoTrqzh5QlI8aH4rDz12P96jLhWwLUTwpAGTsY0Z2orh5mSdR
vrbCqJ4Z7QOVTiAFJHhqjL9ZxGnXeDzjYTDpVNSmOJa3u/L+tsL/PE3Fp3vYt3WgyMJqgLJS5Zu+
dLZ1GniEE2J4AUn5pBHwMNOA8MvsAvxBLCtg075upyNtW0hDLWpz+bUwQYRwbu8cXOym1Nt8zjYp
AJH6HV1nrvSTJdAWXEDOw4dR0JmyUmmCWGw8k8zhjP9NzjtohyDa073vg6LH1/+xua/sIPZ2p+eS
9fHKZiJx6PKw+IAtagcrcT8h33B0qfVMdjLsWCrdm3JFGOTfzcSXx/DPgIg15cgc+/KOFX6hDqtC
u8SaMc5HUH7xifck/iVI6Ug6jvfK14u6E7kXRLDNnXgU2twoLmXXc9PeA3vDhelIulEflW8gzuUr
bJVWnYBsRpc3uMKsoq1azTP9uiVnOT9XGGIEzmQrOI4sNr9/Bi/iTm82teeTjJFKxWy+IM6rYe/M
E0p4HdEdplKfTZDUBpv9JBvdWq5klDn9AaHSBoIMkC8IIHDJ28fojcLmKYiTDKNzYG4BAlzMGvxd
KD6jzEyaDekyNUTG+BZNOFLBbdqLtPttMzMCVtLicYf5OFlgLYbdSR9BwxwuoXGlBwrrDGp/aNEp
jJXtmZJmPoxCy6/sbcwMp1PwXqldtN5oVhwToMFXzXwCXYoJOa1p/Ny61WX/LUuMCLSKNmJFrXth
NnamO+bvsZAOYRMv9k3OrZRKZ5oYcZN7KdMERLK3h5ZltU1dmAgzCXDb37UElMw0lq5urdNMNSQ/
2Yf0bqTdnWm2sD77ZCDwvGD2sLY/qS4hDVGc6qZGFseewT88fuQWxWzgnwN0rLV0wsp1F45wI8KN
/2pwzMC4VU2EH8oxC8+FKh+/52gbOobawfkvW35mlVDHnz3ljVFTywAaYsztm5Bw3Cfg+8FvHq/V
0gUKRAsbGElepaQQyBD/XmHlpXjkHgIFbabRWMEr4LUE2pw1hlfZ+6u85vJczI6IHDBGyb6CGpZe
K/zVVxKUHxnqhvdwnrqdL5l4yfEqfr6+8A6M58sQJ/jH01z0BsFyRaVXGeaYuthU5g5yQ3jYper7
gzrDfH5tTwAhsi32fSlsAWINL2boCyeZHR6h73ZoZyW83MXIGCkEmG7Mh3EB6QhvBFxgembXl/ln
hWvekTgDXXuhue8bnc7QrpEEbV6qhcpUcBk4J2KRA8eiK8hwgSzg+MCSbh+ON+1eRAwXOcFYQYl9
b9/iw0OM0W8LqxtFFtKg2dMf4ioCj5pIEcGhXPpsqmKi9zWwmLha2CL2bR7YnFFEjF+YULMbk1Is
bFUgekRSOOKJbHbPDUCFs/nJRxwbCZ22E78c443ofRoGvoaXz6x+qIG9N0HNmtisWTshPPUrX1GH
VtzPyNkRtxXA6boQqUO2qe+qVEEjrRUx9pRCgp1bJawUzt4L7FVn0YTqwFGMHpDgBs9l1tqZfbcq
ZcYMJfLEv5gBZmZgLwK1mC6EFd740G25yyKksZ1sOj7h9N85g/GlC0r5fe+Ur+n87NfvkfVtF/VB
zBOZgY/LgbSJhYJ7UHoTnUfLrG9pyuQe9TjLe9t0QkOhX1nDxl5ZiZ6j9jC9EYjnQuC+B4X6nVP0
muunwbXAvQs19mvBiz8U8ccaReB+1Os4QrPujneUgUbfw6R/2yLPYPus9i9ZC4eT112v8RESJk1e
aonBoD3XVWW7e4wKVAhfXLxaHf5nOHtwRSwWOD4mHDfp0wrHTizE1tzmZ2twYVfJBk8JdZw0tzig
2BGdxGz4V8gI5IfDc8vcQZIPlNEHM9CxU+SbKe7iE8vEhKM3N14lcdEyhYXYB+94E484uRYAygTY
KlApFssHcoijX37umi0hYxHm0MlHP9q58kTiV/4brZDWttGZ9sLSnuN8xi31fOd7uOc39wCHD8dx
91hS0uMKGReXtNrwzjE34Jonnis3151sVEANrZFK/nP7orqh/6DOvEnqVQk1Lm0L7LaPuborUYAX
UPLi1cWx4k9CYDCdZ3YLv7sQZhFfGK8i9Ru2uK13Ui8w68y/+Fqx60Uilo686Rn2RrDQZ8cMB1e0
cad+DtHwXOKO7XkRBaqoOv44vbJDve8awM1lMYpqLLIafCziMdLhNOuYVIn9ofDk8XqFsFQKah9/
u2V0YrraxwgkeBqHhOuAqMB+RUL5/ahUA0l3Pyq8HtfyznfjrVJdKRdRX52k4aytnxkgZk99EUMm
aO5Z+MTMyHIcjXJ6dXQKy38KShBWAgAQf0itZzMcLu+mPTGA93AqIl/Srvbd/VEa4Loyn9umJ6lc
5gWTha9wUhL5x2xA5F6b3PQFrJWJok3qbj78/8hfqbKd02q6UhxAYFSWxmPCpFtuT0ziZTh9cT06
qHKEwO8JjCumaXY68rpOH4HZEMl6fLdxujFPpQjQgNoS1UjV3fgegocOsFSgpFitFwEprdYtxdvl
RBc7t4B/2Yxmd0srwANht+e1t2SEzgVXlXhtyl7WzfQQTRfMpfiIM3BUQBm84MkYv2jURLf9JwiN
PH6cacJVEQdK9VnbCFtRcSHDSZ20dzKQMhv0jvij8cqHG5ZPQPr47VV/sSvWQxWyvyo2ruLgGWKy
f8qoZ4+3LQddqpgFJ+/t/cR8+uLIu+VRPq/eNLc/3seqWEMTZrJ4ZaqZJCE3jxEGq3BRs3Nq6xlo
SAheqPA633gIL7YZYfct6nLHPcLAYY1qXKPNx7NMnN3zD8LVgaJYv8TkMydpQ8usrbLA7hP6plsg
bB9TifHITaxAUqqYdEwcBtG4NXVj/+jrlKWM/Fv4a+8Ktdbv6BHO2VX7qB0RVMEve38OOytIUBsC
S5WPydCSdM0x+Cp5qFlaOxRZ+4LVBLCMrB7lQM5sYqDHCGcFHPfVBjRxoA4T/Ev4xbtbff4VoMzS
zy3uaBYE08jcO4y8OpEjauGxpLrM++CA2PYjGoc9JfE8WXtiQz1XlIb+gDSu1cltXKObLKCUJjIi
p390vp9Yk02/VbTUmiwMqqCVzA5W+wOs9u3wI80e8xm00lDd91K3wBDcvZI2mDRPQ1jHcD5+P5Ma
iv84/4oxjyk7PYzJgLksV+iR7UmJgCjeqbYjsQUqFw2ueyxv9ifI7Vqjfr/0ldWdKTdIGR8A/jgj
Xazi+nEGkDZrUHsHmhq0Gh6UU5DF0YabxjJuhC/TY0Tx5CndlPPcIU/Zl3XC3/hhEokqEYxxGus3
9IQmDfPPGZPSv6kgn5PmGOrdNLxqsAE0UhH5sU5wKdKDHVKszS3vz9JCJuXxJXqMfgUuRsS3HjSB
qQWmvvX6cRr9EPQbJvAuhng2WcubB+bsbn7kvuZbSsMckvu4YNoSCfbZQxecMluiP2Oct8dpITPN
urqLDJO6AIjyIyfi2wXx3hCyXRSAEkdYE2jEUinZykcKx2zvIVLMo3F9JhNpe7hKgYxYeZtfmbzW
PXlG+8j/6BcEI/Xd636tjWLb3mnPXqrLDNaKXvQ8xONudFDG0aljsg/a2U19zZattOJQBL/zlO3p
4t6mj5DSECekp/C61czGAO7wM7rEDyWqe+A3X1/ueuRe4+ftkfZ0cAt79f+XHvseKd0ynNIFP3ma
fZznk19UfA1q99ADnZU2wdYVy3eMl7cyfKfDB2n3ovxdMODmkmp2ZLe+NUZtp0XboU/7v1PgjnLB
WeP5S13Mr6Dl64re2zGOyifZjZmAh0Yb3CGfTeWldlHAxRkP8XyvVOAE1wwqjlRBQIad1j1K98+I
fGrT0oLJtqZQs7pmgXlZHZLQfz4k7UYBGA/NdDBGETPz8V2SNuYLBXIccqi2UQYz0af1KAhEQG4x
1RzbEu+eOMDqi4pB2sTFfqunZm2GxmofBDzi414e4jcgOlGlNVwKTdz4JVKgwbg1DtNMeqx+Iy4w
ssdesZHkor+2q3sH7Utgtlr955HVG4HeR7iqQYpZysrxA6FjSN4mFhxS71uoGE6T7cvmIiJ6eXjB
ZmI8Nw1ocnlGYmHZuVajTMolmyb/I0IeB0bbNErRKJo6IyPOUJ/czVx6Q0kcwrwBRn3vOQpZsnyw
xNuLA8cTNQjNrYh5SXx3M9MaNydjsjto6cQw5K+Lpd+QI0h3KWhZQ0kahKiYw/eWk0LI8vUOJIiG
etqaqgVfpU6/qK+AZ9IGEP8JV/uDL0F6TZVGVZTdJtrQXVkbSMMD1C7vZqi8XiyhNd8rXIjt9x8x
o6UQEb2H+pNSKMvlhs8OFI7+I80Dho5ZkG7YGAb5iyMlqgYycEAg1s0ZzTh8aYcyH4a6rhm0JVK9
nQmz6TbeJRWfX+S6rZ79cI0hnMeDzeJloyzuV+mP1MQbXVfoWMxqFUNfiE3PmsKBZ7vz5RT+dCJl
Wl/x1PrTkUc+BZnL4Bb+8k0W1YJpPtrC3ZIz7i3XqGAwKUlLSJaVZnZ6p/sO/nFtE46I/JlMoBKX
t7iAvEfF+/QEhmAunhXijct9mcwWGmfDbSR670plD48YYBVHj7DGg1jPWwt/GoIvsIGWbUrr4uWu
rwAjoHhFSFvXTmccPFIMlNSnx8QWU6rLXyWKb+lXSBF6Fy56qWmMXDXhhrH5b36EO5+rYB/1ZxRB
cxUOjEM7JDMWhxZYsJF75Kdn01JwOLdOj+1EE7+oesiCT17tF59AbBPQVHbUj+EFhGRUb7muqJuI
KQ9EFENLo7iUZPw7WKL4inq8imImFNCNoki9KY3Ij6EmR+M2vfGA+oyQEf+6JhZdXK84uzwXLewW
/a+pMUg1dcZfaC/IwSnC65sZClK0/pDY1EOFu1vkLaK2VZ5wouxHSGVh8Wqfpvl6re9BNgM4306b
2u7S2W8EGIicAE4G0fiDlA/MtOCzXRj8wccc+Zy4asGWnJvnUJqjETz2wnFJP7m2faiA0W+4zcPu
aoub/+DrjYoMnxK6tf8eqwWUqGMEAA104l5ZpfoWofZZm/ShSmLBfjgOFcNGLm9a+B99hauGRohi
AKjMZtv5RGL4vJD1VGJUNzJ6IHfMKVcbG/7+gOIV8H9Y/k4gH8UZ8CDTVcxX2FXem83qhjcFS8XO
AciayPsaoqmy+VeV89rxMfZF7c6wryht4izL6P3KlaighJgNDYMK5a+9ecmYG4kdCiv4U5aXYJqa
at8igTKXnjKFrP3QiFAbuqwTQM23uXritUvbaiIQWaURJ4fxmaA5lxtzJlaGQ6dJwXgs2+aYPO1e
PjEdVHzRGvNWCixFN5L/c4ZkvfOZbnxdp9Ot8WF6WvcyEq7Gg+A5Ve6TCOeislnEMSuB9WPWVvnu
ARlEUqCCcNh+4LHC7rDslUrjBPwNEDiTinSNSEo6e3Cxj8ikwaYQd9ZYxh7c60YFd0xRvVtsmFKv
UJjSOf4qxvx3me2npBg1hTcYM22cibRJQ4HEKW5I4y0gS2mVLjhjTeCjpoZGxI+9E3iRNo5MzOtz
qkSYtIH01znnHVakJ/Bdu1EWFLygimCClXDCQffLunwpH0vEUNJzzqpbQXetZgwvqZ3uoL6i3bIY
OxNmKXCkVqpRO3O8rjeVo4rp47RS48KCooCBDfMlcv9mPamsitFUVBRdKW/TRxc9lASNYfc07hCS
UZuld4JNJMa+D3xllRlrjs9j6J1jyp/33ehVRDx9LRCsKop3CWWYJiOoeAKasTDNXlF2v7ICTr6Y
2U5t3m7YbKwHYei6Gmu0h2yEP9fXRFk0MHuzVmMbeJ1NmSKFROYFl5g6B9SVAcI+79hzeml9thOs
Py6fiXWqGIP/Xw/fhkffjl4NWgEePFWqCjN6auXe5PiqPokXkibL1wfgrUJhYimULaJqtm49ne4B
UHA6SRFbN9kqkVA50J/Ca0+KVYabw28EvuO4KgxZ98+qjH5dzCtYv4T7OziqCJo5vzvjn2+OH2mV
NKEO9+LFFdUcjI1nHRIV3Z60oh9SZqWW8ABRCMYK7Ic33SM5coXEyGwOTgG46WgjLn0NVBr5iQea
5XyeWVm7ktTsfKfq8uGMPjQ+nJdor3NZHfjOsEaEgGchruOHfHpntq6mzhjCobIbx2oATayTkhgt
hLsqNaaM6ponjYsigFv0SMJsjMoFmy1NXQhDWkmSRCpfMIxBKsDpkkXQo+YWOCtkk9/C+jqq5wlE
WPhkLN2RIRifwVtuUVMFQbqWYgRDc6OY+N1njmL7DJBAE3Vm6xYVTNus2EXcFEEej9vQbIodKTiP
hxRvNEbnVFlZlXRQLjvbEIbvtgXH8gX3IiQeTpxa8YM2Hf8tj1681l9cZPT4x3sGdahKQi+cZb72
K/tBc0yS22BH8T4bMGqTGFsh2IWTc0oNrbJ1wDsPQE4Yj8GOhG2uD08wnXiPDYaB99waNrboxNJe
rxmPo8CY8/LrOehURv6pg8E7fF5cEiQRqMqd77OAAsI0GqcKTmQaGKU5B6UKxqr7mg+b0uf/rhbA
6YuFEg7BGXrdcjDIubLxed2zH3XecbA+drUHBZFHhztGzIMrEYxBo15HBLSV8snbirCXkRYcIyIa
isRYtB+8LZ9IGxRvCq0FlGbpdj0iJzUMRskUjCDCIPZvUcH2FFEJI87MQTExeWAb/JoGhdkzzf76
+qR/Rr2q6NjNXRky5WzY7dNmsct5LHudEcaerO3CYjKdjJJyATeldt6sml/IcHsoCvf9p579CVNH
dxMFTExgYViUFj2hE57Za84zz0R0B33SsK2p/75hUYT312fb+vcG1zLRtb1C16NvbZ8dI0Vakej1
X0XX1e9hJSCRF4xreFyO19YorWjAptqIcs08yLdIBS7sYWlCIvRi7XL5cIqCxXnUesN9YipessGq
xRqb65Mjb6YPxFiXxRbMcV0Lf7wcmVMcLW03NesyRzjAqbQDI7K1AcL0jhGaqQrp5FGLNJerlrN3
VuIq2zyeyYGv0iPLQ831PzxlzhUSxWXWPnPKP8KP3YjC7XHFwWkgk9Rn7EUw+WqlGS8aKEXZzJ6u
kLlvntOY5qWAy8gbrIKNK4d2kppsEB/L6l4vYY9+YLbKT0uVi1MXLwn0LQNIIu1fJ+MkoeCVwhcy
MJCEPVyLohNiqELb6dyzYB9fD4e0aOZcv9nCMMTXlP+HUjyLYwLpUfKQ8rJe+6ipR9tsFG3W+XN5
+q8oDvwxTrkE7SAhyMZaq2qC6/6mfVk0VQEEQA42q2h5KwRqBSoB/02LJIiE3xMt2PKlUKLmSmup
wfftYUDHtSBGwIrOlk57TFSUp/E+NKaZSJbw3Xv+N5fE69yLjml4Z2hpSxWhEqe4IPnKMy1lKHnJ
vrhXNeJtlaL7SeoiBwUY3KyadkFxSLzj1ZY4FIqDPSLVLD+qrgKE/K6PshZ69kD/SttBTq80XfL0
+OL0uRveatGDi01kmeibDEIdOK5lpHBPtxZaW0Uymafzh1fkh0wvvNpJx7qR0KiFh2ethhjX4soW
DKNghekZ+t2JR2izgY+PuB4dtltqxV3sgbQm5y5nHO899rNSV3Fn+1MX/YUWPz5QnY3oAPHYeNfo
XayDy+l4ByG9abg9oDA7XakbR6v+24+GLJMThPLh5YzXVbvBl1J/nqORoXlfsT3d7z3dva5GEuVl
TgiFnFiGao3Y9cNd+O7+3JzfKRIr2tXokEDw1G9G9lR7un4/SF3mcfsWFMKrCOdBHXOuhgDyvayH
5S2OvVR8lJeU+X677tt5T1qcYPfxT001DdMxGnTYfekk6Bf7Gr6K5tDZjgQ0OIVjARNygO+M0fea
lKzDdvDomKYZcnXKoM1q1VICSXt7klNZqJQgaC2CbEYLMr1L4nuQN1zaYjefOWu+qsIp7Xh4hwh2
hyCXDONq+5WT86uth9t9ZV5TLn3+C7375k82mG0V+SP/9R/UlriqOYYPb7CVPB1i7fAMX2s2xWXe
iBa+npU9beZeYd+dR2nJDu4R6uYdtmeOj7I5KM77JJXB2turnGcEdB866xEIO1VwB/rDmXJCcBpX
Sm40wtVXhhHzz/ANchNpboIu9uCJDsXlXykbRKSD3rvBhmq52SfN6y3XRcYiDqErAWmSvMv1iD00
5tEJQ8vYImai8vGifdGsEoR7dDmzFyS64VXPxnF+nGErcoWQJ09Ekl2PC/k+TFRFWua3U/L2XCjF
O1/xHWyrEDAyIaZuuNReZwDM6nChetUsRR1T5Gwy9tTvc6EeHIDVHhn5rsCdwXyG+7Ltod7oqSrE
64aml6iDpOU6j4Y27d5owMPwHK19Lj6eTsCBjvL4+La389sPqqXiaJydgNj8RsqUxMeT6k9clJ7t
tax8MO9q1bnMAw3kMuwbYpEiCXblzs7VnzTBtZ95QhBmHkM8tOn86Lu9NjjQ8zVnwBE6fAlAc6Wa
H26mJPvj5Qmx5APKkwr9MJngYn77YMZFvtmG+VxQu+vtnbCYQrjmqQuWrQLii8krnkbu7AI7hfNX
cLBl1bfHKNipW6jBBWje8BlaWTrCiTRVLuD1hU4O65y4SFRbqa/LDAAxyRKa8djiex+R8up0gbAF
JB9kKmVZrbsHZSNJaYgcXjPNsRSmBq6ENX6HEKTD8aqwcSuhlqL5KWJk0xG1eUz139eAhNobXe4f
vUsJAWNoP8O4MiyUzmdwYvsJfmItl9mz0JnFQ2rrnPCENX9tM0CTmsDBLIlwCxvvpu1UR6LMZCht
FRqW05TIZrVBiKuoUIDOxDgt24BDigycdLalg/MBbKBIOKGtI61eosRnFvvrGPKMqzTu5UzLBfpu
aT2UdtpMOAw/S+ir999biPjA+I+FSX/583t6CK0+5BZuS/yaN2KPwaGJT0xAgLKJQcf/7OnEWjPG
EPb89LMJFyqr1HFPWtqA7FhKghZnwPgS4CROHTx3U0miY3zQCB4Si3TMu8HxDLOFWpOz2Pi4Bznx
AqNh5Hd1GsouDmr4lnorg8Q3EJltEWa1T0Yup555QgXPc4OdWLPJhX0PF4qgDINNaRCEuvCXwtN6
D1c8GvHL+R4nGadjFEmBKCv72D2lMX+poIzNcwEUAoqy8+nwQhXSfM7y9bBn4ARHFEt5djvm4oAf
+4kbBkHgqANieuL4gjjli3ZiBPE3gUIx1OW/1lsRx+C5Lq8LyGM0n1/Pt+VlNcYQPGqKFb9L73xA
QSPXO0oOOZ/iXpn9a1NJUFLZew3bmYV0TCuiT2VOsivUU6jcbz0kUmsGXu108ljnar3uLNwactbv
59Yiqar+Lyo4j1pq1ohic0eIQgOqnj2cj2r6xsAUILsxpaXsyJY+GKhzyqFmgf/IcJI0Kxqu4oGe
LAxuvnDb/Vbby5mnNnPW3aGpHhKpBIWKgoaGXBL/qXYQjuFPnSxMIK12EU2me4Wqz8s4/kHj8RdK
lNl7ykcGXca2LEubtF30ETNmu+61G1010plJYbHqHRua17+ID4FZFiEg6SJxIL7f8CA4wUM2MCep
PVco9s2pI3pGvTrAaMZN2FfpiBP5daOU/mXJLArj56aJr/Zh3bL6OXrcTsXHx6ahlVGbsphNefhg
KfTWNI1yP8YKxEYr5c7QumAB1ymHU8eojD2oMHc6T+GMMETYOzFF+qX3URVlWUODi0aV+p9dGnGZ
h1+TmZ3mAdU6HxQskVnu3SPalGg9newBT+yN6wyfKpmfJHLlZorC0LI5oX1e9EfDlSqNyVYMVhEs
9u0Jg8vcbsjl2gouvVwzeh8Q1lB5YYfc2sCrSsWH+33wK2IF8YUbCPkAqTmynjnMechR/i8PYKzh
Dty7DM75yKVIEgLeOYmL3Zyh1/AaZlax5xvvthjIw9edPjAJ3LwmluQZiYaV68uOVRN1Ilp9j8sd
r/ijitcfp17QlehCRUrXzHQpWcQUYgAjh1pXbHkG30DGy6j2qoBmG6ir+PCQDxUrkbJ8TkZP5q3q
HpQIFY4yR0cMzn/P+oc9Kwa/bElglcxSnufJw5hivfd0f94D4CaVnt/IQJumvATSp8TsUUj7cqwU
1d3FhjC70TDk0+k3BUrH1J5pX07KuVE8Ufn977zLKyyCo780DXoHAssLObLpIaLDmX7ctyCuY8RL
Psgjoglo1LkU/YKTlfNGgBEPEnPXYwqJ7ql+392u1uw4uY0gsS9k7eOkV80wOjbasgx0tnFqXwfA
1/mwCd4GskIAGrScRvVnBxOC8yCtMk9AbBh7yLJmY0OtVZa/gGTZwUMMG5xoCqbOCsGPIGLwK/Jq
HUEhRhXr90+yitkhC47GP2KcweLiV/7vRXC/QSPJgnSWaGd/nkbShERPnks+Wbwjy9wJHlc4TlND
l2D9Tv8G0INtmD25OGZcJFrgzbvLJnzi614mVcYvJbt9bVpq1U2fNH2Wu2vsko6QOujgEmvguQBm
WmYojy3hN9kG9YYra7FLONne+SnFq/wmk6y6sQQ6X5Rfm2j+2Ayx13qxi6SiFc9FGc++Vz+zxvmZ
WXCO8K2YuwuD66lqfyMzF7T0n3pTkXjPYUdF4c40D9azt+sJSqywUidJtBwXnsI/WE+wHB/tZm5w
a1CPAKITKaQmnFz9mn17z5OyCqwjV+Fln1ZzzombLihQpFLdNrdMkQ+vclEQqwt8aI8ZJtHpdOHR
Fc9Xo4LSjLFadgAKgel0IjRFkVk+ahtaVyJAeuYJkSSYiIXjhdsoAKEAdOjYXV2Cqx8+oNMQUMJS
DpjGaf2DkZCDG68P+rQAQiNSKVIhoFFxybxSyFfQc3tcCa/wfJS/bDnGI0mpYCUjQbGW12jxpgCU
ssnbXPom4UYRRiqVcu8MVnrwVLTChdSCy0PP7uuZrQUrC4O+fl8rXQWefrUydzkIkgVOC/0Kot7M
TmcCn0Pp5mJoLf3qEIs6OejJQa+qzmxXcg+kU51nGXQzAbJylIdnLhPXYYdVApi/cCPH0cOpEfNc
leuHYKQu5lXDivIyh7j3pu3z8k6E10oHvXDE8w0RtzWkwcKdsBVToLQIQkYZTAf+A1sUvaAQVWj4
emJJjpjv7PzJTk+1JpdMIw0Okabz4rcz23cNDvsGB4CxBc7mdbhhwpVddG29Bex7mAbEtX2vOaIb
ZdjPpevsASfU2UjH1GQOtZE9OaTdD0XSyaOvhvB3k/4J0U4D9uVMnu+a1VvbZKFJ5/fdnhnW8Z/Y
WnFq4CCz3YRsN+JLXZh/f96bkko95yIh1Ibo4Ngm+udGdEnFpew33qjJnyORtzuBwQwQUBzxatEH
4xtv9f1trLz2IZObuj5B0ZjjHv68u0+Nqn2WjR/bAO4Crx0pTSs/L341vrI8wkbvtXXx6qOZz1fy
AJ3KdRuljnKBbR5tFeU2qScLOCzGca9xVqo4w/z4LYL65JATPIOw1cZjT4CfDCTAelce7wNTKP7r
Bk34Y/FJA3IKaDL2VE2YUw9iPgqD3seQ/lhz+tyT6nf2AhNKfq4R0j3FwhQ/diEz9kTtDntw3tNk
iLxfV3RYDpZEajjX2MYMn4xRhB6RKJbNXW0U+hpqSEko+k4DOpdNVtjFRWuXqvrfgO02/izD+j9X
FBlja2zav+NclOC5gVZHSelXy3RCGBUDY6x9xSj/Wo8R655gGEl9bBX8aq3zGDdMmQpfJiEzSIB1
jjYTKjdHlbLNQ1+uKklRhHj6YTzLuW6hbe3hUXX1mgOSd70ViVj+6pisSxYH/sLJPRg5lU5Y6Tb3
NCVtsSzr1lggAVI2k+FVMjbLvMyoEKVNp4UjvHqaGVsI9DYkeD6sB0wjdPWla2FwnKSgx+BpqVg+
UGDx2jtK/w1FaSZWPAA+YioJFbyopLUI1EFg+uzYKtK8yP8BvxauZbnPq75/NXmAwAEnU+gukaWH
Hor2KeJ7apxsWJvp+8JGuOV5zK8P+yUYXC1/WmjpOsGV8QD9VrAbjpDXUyo4gzMq/M/+vXRSgeFT
mw4ugbDN+A9WgSDoyqdm06Sm/B5hPjLFCCZ/R1f9tfH6gW7GjMZ7GhRqH5puh87QSoQb/Hd3dkU7
K/j3CWiFvCpaPavttZq1QQtfrj+sfGyFWRAJVoKDtCJaqLSXPy2+CIohui2xn36Zwv/NNwMQrEgM
Idn4Qbq9La18F4knpleUd5lMRTPosgfBXHE1UYMa3ma9lrzdpxp9ubTIX9t74uU4FqHxlByB7MFn
ckbWt2vRP+qU7uKvkcwFJEeBHyrriXhmVgbezh6DTYqCS6KMuicl82c5sC2V+kHZr4BtYImOVfl9
ddTee7fE29hH7jpcfwy/tgCPezRlr4DKKnLXfKwE6qh3O7U7+6EHJ5ITwv6/OYzTePKOvhRq5/3H
1eG0c+D1bLwKCp7oEQgizBkdpkGBoArRrOd7I4Mpdi9krXVWd4Feh1rYCjIjJr7MSbaQMHSEQiAW
JySF7/RSHFV3woZ3GZ1SxgAz72mQYaPxezx1w2WKO3wyvgiwe1xagFSusV6omWBvAp0wZLagBjbD
3vXeb1JfKZ7+X7UONXI9gaphiulhcTOvzGEwsqP8MyKdR6VS/qMiDo6QPd1+RB82ipdQ88kybmIs
VDnLx16IpeTK32+uC6TFrLyB9PgCF427P7BJitUa2qrxBR8u3y3mZLIYIBI76/QNsN9enq4zDKJf
pxUcXWTQJ+3HeGU0Z7rM16rU4K85FZP5vjRvxtu9iu1ED1g4y1f/SYpiUXo481vvRGh+iBjaFfzH
OJpq2vjhjRQyJ77DANHraV8vE1yDeOejJHONoSxOuAsVTGcJz/DDW49X9M29Vzv1EmFrxNICNS0w
zDgmLxJHqlpzJ6pdvI/TpHO4wCIUJFkWbL6GRtfjpJvg+Op8JbrPpgywYS4qmnEvTo2zS+6sf7hj
ZriIPD1RCTSuO7dW57JdDZaZQrzytVMVOdDpDAntHxD5NqT7TH1HGfmfRrq2/SFGhZ936NNhy/NZ
KtOt2S8MKJvZnPeasqent8u9cAwtCSywJR8odboodRHJzBQYirWNTt69nzM5o1X8a2LJsG2ky2/M
o9ZPV4sfN+DtEtJb/SFgNil0Hq0n3R15ZsNcc2Qnx+jZZJgGNVpmeadxIxBaZ2OpBgD+q61S6hy1
p+zPWxrCQjUpkSealzyYrEJhiMewC3q50SS/8Ww6SdVLQfbcNc1bKWSavFLJQTmQjpD5YXgBDGk4
zJHGQbrsrPFVjfEvVlMn6Ei5BjjKTtu4XFFajJgeNmByBZR4031mrjnGRi1RqBA1K10QqQSZRYyw
3iku60+D8QtMSqsn/sFG1mUw/wNpDm3PIXv54a4NsRP7hCm5b1TQwmEiXaVZ1B8bInr7jK2WScvT
jO6NfKadGGu9+fHeXsxrLf77vaswx3rQUyocLukGnqmU1oZAS4Kav7aHZiWi+jxJAMxWApnhYn1x
orv83ywmw+UHONnKH2VMlr9KtErGZ7lJUEK2JclxSzCgufjFELL/70IeVef2NFSVOYXdH+5nPuB8
+DAuYznIXo3JRB0fc1umM2b8GE5Fs/Ssrt3QQmRvXQXHorxs7h0IXQBy7bdWcIu9mIPAc0oEDHs7
HaN0cYv9uzhLKxu4E+CwKbUvsV22BG35pPnnnW3DGefkB6lmdMLjBVPPFK4SIPL69qEi98c36d3C
5vbzoVN8KBHKECM+J7tWsOIXo92DfXbu2eoI161PqjFviFRaIJUbd3B70HEEMnn8GxoEELeHQUjg
e0io49Y9Ws2RB0FIhJ3T/47T2VQNtwjZA2FlexJLuNYVhlGtqrlLcc7KaSK/RlPr9O9gu9cDZJsz
6968loaDY+66Yp1k01EoPAsHM4Hy52mmzXDQbOVm15O7viS7JG7y1q/OsnQnPd5empMnO0XeYG8W
3S75ca1+LPvv6vumg1WVZ/uc1kt/MzMJowMI/mt+406MiK+aQSrX2UHbAyyEJUJjLw9N2R2AhSsU
3VJs2AOpUYXV2oqqG+texikq0aXp8AV32LWXJsxkRFvqbWPxrIo2NC6M/N/DzmFPOkp0wxKx21dX
gni/Bn7yOfsrI4Yy8JmHROBA6nPhnmNfsj3U7Bd3PTDIVvLmU/1tB8KQXtiPQNnZqHj9IOxtUYtv
+B1S9TY64CzZIyFNggafzF66qqutKta6dhPU6jci1N2m5M+DGHTu42kHpqvyb+M5Dfsd5aTVLGTS
n54SOTMvbbsny64A9hG0D4+Ir7xWEP10sSRZIUtm6zWOv1xUwNNYht3xgJ9+TFxZbmf5isM28Olm
FtHjbgft7jRx54dmKlZf11pmuYEv8nj+gVZ3i8txorB0eq/nTmRNf9r8uZT6Xz3FpCpHuGPeQ8rf
bcSYNNUYtdRRU/e/TtvdxUojaHfGpEt89zX6a5ng3bvxfyaI06r93cw0eLABbmhhmA3jO5Lo1hw4
RS5sTUb6DCe52lCyBAPgcPEIxl+Uq7up2Rd2d+XApgRz4m8y7V3cVHhH5PDEwulz6rqTSQ5aHIFb
r0Ts0pOtpiIzL4xW5kFHTFH0dtRoxdto0KvqwFjfjS7DsXVVCzELm/VaZOEAZ823O4zIL0XH2mPY
11Mw0Z195jlzN0dkTldl+Hxggg2nkv755vcdZBdQ8Ke1tnZiedaieYgtkdwF5t7rDYcp0QtZp11W
kCqZObMz9lwht/XcQ0CWHW7InlygaSyYTzyWl70vLhxLDxTIMdC7Naij2+118dFUC1cnYhUgGOTg
Oo51c3O5ImwTv6ZW66cgks6n9MH8UEHSy8oN1FkGL0FFZDWsO5xJzvx5HK+aXic8qUNqQGNzF8mq
pb71tsDyAvV1HuxNNaQiZF4JeQVBrjd9BUIW+id0qrFDBv9F/h1tTi5NMpF2OHwRqj3v6SA6aD3o
JehX9NQDr2GfUXJnVDBHFuyOHF3U7cRAl2TceSjLZhBdIgxTnrd6tZb6IEAkmKX+UmDBMMBQOHge
reC0m2EJPmS4cUfnfDYYWkqVSkk3ocgokzb7I9xLrxHXGJ+NfDf47nPJ9V5++DsA3qcGH1GE750H
nUpPeNZogiGK9g4U2AwnU/Ex/FQZKcnaT5FUfC7MJUxSrRykoFnc4Tdf7R0uFpf5g0lmE1LmUhS8
VLjfV9dge6jGeLkBMt+kdtU5dJr99P8nIGbB3x3BnmuoTyOQgDN87dARUA4Pk47rSIwJm1JDESQc
bt736pea5QJ5qUVQmrh8WaWwi8tYLRnZWTDEixHhsAPQ3D+NHv+JXmqDJWLctHrR2e/748a2U6Kt
jkOJ7iIXqkbRF4kCFBaphJl7mEO6N2+Y6vnEYnkR1NNtNozKZ3hKDPWPQOSkN6tcZXT4IvXmV5pd
BaSqFT9BpSILYepR5ZgxBMDPPT1/cDkgG33/ky2X/AfGvXNNWJRAHP/Nt3BmB8shD7yYit1w4ciT
2ruUZGj2ZfiIEHE1NZxpLqhTPffs8hz6/VJmT/p1rZG1DliqDyzHQ/l8Gmde4shXYwuPutfVkO3E
kJuskXa8qfc51hUr9GDIZRSC4IAmzsmbCuBW2Np0gDinS//gD6iG5/SlbA8Db+4fRvL5R5UjJUbT
Gz6BFuXdGabas3NNcmQL+Dg5xxAjQ8IdumPpbOgG0Q26/6OF66k7VLjOGLgIQzm954WOxW+6T+Pv
gbrXsHdmrYex6YNG5De9ocPozznQDEw3r+8ZAV4AZrw96U6rgLf0WY6eqo1E5Qpj9IAUOjSeWb/u
oZ6jEE6qjR+Hyh/m7AZ/TQJzVqLZNJ4HgTPr1EOxzwm/b4GVmXIIW+oIWItBjEP3JC4AkgFgCEdz
W+m4xd27ga/LEsRKR9QT4y+LRHN+VGjlZHl2n5XlEqq9xbtclucZBbHWZxS077o1J+9o6FPvsKm2
MZpGTUiMp94J+1W8iFSKy/5Ty8iCGSk30ShbfqWF/CYfaJZH9n5OXMduCvZwtQIx2EYTqNE+UOIu
cDuG9zbCleZvkBhiDPetYjtoLdU41j1Uodx/jS8o7zMc/SItQe5zQsFBjCs+u/jZLLdp79bIF9uN
6tEOzjmLqCKrd9SqjiqlI8AqSZjSG8zYj5GdcgrR1xaDcDuVyNhS6Ba4NqGqUAErWNTedbcWwTWa
gzOif648jxZm+qAzJ6IwreTMaoI74obo2J6mM9UzZbIjHHumMeALu72K3BohY4vWEVI0DMtV/26/
R2LDExxUJ2SGZ09TW7i5w4WrJipU9guzAz7i15ta2s2ylvOOupvxNAm4mHGRvoyTjJfpLkpTbYUi
coHEo2nkEu9CuKernO+4K7aIb9nnLPV0ogs/O6ay70iBIQgkLpR1MwTvZqVlFGI0TJE56tAPbGWC
iSuZjFmxlJgtTBlqSHcjxO32DEuxs1FvBTcupG5ZhLw2KK7wRMavFK5D5JhfPqxj9IFi8MHbBYHp
BZ5LSQgB0ueCFtjkqykxJsk+0+BTz+TJmolHYUtKTuuh+MDSFkKHhDRr9yJzdisok9OmmjAXjBlI
sG5M+P4pkWwUOF36Ietvt6v4dTn17FG0YZoTxAPo5Qxk7D26klsea9Zv7EZgwo9H/KWtELAFjC7g
gJsftmUw5YPj1a9W6zrVh0FHhXW2m54FC3rGnDE5ehT/NHdvQ8tE5IEpld0GewTvWnNh0zSS5TWu
a9InPN8+speVC9+73HGre43mmA1jo38co5fVdWQG7PSscEa3fG8i++6wDICbUig6tp/qGZE8WT4S
k8L86acw5YKQdpZ3clAcxTX3KQa+Fu7W8kiPiQranuj2XqrBMdSZWnBBT9olQZ5PQ1UnFn5t8SMb
3Aj+PAyHtXWafOTuG93wqCh3tSMhXAwXp593w48xvRIufs0+MNzAcEwn+tAoX++fGqCBmSEZkgQw
D6Hbpz3JWg+yIwYLMJJcVVpaMaozFi2YxI2JnUa0WmBA/beDPlmqA4rLvgddrdyxxsdeKc6jE+ZB
fk92AbBTWmdOCLPXo2VQs4SknLzSaZ0EwYbrksLM9Ea0qVy8Gp6UY8mW+OmG//1hSCuPeP9XU9tP
uqKhtticwGc4VuCXW/VP1B5HHFlbIZXO23KZ1ZNzk314BhAximMWmVbP+ZUZ13egKvVR+JP3uUiS
0nQwfxYY65Te09LsXnINN9SeGB0jNFa2LIJPKCk7O0YJAvKCK/x9IBYJmg2pD1T3D8ClGhfQm+Mv
/ThIZ8i85vLRG4a5yJaD2paryc3v0RgGAaP+YVvdZmAL3HhXswHmIvmxVUTFo1CE7qgfC20405Fy
pkcAcm/iwpR5Sfy4cQZ4Y7hxyEXesHyZ+id8DymFE7J6SwxE3XnLlyZOZT/JPtETukBeI5banoNQ
zcfo0WvrSCX1LjGM0YKzLBknJQJP3GxcOloTmVXqWMJS9hbz6FLGMxYmdIEydWvAKvwZR8MlKZdG
KRxgzyFFbElzDihsreMKQJP678dCvGfXngjb0k6TEXXcbx9vBbVNeVbpIv78n0dwrGMxUpHMqTYy
yR8Wzx9evgs1PrfTNgX66WEmSu3Z0kYOwsCHbedAlcFKXt2p7ZYyh0CrAhkexF0OLPMVxYPmOGAG
3wOG5BOaPQxz+qdhpPXGPZ7Him2JyhTACfKxQORS4+uAiTXLwLn59dzb0HQ0o5vjD+6C4JNgpxgN
pKh2VSLVVhIz+cCyFj526oi5Jhbo3ldf1MkzM14waG3RFCKrlbxh+c4BxFsrn/duAsFdt+tkqEMu
c3B+qPWYcgvrdq5txQHYYVY/+xV07pA9/X91/sqVTpU9y5AD2v3zqMfNqVlfAFx/UkGUzINhiBtf
ZXP1Trf8vprIHPveW91FqVeUN/yd6yiDPw0ST6fjpqioQiAHGyfr/xk+b29oDDUjpYro1ul7VT8Z
y9TkXhQJ8fi7moEVqQ8PrNpyp5bbYncP5feNJEj8a6Ep5XDt6zNtCQYLnmom+VKC7Yk6wZjwmWcM
ahNMn0WRwpvfs30KxOk6oZcvDLxYTwbr44UIJxChk9bLfC9b5/KAInSBZ9YvQz52OeO51VYckwIz
GJ2JO1eAsSBnJc2EIHumovKFtktBzpXNNCdwAEZmXV/MHMG7wU1cS/jOLKv9Js31iAS4dWqQGH84
UpJQJFkqieh8LCkdfcolbi+AS+4HBX9T0sPb2pFVjl/vPhh+Z2jA3PIAYm1WHa7OGdrYHjo3sRxn
+Abv1GALBlA7n20wqpR0ius1ygNArIUMxeI7aCYWEnEtGJhmhcirSGGPKt1szhw/pFnDeClkcqeI
eR8Ns6Mt3y/NenY7RbbOnMIVjATvmIj4Pb/DUzG4ur0GtB1DWFx9by526FssVXixUN328thdH9r/
7qwMDC4Ub5XzADc5yZCQtPYxRszlAxZBccB06RjiOzeUj6zNWuJsw4J//RFwvv7t4wI8XIWFhoEg
dz2sB3DMiW7JxpOvCRA0dbsYbwYEJAlvqV6tnTbhDvk6Q+Kmlv2OflBmYnFWJWErwnLTn9gv9/Yb
JzL5TGpgrdLcHekmhB1vLl5STrd97ZOcbof7HS5x9794a4OK1QN5zj8O3stnlktdwS5ljAqmC37i
gROxzTRYbynGfAOuhxXZU3kG6HLrDl4c6M/Yb26pkr8dJxn9dFKst+UTOUhuCHECudbcKVZRAJDB
B+atKddgiiE4ea46CPC9L7jo+Cwl+86JcaqQnRcnVpvCaeAvCf910EwHlbtRyMob09ptmQzmA6zz
G2MKhgoOP1ghmsAqA9EkP6rVa1GYlGTi6Ch1ES4iTD/xW2cCMJ3xtnWGbTEzScA0v0Kz7MvFYBPS
VB0TV2wBenJXgxURGem1LNoq5VIXyMkdLh9PPpHh/R3uV2TqV9nb4B2m2PI0BoZbY/CIqSG+ThEa
FlM1Ddw0qOmKaKnnJw9MPXUTt+ZUFlFL6zIHOK/NIveJAok1ANggqdVC3G3K+y8zWe6t9rFPZPL3
NBRKmIBQjLPud5Ub1Y8JxZMRfaeoBstan9RMSTZdIMUQ1i1EegHmmNXRFGmpde4XisCgxdP/6orX
lW3lBm5RMfIDkRtm3OEMxh2Q//y/Tz7Nz+V+AJf0QGPW0/Lw2WUD0qK8Z6raDi3G1wLPqj3xK7kv
Qw0UqxeTozpikz15jqTxBzK24CoI4zCQBZhPeeb2ZLDN2I4EmCsb/qPqMQ9gFx0VWU27ohnyjpbT
qPzAaNsuR/sb6yy5NghMtoBJtM3r9Rdfm1uIIz1o6MTGmUXUQIkfyut7uqUgcIeXM3YO9wTCVeMo
oOy45wGZYOO6tm++ax5nzim3irhDbTQoJ7ynZpkFENvunl9Zd20CnEECa1AEUjudnr9oXchWqO/M
loqV+8uCrNYV0mqB8ujS+rmaVsAFmiLDbcCJikAdpmYUcRjDN3yeKxWdyYx4RBNaIYpZC9pFU3Ma
KiNBeMQqW5Tu7p2cHdiT5PsJfpS8Gq6Q57UWQFj6TS2IcG/4oI4hi9rO3MjNqpafdXiasHFyRjsK
yd/XRZn4KllWYk9ueeLvkIXZYA6SZ9v+EG9qytK0jPmWPGU0bjlC1opSfP/h2usf07t3M6nBQAep
Qq9+qdEHpiDpgfEf6JxeL0s1H8SorXys1lOrhUrsmXTQ0FaYurVw/Bh5iITOV4+0SVykFrz6o+HW
VAwNSsjEuZ4fk/zFoLJ8SBjnP+V8Sy0+LbrrHL2IIcHhksbN7Ox9FX+Pu0Ix7PT8VEMfMccMjyfi
4opMZLM8zGwLqTBvdCtCyWTQQCBuQ+lDt90JFUQsGuRRy9yamIFIUd14Wpg8DRCFV4JSBnvR8Qyy
BARyx3wHka3G5bNqnxqxfJFXsdDiCPL0rUV/AlP7/MOmjdAvBTfqs9wVfPv/yNYorb+cx0hawl5C
QIIzUniohDThe9sGJsXScxtwnqbjXHVzW3tzcMbLeVIAJIRf6b3KTBKwEfBR8KKqbeEVWcaZ1aJ7
2at9uWI/phK+aSfqosgwiyDVfVfM2OxiIQMDJFdrTs/1La9X9ZQ+q5axX3hGK84cZ9oDOdlAV2L7
9zBmjcbLohx06ZzUKNSS6rw2Vcx+k3kH0LU78J3tp5e98m09e7bf+NFDoPjj2I+ubrKRnQBU6wQu
dfQWMUvmLK82FA9wvqM6FYGNb2auHru27jy2DOGt73z7Z/wYun6yCzXi9WaAl4uZKdfTdHX/FhQw
X0ofzcYLSUCukHL2rpN5ij5hff4USgkPNgJhiW0c5njatqGs6hBckoMgbTo0FMQ1aD1EE3utPWjs
UQVaUkCGlXox3PEDF3cyHy705X7LlaLxxr99xigmiTvCLpfXDxA2n3Wcwmo7zrI5dXiMmDhi+/wm
R4ui8vt6IAUuvRd6m0PPoU0x0orw+1zQxTTQGtkwXzqjM7MqqeAEJJsWTcd4dhhM5XpCSziQjBPt
mPbYYl/d+ngC23c+XArLq9gfFtdextvfZmT4dSFR9RvE4s79y7WcgZhsrJNECIA7TWwevqxJV32r
KDdZzq28QbPIm2Q+8R/aCoBFEDCOIF293x04AIB4FflOkdFnLAvwGL7zo1+KLi2vJnzMzESrYiF/
c6WZtdLAcrXdlordlI/pzdCqKUKDcpHg2LNuFQktz+xw9ZrcytSUiZ7pzILNqtaevKgb3mFFfyGq
fMkyCp+ucuJ4iNf2H39J0mf9bihGgsO3pMYxdeEoAEFTbAEYhHz80Nl1GRqnks306KtpfmKKvDvD
jQjcY0o0wL+usBLCdpxSOJyFnYd+RF3N9QsjIp9RlKlz1BVqd2wB0ebB0oCpRkEw8zv0+jNHHBJT
Z5tE3Qm8cv5EVj32xe2nYhx7BZR2BpMETHEhQjOWdLwh6TDQuHE3+d4QLVJaNLF3rY12HhFVCkJC
kH/ENiw5LkKNfe2TDQs3fODwNgNkNkBoKk849iCrl5pdd+nBlN8t500bQFoAfoh4T8I+DNhdcYxo
HHhA2Ww/bl1M+enFxpGCZTKiwZlSQlOlDo4E8BT/Nw4xQhndgXxdK4+bJ9JNy4IYBogIhatX78R8
mPwRbGwK3GAo2ssNzcvn1Z6VfKkQ6kT7IZuJPMbltPyNFHOIiiUSvU+eMkAPnvGD21tA49b6NK2d
xCKCTQ6qVxKSy+yPFmE4DuFQIN/uiF8dV3lrDtJ38mP01Fpi26Ch62jin3Z/5O+EM0hioBHmzUeP
HowW08KtWjNg1w2eT4UZYhXs6lYvPIUPFLaQSJf0f2lEqJSAFZib81zDhduqhdd7lCfzXp10zKHh
aXt4CpOFSrsNBfROU/PU/WIqb7ndcE54iYTBmyzlIYN4PGF1KdxaBrWdWCWxWOWZfo0glXZq83T6
eNj2k0K0E8I00MHWSbPPiW2TWCyJhkXtq6Wga8VeVLLEQo1NI2m3uQpxVezVlsgf5nPmU2KSQguH
h71ny3U2CgXJN1KhuDNIfTrYsn5t7ZFHnZWSBJ/rict4G9g0BOJtFig84nnN5u0MthYEFC52Sd9n
YCxQfNMx+hnR6Qp2GjPFBHGkYUY2NKb/otFm6+c+d9eJHVYJl8qeMLXLpPTcW+q1lcEMivKtlQIf
GZ/dakKlkzz2Op8t1m4JaLTlDfYlj7gFyTc1e/6rYGa+sxEdI0RS3v1ej+3RGM+tx5VsYp+e4QIT
Ln91MDqpJ8dAJgQa/ziiMe95KzK5MxhjN9p+U7i1+US5am8yAtnO5b71j6abrjFQDjcrKlVR1E+T
mnsAZizkp/i2ihlz77HvyKZBUcGpPIedZPekAmv/+3oNnR40YtjsxIcnxWpOD17zqPom8aL4VRP2
cr/AHRjsTS/dlOa0ma8iq2trgnVcyT+/2DeRyvYtYc48IpEHxn3nPgeJlF6hzoHjMsUHRJFNMYt+
M5qiTCJfCrkL02t9opm8umhms2rgYB2/XfCXIbC86OavZlrtzxXOyUJnDjhsPpakN5UEOYGwsUGL
7dd0ofLwIcFhjaM1kajMXiLx8bS2ijlz/ZduagfdVws1g/ZqPybWq2/Bd5Y3kr6CF0PmnHbzUZk+
tBLi0p2+NaraAt/TPkDVVsS36Iiok7L/DwNOkSbqFKeucW4ZI9zj4l8X+qpIbSay4YUmkTCCUlOM
r06cutxKKHOdLsDaYPe4GgM2hdudbeafNHxJ8+NUrdBvbC/7iWl1AY3Ib9MKTJolQlMjebaxy4X3
ZsK5wLUs00Myg1me0uAePnBgCld1SG/GuNmAAIfGGVL5qD/GWiFEhjSZV3P2v2txJ3PLRRLqfHe/
ZYj7VVm2XMWhBzihh4Dzmg6fr9vfVfbkqr2Rw40N6EugtuLUcmeYPFgzJuci/52b85FWmmR4TvEi
btUxFtC7s0iU9kpxoDALpLlkV6MKq9MpG3W4ZObKTzvjYmHOM6LRZ6948kYl5W09k2JBu7KvGVWQ
Kb4FFtLN8Zpe8Z/mSbPcoxco0TGeXP+f2z32vw0D1ox37B8mIc5coguvASp8DFvXmskLadio6nNh
TkpSh2LabgSSrpJmiibEH2gh1NEjPRKgRRNGX2euvQNiMdVIw5sNh7ZGeZ3sdTW/Y6twhvihJjgE
erx0Abvf1D1FoDxDpqUGIOcOZC1Ro6rZ2AiLQ+yVMR1Obo5cgIWTGFlSYjkT81LvLARyjXpo5dwS
yV4jqOPo1SWczVJh2Rnj7kv8H+GhFSQZkPy+hh1JW61OW9RIEyswT6GnokA7Lw+knJN2Asl6b5V8
3ZejMkYywRyh1sltlBtbS6+Ik7ZVlvDHgrbodsmV+OK2UjCWcm0ipKO3Ua7xYNThBHPF0ZLY8Q+E
mQIZH5xteiR6dAGueTJtJRD/uq3n7mEu1lPEZCgnQEoSNC2bZeVz8unKwXb/94EBA+ZqtNhnrzh5
PjrB7heNNNEvFzT8nSdPOV62t8nY6ZihSND43HhhVb6zOQgc25tjSDC7atK3gVGBCPtfBaIny40m
g5Qr2IURin5oUr9LCaGD4ThSdMy4jqjJhlhXwZiZTesPm2Kq3szwz6K9hTdjPoMlfTj9fBoUzgJ/
ksEb43qnqrxviqFwpSQQI51c7xgO92vWS5D/7IOAUUXsYJNe7iLa0YSu2lgZScWo1OjzmAEd4M8H
ul6H9OLAMHpeDsjv4g/DVJ3lkTpH4A5fPkOE/habyCfRAnsvzJJfophl8NIXJgqHkNGi7uAOob2O
eBZk3CNITyLKe67UZ7f+ZjdjqZMj6JPgg+XqSq31kYe7MeSG+2ZWngvCupMxQmIwwUJLspsIG+JJ
ZAjmmR2lc2TLK7nc5tBUBU2UXL2OqOczHJQi39SE8kkVS8JUCNjQueN7gwhhA208+9eQB231ArVb
m8ykyGPgN5816wq1PPWgLfGj0TLx/CJkPGubstbMoBQI7f62SOdtBBvf/6/gmBFQS/g7B1nJ92HP
Q23BVwLNR6IcxdNpu00K9Jo11Vb6mRkc8JlK/sNiZom0sGIncHn8sGwy0OLNOxKQ9uFQrccujBsc
61bCoM7dnm9a6/EIGW4q07khowzWJN65XV98sI9v5qBgcn8+dvzY8ddKzptwh7BlsIYB1us8dUL+
eKGrBvPhoJuFN2+k3JolRUAIkG9qdH6+z7SbSk/drJehfkYYFoocR+dWnK3Y7qN2ifQc+dkrCkUN
eCSWGAWFPUP3y+OZXwPwdYDPgu+up2ttCjUwfu4A+zhoYR6rJWe4gUk9Y1bYOXp19TdOBt+pa8qn
9M10xHGlvlvI2huR7ZCSay2OtUw4UbggaS73GJLlE5mhO3NDZHvcjPILFevPnZw32GuIuQf4PHKr
7216+qXS5SY43EGmvE6wpkqx+DWQZ2oL1W6nXBD8NQvP6OaNtcfBDAKL8t+hqj93+DHH7W/n0kZq
YpQVqGUmuZGvy80M0Ol3ykfNQs6gu23twp36h2xD9ocoiD8NqQWYfkg9UjRsEZVdO00mWNMvid2f
CNv6SJIWANhKMtufPZxVYRykr4rz/jEaQCVr7vnNEvBHFUnPcvJHmTHM1NmSFOvOJSB0yTUwpZeP
lHINA+LlmUQtpOE9bObbdvfkEohCsysDcQ9mNNC5D3uS9M6hvwCB4vifZlZwSiZZsJjWA/qwUsOa
6NYEX1LZ/Luh06JG/RpLoll09IGbpjtF+JD3aqEY1gOskURQZr2pFZkTbu1Qrf7lhI+ApiecV7x1
bfuQHEIWfLoeFnxHc8ZxZhkzWv4XRtSYgh8OsTHorUKj9Xig3xjNa+CIgPbjjS/ceSQ5+7cn75cV
/mpglso3wLOXO2Q51VdkxfyYbHIzS8vWronf0SreikwMr03s/Cr0lbT0bfneF57Y6JaGF85lFTAG
er/g1XkiDp9yy6yVVIhhiCZOZ7Gf9jUWiGa+4gTSxkI17y0GE7/30BlA+ncn4UBV6zXe7/Ve68RF
4yLsSRtIw7BG6BJyHaeVRwy28Di1p/F445uhXh+RTpBV8qsFeeFNyUxiPLA5teTgoE9NV5bao9iA
SCcjA110GF2PKR4xqFFMdm6ItuYDtH48G5/y3ocrK5p74STJZZT9dT9AK4tI/EmbKweNgseD6Kul
R92jPOhqQ1Cpxt42ApIy4azAuNebogavLDdrhL8plROrBIuvYfVXn7TXIamMreZ3gn2HUC/8Mos5
QlJWG1/4EFXJ6VEic7+AZVdV8iht48nbjDs7domIbmLEG1L80dLfnTqxV4+E3T537+gOnJyAt91T
RFLub/0bLvTQNIUxqO/X9uKPEpQBtETV7LJwUJWHLZblHXB96Z1zWZxu+r/63S9e2+b+COBoXKk7
rIAp6yh3Y219Tpq4G5N4j05625pJAjtljnf0wihAgeEKamcK5S5NYfz85QbZC85a6o9z01lIUmH0
D0uhJVqqyhp/tqUCS8A+RjaOE0zLAFxJEK7wf9Rsvg8tPApYY+aY1qOwf4Xd7FTFqR10ZxqaFHlD
C9rQrNEmPOT0/v1ptD9l3n6BCEtZXjUlTcL3wX895gboW3E4PnT6of26BJpMWPjmcvbIJnbrlBQQ
rDc1HwNpB5pTt+aMUJA61S5R/nbY+LFyNVK3OuiEgQw65jJ3IWrVKZdDG/5VLtE5BJp3upLHVcvp
BVsdg8g5ct7liZDIiGyuq0CB5u4kjYUsiBaRzYAQPiEefQm1m0GDcg7t0HxPd/3FfPkry8AqA8P5
Kj5TEhdZRtIfvY0U5M15C2YeOBaz8oIupK7UexRydifAicLUjCgP2KZV4q1L0VY3RyAe77l+yX+H
xz6K3Iv0mW+zGFd4eqchmMdz3xhgnzJrrK+MwXDmJDNODGGk9McxzXJU8NQ5aviEEEWEnmYPMLAA
tO0XzjEPuqrVapyBFegONC7XLiZKWHl16sNIPpgTWitY2CpFOJOSPAWmaBaZmzk7K4UphQY3sdY/
nFZ+m5OfMoRRbrhWgv3mnDQxC1Q2qZSMvPRUbTzrnujKGXm5KAJ8dsSEkaDhDOVHMGpQMP4sTqPl
1aQP+PzsY3y5mveIrt3aw6/AqyUd8h47Fbxmhuytnwbzjvn+ZPYT4Tlky1OmENwZO0Ul3+weFujy
qQjJNfgVCg4zoZrNYnVS9J7fOjpc+dzT4bbceFn38FNwrY/vQoX6fJBmqfSvrci6FqI4Ci/alYeL
7YF2UMqwuKn5J4OV+LV5LPhwybhlbbN9I+MhF97PwLUQX9peDQLmJ74EY6q1gDdSxWxcfVfvLwyI
kLRN6iX+hdCf3WlgyQFStTts5eE6OeUReX4Ub9ubImjz94ZwzUmQXOd9qRYGLw+qSGOQ25T91mRk
TDupljwB9ifhDpyfR71rfarfpRxj2okSibSFLDtvKwl8ZDwH/G6TXozVxiBJk5taGrOlwjXteyl9
9OCUD1klM6SpYQNqVHpcVwRj6iujTOJFQc96Lyhcf7BfGTJieKV4lq/FI6XpNoY+H+D/WdHllcj+
kFw7t1jl0mW6r1zN6TPfFYp3ZYVXspNbbXJTBpQPJrWJZDSrX1yKGbvVScCZljwiZ3vxBp1lrsuY
otyhpDAaW0ZccFPSzn1GkB2SG2XIQCD9rbM5PBJ5gsJvOswuV9i3dyFOyk5qPWPcb8jmltQcnJ0S
58Cz1DyBa5Vjoj+rz9uNMpcviTZbFXs+WvtETJUFdWfX9lO/77st2wpygPTC9UNdltg1bhCZE+ut
PZ7djRQH+J0ZUMGmOGCp8oZ22k+o3Np00Wc7HzydI9KmovaPnfsGwgZx2IFDPdPiuhX3d3ohRhFh
odplWznwbPBbaTBlBwH2nAfpbm0O+ZpmzEoPn+iOMKbF+p0S4Z9mlis7TU5xB/Tx5Rtm7Sw1HcZs
Zb3hGO2wugwoW9838mtAPHt4tzvPFlfdMzmm07WdQaPSbjSRh56l18uapGV/gKNt1yd9xGFLRTk9
5h6fj4NzhD/mUVAjnlHyuC8x7DG4tBJUjFbCcpiNYcJecJ8yhm/uf3ngICzylXEDsok1GYJwumB1
d/hkmtJTbeT2ojGqEDwB4L9CXGuZh0SiIalsjX9iNR5JYb5cB2KnH+PF4TI/uG8i/vNRy1yGlUNU
NhRWRw2pSouIgWjxTPQmERLTcuPPZbhXJ/ytfg3r4u5KMSZhJ9fMD5icBXB4ulg+jk3ryvVE8pcN
l73xLLnI6DAKn9q72LGH3gdRT6O0xXwNZwbkHcrqRGrJZ7Hdezy9H5c7t/jetDJD8NdYChzonhUa
iFClqq2k217X3nDBjodW7lBLGx+ylQDOocIaARMCtqR4T1+u+WR9M/aoIVXGZi4KEpeoDWPPtH9o
bdKhEv3RLfSZAIBnyKBrGHnwRnfbIYfT9g38+zydMj4zdoTMxtB8fW5km09JQf6CfhR2jrGSy6FT
z317Bst1XuVas6BJL9CLDi9dJBY6PCAzyRyUI3wzZjtHPV6QBl3S6jvjtGnDJW6m+N/s5QG6W9n6
LmE3lL8kuQUXY+PG7zGFPKXmE2Eg0XXD4dpSTLUvgoHPTEdZ1cKXQHBDkuyq84c5jVcwlzuSAv9J
NSz6BdErf77x+OM5kG/i9SYTH8wRRUKW+oapWCrQFMTXhAhx/EjLOpE/fRCf5wbZ3Q/+A7uTJBw3
oA2Rd+WYLf/9t6hXShbG9svPcPL2LB6nKfBqPuPcVFdgU0I0XlQL3bhwWabXzkoyBHyuivr6tP7T
0fcenG50ZncLLPCwHe4/tbfquXyn5xaZ9of3vbo8HHaao074Jek3aYGpfvp18Aoc5ozyyvZMmy2p
z/qVR/aITPNMtP+4/A8LfVxrKrksJMKeMXrCnFM785np6d+ycoLu0fe0q77x6hg8oNqW37jWDDCg
5XNjj+U4RaKxoScx1/80oo49wi/NlpC4l97DhcZO56/jE4xH+CNAWUfrLB8DQELuZ8ldpEkydKw1
5DQlEcLqMADeQgtdaz7FRY85Buz7NGqjYchqloP8zDPHC07D8Z1ABD/n5HonSSUK9zxz3hWyeY4x
NyRgULY28aFhNjLh5vhjFiMEF8sY5xu9FszvzDTy7JNSRectn3g3eZAOMOfnssRjAqlYmaQehjnA
FuwsdbXMshEtearaLbnT+hh6WAc3amAXf0b/JEQzREp44qGoebSYyKLXNxNsMx7C802yhfPg6I9o
x1rb7R28iTSV+rgNIrbNySH4lIVPyMKLu4wiGG8NnDvUxpE+G1zbrwF2jSeTae+EHDdFIwrxMHT3
Z+Gpj/rnV01jx6GV5gFEuYTIE/+eDSjvlinyM74JYjrFUEoreg2tN/o0RAJ+8qd2fD8dbzjHV5kz
L3OhAjwLYClmDFL71TsfL9UxAS9bsMWDw9QRrb7IMTsyjcXNMgan1WgkOZZpiHdr7Pi6t9sRIEtg
VOW6eUVzxXkSqeEhTVYtrLndQ/8HoSgefWEq5JJQJlhyQbv5O/6LfcakCqClPpRWX0Mj/4EFPhmN
RsQAz9gCmg7G2RgMA8CQhObUcQ+0yavPJGPv5cf2vjlb+PakKhI/siurFmu17r2+51Pnf4dH8pwx
U/xGyAQFZf8hEbXmAeWriErXAfeXUCIfbyIt1h5/xTCPpUM1Nl7VCspMryxLldLsjKKCVWoFXMmv
pdkLDxntlu3fdP90R4ss0Cvoz0gF1DbqQpnTbnOiAZoWaWBnTJB89o7+xRga2XDaV5IRdMezZu8c
uRPzPtab5VvJKJF34KAgooWvkhTO0ItkXnzWzopQ815BaeMViLOjEa8NZ8UQ7sJo9BEu9CCVlJNx
j/VXAty5nQsuK79IkJhXW9qFtukjuG5czeg02rlro6YBFSpCguA7xD2HgTi2h2/1oBrwlwcb0IeX
5/qpVNNxAgTsnDQ9/LmNrQS6+keXOAsWSnk7ktgTHjZDc4UfAt9lV+owqMnjRwnN04glaIb7H0ra
glE/LaYlLEGXxIbVts3IzZi5M7vYm5rytUrpa/jiKPjmaJXlrwGcvu/G5LfVbDNywIUlqv7W+Ph6
RppxxBu18Kp0Ic2ePTjoF/Aey58hIlecaQufzk/0D5iV5cKuOLSxG+uMmzXm//9VXLh0kaeh77lF
6Xa/zKp9q6soQjfrltZwCZ5HnBfvzEQTBA8TuWLGINaO6Mzxh1AgkvMU0aJ2alQRjNag6AwrdcDr
ajVAgFkV0TPzcOWJKZqO7A8E2OtV+wdGcbmXqEvaXevlbdIZTZryXIPj6mSNEI4DrrlPrKkcVxii
One8RiQSn9NM4vudJqcwVePD/Hz4WLYuuvpAnW5HRMfxu5a0hxPPTnyzRdaAysgnv6JDtdRQRg4M
xAj9qKU4sQBJGhj40eyca5BDinnJZfJWwl2uS6x3w19AcNRroZssOPWGzNJiakLoKwxeBwtAGBxC
AbcITTlYjFkLl/n/tIsgfbHnZkke7KfMx4fdrYKIUsy1fwlG86lj58BtLQRq++Hw5I7UGjTNQlf8
aZPb3ZNMXAGxJ3uMUO4yGhsmwFYQ2EFuJlAYrNxdRSuSDA5fTvBXVN1b9CEikcII6XRkm8Cg1/PE
JAL7uNHcWHDCMb6Bxqlm8sqHFO2Bio/9Ll6mqYMv4X4TRSCzkj+6D2RCorhmqhmLZ1QTOdWu81P7
BcPC+KjDcL+/luSOnpXo+NIPt6ABneGr7mj0orqbk3zquOieeQvU/jH5P9GNR82l3OfiRK4HJZI0
VKABDOQPtakn2FauoEZgsKtT2r1fVDyFOUOhXVRYGSuEMXqNL1Yw+zJOPIWjtdvyf6/X4xbLWO00
4N/tLYDSFapfinw0UM4g9qEOSabMvz1JkVF0bPAIIycRsdwjtj47I+dKIvAhe9oV93bFt4SoN65e
IunALXEnIFuE6D0nERIR0qWvXY7jT2TPZOr+uMsMH0Ql8A1XZP2vsnSwv56qqfJzqy65BPGH9vZI
ev3M5/rvXnqsGGs55w0lb1tqwuDJ07zvpA2iepWYIvte4pJjK+OdMpSTfuUZMPRWauMIzTRi9ztc
5xfO+ezcNIgJPXWWxZcBpwyzfAz9CJ5iz2u5ySis46wQR3MOOR5bvLw7m6W2bC5yZ3+VbLGSAIaX
2WYx2vapMsUxvPX4DDEdY86jsh620ZgUQQWcszVml8owLgxfhmZ/gLgi+c5GY+z+SBWIwg86+lrF
30zYZtH8XDfm793khuKFoGwKX6CmUA6zJwhvIc0sgUUG7bvp2XcnQg9pw6w45UPoduVoYjLlqFDU
bVi80NkdH5AFxi3uxChpwBMHYvMBfCpRgrY/k1cT3W/5IG5Vc413rIBuVhKd5fsXu2mitOSzTwjs
x6vz2ZZWOMQdox2ZSfANfreZ5bPhgviV5eDra+gMGeVitLr8yOctOgME7i1+vqA68j9QlKNnOPkf
VK7roI2GvYxtHWwTjgnUOLZsJ4ixUSiJmdEWo665MSc6tkrJUZKRHH9pryZfiSxTTKw95BFwwr2Q
0aPUUTOyTOtlE0E0y0BHmncI/axjxFKyKXJKuE8uEgN6RebBhjNnoe6PySn3xlD0/iLlRNWdMyUl
nW2vRtZmbI/UyFfoPAia/DP9uleXCd5X0WiTBm0wwb7p9rHfsswK6KimNhG8MIU/YQQ8zeHunMWQ
+ALgTly3lg9lwV8NtfBqnvBbhNyj3h2E6Vk0z0qnnbsMhDRNTBnY/rlp2O6pVIKBnGUBQeLA9OVJ
zs7WN9yRu68EDcxUWnwJAH2in5zQiehpEs2XtN8Oqn2t9ub80Rg1BEFop2Rzo/4uZziveWB8EEKZ
IvTKyErECvl6RS8mWYaVtDrNfl0FU80ZsLn0ikl7LGUkQ/TdbOW9/SVollrcjX9BOag5/u35uJr8
UnV8RAs01s7CBf7/UUnUROiylPPIMMK2DQZtFoa+R/WV0ieyuFBTSfA1MLzNbhNOfRqlT5gmChu/
Rgk0ukLvPpwko6T4FdT9FC/9frv2tfRP3zBIXvzippOdx6ELdFHQqYl93YsI6JH8xP4z1K+8+Xvk
IadazYon6/VDpNamGRxTNo74A2E2fHI4CJVbtkLTh7AAyxyK4WH5qrfUU5w3Iuas6u1Oc2B+s4M1
unE4McxTF9lDLsDxvImFCrkGfcyfVxcvYf7SJ0pPAkqmk4lQf2aH7FTKW/kcS2VyGwQ3pMRa3bH9
GrWC/XgRsZK5mtVqPsMXBDXWYCOzFn/XEhdSSaXlUCkryP+/AMqBOZrh/gIESjdPofe7RkKA2quW
a3fRVamGDtxWPPfZ1B382s+J66Gll/3lJmZgFuX9Vvpmiv5CRKca9GyTUWhp3q44TAUzV0o3GiZX
qohFLBTeL8A82JN76wZWWylXL6OU8dq7haSUgHelVZieXboIhhSZH7tLlsOFFbeD5ZSQXIhWQJJk
ccJvUlrkBmT2GnBrwk4mzGng2rvEmBW7kI5N+tr6GrMLlgOScDDCuScdLHhrtAxEfOK1Jcx2MeXi
6xvyH0FEReuOkDpXxBs2AdTg5HubbtY1gBApsVrWMJb/evniF8rFg3fvsWhkNHUA44/otPIdzuHY
4NqBbgpAm0nQEqId6c93m885KOpdZUxJZT/u8nkhKL4XcKp8zPk9isJdCD9k2vmZZTxraMaNOj98
UI5dpmHfuYJiSz8Pl2gS9CEo5nYGZmxHRxLnRcJGekM0XA6F4H2qRHRpNd0OVDcPIN7bY4QSZQP8
rRD23jXvqwvGVeGNEAp2mS6ffBhCNWDePoQ1SByFdx3JQ+tEKFHWhGK/p+MeJ4uBXSATXxSAO5xP
PLOzKLUPLIK1TKzpHGQk+LRaF10qE89jqWXiveQu0H49eYy0syJ8qcnctXRYmJE7G+Mhc9Fvmuk2
8UqE5VGSMCJz34P2O26i26VuSy3FPaHNtFnh373e2lqmPKblLAq0FkoaBh3Qx4NXVQGJgq4JHiA9
WgC9c8/eyGDiYJILEukNVijVXwBBe2GALcZooipGA9Lj0Fus7FE588QEsKskjpFgqgMVyMuE6FZx
4nm4B4rAiVgElRBia8pafjcLPf4vcZDUOaJd/2wk6J8GeiOOf+8q9fWvcOeLr65KsjprONSVSeBd
zaUnVVvwjF9H9RLVmQT+NM3SEmTjbq/B08efGNCYD2QN7tf1JhahJr8e0tXRfLZxU0m1w/G+6+4d
grI5M+bOD8vFKzW5zUyNMeqISrVjcC8LAIvu2GJp49GJeGOYdGnqLfTONJKc3FbHDWCGWWmwHknK
i21qd0U96Q3arWKyZAx+kdiQl90IxgNmevFO1/sDFRwcso66fNOUSkcohvcXyX73qVP8VfszAXLa
zolXeOdXvsZDUHXZH1g8nemeKWfB987VwMfGNVcmA05hx7N5M4o101v1Yt8QBUYpviGI9Ijv+V6E
OHH3XmHHVGTfXJjgPNzKC+T6U7vQRlk7fluNe/Wdrbr1goLqoGxngAAjNvgqLOVPGXHJBGXY6Xh/
4mzqZ7S+pFRIyw7lAEUcsKx6mD0+sKUhDj5oM5RPnBMEifWPGcnbPnHdrX0YjFDODzvnHoyq1e2z
we8E5qrpVFWX7rzb1aNxiqCIqjrKAC0QqBUUXtSdWD46yikyGvj+1idMDJJpXW8zotElCIZdURRR
RnHeKC+J7fQcnYqMNDGRxs5YET1TVN2sJ9Gar0RFnNJIGhHTg+Jn0W+mLTmrRWjWZbcrX042U0kl
L7lNgw/UwkhZEmQhGy8svWTZ84roidN7AzmLFBoVSRM+E/kdQVf8QS3HA9dHUm7KGtaNGk0OZZ6n
UhoUV21TO8ymMGD9yqgGduQRPclvHwnImCgCpUJQBMoxWTHiMRxI6C0kGathKNPWnQvGkX2sSTBZ
WU+4VE1zdV/NMkfBGBlpJoTavglmk3GLQsdx9RbW4t59Rd0JWy+AbI0Ge6dkxDgIBZgkeqkhwo43
bZ+ToV6AD3oGWAame222u8jRZkaOzrQwrzVc1g0z/Awi2dH/ozYJtrVTaiYthkrIHS1g/nbGqbxN
eLYuYAVEX8jIlCTQZvgJRbmORie95RnTcN0Hpp7EmGu+UweVVJaXXrvG8DcpNvKfajlo3i7MsnVB
++wCN4hu3Z2qppSajCHyO/MbUXQXZtRpFuHIKKCbHVLWuHl11nucjsr4v4KWuJk2BU3qocdXKHZ8
xe6nwHnwTMDDjdv4++pcfK3MSzt8gtMcRfH7nplSa6HCTix9e+BcBxkz6whbdIG1Z0r0WeIpPqO6
7igNjdFE//x4vgJDQicGiBqLd7CArRf2cnqwB334hUFnSWEStX8Bn2G2/5n54tOo/Cf4I6zEqijv
66t+W9dHC3mUASw9nHLPgGcrdrDimr7Ani1NJE4Fs25NNreY3VE3JmCxGV5J1ZUH0a0+ddKp73WI
TU0MKXOCdBa1/vL5Rx3w2Y12RBkwvU7xdjzS0LF9Sl7C25/8R29Qn/pSv5K0ohAd1yqTJeSAW7Fd
p/OzQdWEPZdgs5mLDfJDXXanfNtqoCNn4F3NxHXf8VgNeyERy9Cxxdxc+Z09UrksqioS+mwUFBlC
oCxD7qj8t0RUCy/aFg6P3RkJtKfwJYFKUi2zMpeclHQN20WGNQZknHZwq3HSh9WUZc+cIt0RBkXr
XFXcoWxNo/UVwVpb/bCRtQAlFrCCNmI/FEIj37FOlyPNkpLA10LRpoaDme2/b0zgllNwI+bnHnL/
lq0cEY1kFNzYxPoKAuXo2nsZxlwLvRLSvD8/bpeiXjysk6mIVB4lKv07TNQXqqoi/cAimUjHEixi
HX14Fth+f6jwWSBTRasOboI1yhYWQq2J0i7j2k0g6FGQwW51mN1AZsax6cyZmZq4xK7Z+KUQRjnj
J8EzrjLWKMt7t0/bs+iXwBr7tTYRe1psI846Vd1hxXuJsL+YBjd7+bBmXcFeFfIVO6lB5/oBsYsG
91N8tD8e1sIl5WukO1OlsE/0H7zJA9OKsf6jZ0AG4Gn4oXfsiCQVYfrp5uONyzVIxXnStYszATQA
ywVBMIoabDijPmCeM1aQXm+c3pNhsUOYlXvskk51AksgIGrCUlCFP3iu4Fffh5kGh6WbH/9IJuxs
dJ47uGwWXM9zJGs7hzRqH05ylU1KCrIIJRcAZCg21fYUtvdVUO4SXNgSlbJ5/+V3CmqUM+GbPWQ2
/MZd2gYusAO9gxe9QsCcOtPY0BQwMU0iT89H0PbMh6m6m6KOb63LnwsCGy29rmBueGp8NU1s84py
SFOSE1CUxWbgmxmv/8pCFhafmKaH/SPDTPGcbR37Da4TPmXllf1mW11oYDD6YG+DNWYmk9J9S3JL
ZhGyZdD8kCzpm4cWrFc2F5zEW8FJMrCuo10KKCIUDjdMtl0elLES+zzBoxHpVUqSfl4TT9ozneJN
y7y0DKFvjcxiHCb6swOSY8uOG9SwRru8zoC16pfX7ncnzWDi6H/qS1C136c8pydJG39QHNC5rwxk
pV8IrzRQbDocGCkOnD5ZGhL7uYzPp/sy+fcqhMnlNAxR9KN3gbmH2qUIJtVdvAZC7moxRnUet2Y9
hQ+MxWX3SZ7v9hynzFOtucA5hXkmn856Xqh3R6RXY3RoVsPTUf4rTna7k98+u7qIWu4oSClypYgE
Z8CxqfS1jQB3g+Mw1XdjZu/VG8G9bzFygQ/NL9wG+ovxZFfHRtM9S+WfsdxpVgayPqF+9khoSvt2
CeYRXnDvg8Pn5pVyP0ysVgDLkIEjga2416tFIZpVGvHgDNuXjPrxNWmcheiBLzxyWjG1kZyK/sn5
aGdVsa2BNMLnGDsJh/Fvowjj/XfFVpnEg/OIT9lioMmmwne8SX3gqa4uGYMMa6fHn+AGQXGiYsRn
Uh6EzrZ657JYfks6od11arnToPKH+6GxR0yOphYqNXxQpLjMRrm1sSbnCyFJ6t8/LeuJVxXxjONy
k3nDEXx7Md+3pWmlq/r3ROhkmogveRnkE1SM4pDOCIAcKe/Ats80wWOf5n3yTGDORGOmb8m998Oy
fHs/eyt51XDfYHp+pWOhpcrGDBiJNa/xqsE0N2rNvExH9vleDpe6OWiQnBAdlrX38uCWuXko83xv
+0sCu1mmZYdyvRZZDhsYECEAH46DIIrVCeJWteKptuhQJYVEiX05hAgiKM3KMoMlRLkz7XiItyoz
Yjni0Ua4lbFoZRKUBPxt/J760dM6PFlnK1fwEbFDOZWaHVmLDTw9n7ywMpaPabIcYlY+iYORZyvJ
NWYm3l8MvuDv3Bq1dXeXmVTo2I4Xo/AvqWPn70PH+ieYnCA9sf32gQ8KKgjmZv4MfUeMC4Rrca32
oGRju4lFrBZV3HhdXlrqRHMpOlmr7KUZqKVk7Q4eKFpjy3EkyTy65gd36dTN3LUGt3DRJTfCxvXT
MEIdBjX9HMaYD7wn2o01+7LwxUrjeo53aUa4sN3U8G8CzBxQWMmFZqoT0fluRkf/6fY7mgp35hmZ
ysykKP80a5ePGSfqCgVujh243NE+9uifc08GMlBFZElllLLviFkZ6xhxC7wpDF7SO/eR1ftT02P2
mQWevXYtGzf6SVh4I/zkdZA6bXkKKTWSdXuekl7h4nu7yNOMD55+fj2r7/VWI635S6zQWpjnezWl
seAkIDoExi3n6Lqp/JhpFWuilbIimaKZ11v7zYs0lc59FXSaAf3y3VblU9m7qgVwm5/ooecJYEPl
2qRtt2/hC3qFyQTyo7TNtXyW3zxbCsm1p9jtPEcFU5fxmIrN/tPyI3cPKa9w82MoeU79Y9NrUSj4
bRmiUJ8HZOJKKhkgHnohbBLYlJJg9tOnbqGtVddOeMB4y6iWZfN68vqZ1WHkVs/5UNuynk5w5MF0
D0Jbrt7qAGIg29HtUGQ04r3c3nC+lyvrRAX+Uux6Dw16h9ZNAABHg1fXhUdiCk9FTGVEuVmCYbps
xJqUn1Msl7lQkwEeGHEUucfZeDG5is4kSneANrCV4UctE3kFtg2IvMnZlen59rBHT8iFsgYCmKQR
QNIHbl3cgW0IMdLckqynDtBiNTeb/DQpd7LGltLg9GAUbPE2cZpsgU4pe1weeWAaC0jjdyI5S6WG
8Vv0uJYGP8tqY2fF5fM8e/PeteiM1/NY7nQLh1JenD7Gn2JMtXWof58VqlXJTq2rhNgoe2DOszg3
OypjiiDgsyrT2g0bEbyISbMrnvvaXAdUbPkJKRVlyXr4CdoHD/aEfE/9ratxoDsq+9gZF0cdvOti
1cn2AHe2PxeyGAYSC8w+ijRWcV+PKUzIivs5FELmpyIaSaPpg4cUJ2A8XDF1wPGa0NesKTouKgH8
ay3/CWc3SWtQ+tOVn1H4mqnp9UH2WllkDcYevsmXu5yZasrsNuX6GMAReUiWoERHqXuggcGFvpW2
seI4NPJnXm2q8Hzul1HxVamrAbK8i8SK+Sj61H66Q/zLtisZpLsiPAZ6ju+9F6HbaUZPgYy9p11a
YnYPxU3svtA1ScqkJPz/KlhGaaijION7ecoT6LDFd8pBcjoDqV0jwuhFoegGlZfKswe+h9x9we/4
ecSYvLq5OvxLZ9kG4YOW0V8+Q6hYTwhBC96YlMt9ZYis/IDLF2SaNfLdoujGmiJP4AB2Z0VNvlaH
6At5URSXJ3wrF3RtngzGWbDyX4tsC4Q7IqTkRDqetFpzlqQVtG+7mNf+Wyw5hoWpwix/qFA3LOxe
BJ9wMaL7WVsILUVm4lJ/taLoWZglt8heqoZnLFX3hmGkYt9qQTtd+YtTJs7pDN64Z3dtKSQNQdi8
eB9HgN11n/NJAFmolBLYGntyumekO7ty8eyCyD2H5VQtr6ks69rnXmPhENXmtiC/E1F+ihYnhLUt
n4M4Pr8gIoFoeOTw/Y29CV31VXdw4hIY+MYhLDlkRDSo22H3LGWg4j+vsYbB0ziayeJdgnyAfQEQ
fFxAlTDndjX7bjUSEWelC0lW7XZJqUwK3UaSOx2HVC7gUwbyp5MnBLHvRTgkpzI9zwMHfPVJ8mMU
iazr0wsKsRWOCs/y3nGckut1669bzWLIU9d2Q2yBSSmn9aad0zhe2zAANE9H+OnTxSpW9aTxhWPT
GknTo2PPxGCwzLHIoyaSNiVDrmUr+lhwnsVfKBBtA1ZDO76tbQChN3u91925gvq1eSqYIi5ZzHeT
2BdFQ52uufnEEgXZIvyYUYGliKIJLAN7Vf0Xh11zalisrkVnbWfpHX0rzPX4toq0wZDrRuwWZvLj
0yv8r5XoOvH+oVpoCKybeQTSaCK0dfpjoENPaQCtNlyWMvAL4/bFo3U17J1V5SsCihXR9nb3QjB0
zKBK3AXgUpitWqKIQp/OkgfrNLUFJl2sa0E7izaI8EG+aBr89ELE8tAHT5FxR/4RDyOIdOnIpVr8
zBWzn7d1ZymrgXC6CHhMcOkSVEnOug9+lc36m35EDQOEsFty10Phk/e+ow++b0jPUT58VeUQIk/v
lJbQkoNqxSJ0iD0WvB/uO1m1AuoZe0jo7rU+wi18ObZqv+6fQj1AQwVEDj8Zp/GoTZH0/KmvoBNQ
0aiYMPFnrhgm9tdNj2X3GifxoViItNwdZBxWPqWL7bsFe/SzR0LZflpWkEIrH/1AhByj8ufGax31
42mSr3UHw5uaCcaARTRbyGa3KJ27jZPrXtT71QDGkBytNe/Y3LBoI1/uwoVihZJ7GGlfotFg3dC5
ZFR05DIujeotTptNYxXrPVDu1H9yOE5U4in0r9wyE4PlrrAQ6lywk8S/LoUAqynfvQaN88z+QegY
emtR8JsOzCb1UY7lccQ+NvHw6oAEgDvDM22WQrC/zKRAQ1S4y2E4TpimSpGQe1GMshrq1E3YdCUV
rOv57HgMgOlwK4w/98EaLqUgu5mPgozXiTZngNToh98aWqzIIwpvAP4aQpHrTjNWkZFE0LstxOhX
KHyYdgCp8YUjeJel1sX/RlZXLXfF1RPLeVmn1/dv75vL33E8+2LgwgQgbbIYQ1ic0rmX6D4adCHl
wvVuX4ToMnGinMb3sz04pWQQVuFPE7u69hkGl6AAhRJTQpbT9Nd96yKfA9eLlW3ymtz5bE7iKlxV
lvpRr7JMzsKGSneAJyqRqh+6l32aPhYs7LX8yqQ/mbkDZJFhzNbCNbztVtBrXFC5OCppAwklTThy
3E4dk5VEIjZZEQ81ViJqBInGlvOmtwm5CcneplddAK9aZWoN8XJJNd7WkXXFEmKtJ8HIupzzyd/K
ZfM9AbDcFW7qlTyLWYNMyejYPk1Z1+QJnL9zM6JyMEfpJtm6FrbLmk2KpUvJpj3cfuDeR8X+nLkP
iYaT3zD2wUEFqUSYnhFBCML0vM8eEf6xFemRORgiPIPGDHsCKzplzd0jeHzsBzrkz3Md+0nobFyf
9y0ij4zcxbV+OMKO71QcnF/qGpS/JRMP1aOam/fIBUBX8F88n7+kqebR/v4pvq18gGQHmJLimFQT
y5V1ql6M6wP45ECgeOoBtmftPQG4+38nqdV8qBlI8RH/HuQYX5wq5X+dkwdu1T6LxuMDuslR1Zof
rNMZcdOGepGl7gEuF9bmO/wL8d5T2Ro2LUux+DZwm+c136xj4PkY3i7UH+e68QUfw462kCi9KVHn
UeyURU+junswXQbzkXD65n5lRhQ0o23Kf7nfQ3qcsGujWBF+EC52WrL2wwUA3ZUq0xPJrZ0bGlTD
LEiiuE/sTsWVMnTshQfBZ8gQ1nsRDFfdrEm7sjzBiPZb6kKLaDNHLEWX2I63bwMq9EeiyAoUQIfq
Rnixl3GKi4+NY1mjTCzzgjIgzO0W1PwGAHPJmLOsr91soO9h8rkFO7Q7IyrIKmNHpWAgP9NlqrHw
ojR19F+SqTRlme3xolNCFn98okgeHrmqGLmPzNE76P0MrTGillAornmQI0TEMbyYyljptVIBOFDO
LZpd323Sdw2SzlODUOP4wvF7U1gNRL4NYtA5KGYq0+LZGy2R0Fq03UmqXzgBQcYXHkkh5/c+Fkuc
jGg11nwLEQlaDDX1I5deIDKGS7R4DD2PtJ1wx6DYRO5t8ZoXcfbKQ1gUG4CZXzTAKCEy0ctqChkE
lgabiWFJqt8Jl8r1wt6jPj0tajNKXzBkzTf66Wz5a9cX/CVdCec9v/DBt4k6j42cNX8Xg7SvzOrs
HsM2dk92OOZwFSs9kIzdOj+EoQdKDrybfrhlndIgSWuKj2P2d62qpFgiT6iUxujrq0HkyDEGtAtt
liyJ1xCcGwdjR7I16VhvXgGo54gltlqC2q+RJBeEW5Y4EeEFetxScrcIrn1p5g3nVHx56Fe+9/rP
nnGeYVekwc4Bkl4j6XTERfFQTh64EJDdxwEYT61xHbubX4VUbqLtasvee9RqNBI+PjIq97M2W7BR
0RLd0zMy+G1KP3a8MGOUlCy0ekKZOitMi2pK0CXy9XG+xFom1qx7wmP42qOJmt1+x+tKynRSspKD
Rrv8nDFKriwowKpLa9p94cozKqPm48PpqEVkV7Hv+PtSCBL//dr2qKzSyo/lAqFF2dS9h8y7OmL1
0nu5p6bc7B2TUAdXcxWai1KcVWu9kchOMRSDO2IaMlkam2alpkSr3E9TfECyTDYjNyppF4GEcsdK
m8A9l0GDP4HS7fibiZQKkq1IGidk1JMEebHKH9eLNTXRc15rT4zHVKEoi9E1uHdotVqEdevOu3k1
9ViqNVm6gAjohrVq7s1jz9x65h/oR9Xf/t6dGc42tYwyA+U5hYBgDn4LWTZC6Wbi4m6qcqk8ZWqP
ivu2NKYkADKCRqf4mpmRwEZeZnM8P4wbK7VYdgp8ivM91ggF+N/ECsxLJqApp0vewB2FRzd4fWFg
WhIab5cGeUEblZy9GNHLQYPH01pRpyUsUZBWtMA7XRZUYI5Bc88nMi2lu2rkplX+PO1y5yi4/PPh
+3gdNSnM/X78M2T9AvN0x721RPuO1UojvqVwOL/MsFBdDLmGSE9+nFHl58S+fHNL0uI3cGzkey2W
km49JG/SWh8RmT/vkFuECdP/mgy9/cLGW8CJBEcgvzzDqBT/Y5SDXtuiKLZ20p3htoQG18td8r+X
XuAQdUmXNAuucNMOYLhUqqA2L3d2kuMHPETMTcLzKiu3YqCDs0hTbmXdu+mxkhSxWrqs0pp8/vh8
etb2UHiNb9O7jBeUO2XikAOmhzxvWTDenxKBN+QWEg9Ot5T8y+2izubaNByxkLCiyhbDkz0b5NBx
BIzWw5AR0fRvwcpYszbYLlYMEM8cc50ozHmGFXgqQVL3fRhhAiPywPqM/AO2wZWOGk0vCvLI4hEP
o7GHJFi+dWhNZ/FtZHuDE+I2strxMIskYFVOLit6NbbUj3qiGoXrKn4Z/k3neAYDzt6gk0jEm7zC
Vd5c42gIInAszhDIIgVA69NNY4/PS7KZab5GLqn0N6ckjjnUk8I7zRDhEF+CgsO+oaEQ2wxauQFF
W7fDjfO6RTlcJMJy5IRqkE3EXfgC+NVyp19MD2Rd+0RnRGTBsYXc8qSGN/osQS++Jq3q0VZHxts8
sHj8GDvJw2hIow85S5eG4qjqYK3dWwg25CAkxRcS9Y0nIfMXXRrCakfYCJqdhvPEC3AsgWg1MFxC
fnQ9EH70J3ZBi2V24hmmwTLCV8unFXwvixf99VB0cgH33zzsM/fPSkhf7rHXrXDz++neBp4avKyY
K0xxc93nGaxF8qKf0UeF7byoNTGHuLRFsZaqGWEupF0JCL9a3PCAuRZXGaC0DKqO6DAMjg3KIDSC
ZwhJ2JfTHJaKyqeOsWlUze/xZ3TCLXxnV94PKfFJ89cH9gt0NkEk8Eq5tAcktMkqbZxOrV9t5I9F
XcKrXj8UzhZx3EVtZ7OhI7ZKJZrqALywY37d8mh0yCqcQS0fwKltA3clKTsaOpqQOVKF47zcryi2
w3tAs20N0wsyZ6+PkNSgNv06yNgnnkyG7b/z350CqCIn51Qli2M66sw7xFaCNeNt6e7sRVbVZvpL
dtf8GqiDn027ALsy2x9V1qlBBYZl8AC1ZVB19Cm7zndUQj1wWLDi66s9E7RgHANR5axxqFEFjKbQ
B0NFRDcP34/2ECclbIFV9LZet524LqTZzS+dgiyi4jjt1Qy9jneQyhfEuM0n8NG3WVbY2vkwfXoF
sZQF6zwP/fRFdgeztktRvP9rhUpFYz8SHrXWzjVTYVYrWLSlp4yxyx+smYjhqyLGLwXujo8NmdMh
xiT2p151Ehm2xLphrWv/C1o9jveSShs3wkmFJ4deh4BZ1StQUZ3d7ijA4ndXUKO8UCozWCTQvmwm
GjOC/edw/RnRE1fJed4rEdcEb1wV5t1n3uZTU+RVAPnnUQpzf+JeyCRzTI9ljiEdpjIS6GYjV/+p
LBa/uad4L4VPDKrIrS3Q4SwdEkr3RXmZrpOj6RLYI8pZT72GkxUL8TQesgpN6Ige9usV2rPW5Tec
58kv7rptEq1mUJwT7kh7uHw5ATS3znilysqyuRn5BOCR5Ck8ZeZvRqtg9ueitBxORzoFAEEbbvXR
UYZrz6A7h6Y5HsfOWy/qexTEHV9PpZaslPosyhIIcqwfbRLbG+F0ifCSJ6ijR1Rx6f0EZ14PV2Ye
DpMXA1VbnGpC682vGLwFGUg2mauXQzsKXE9Muw/wrfEtfvN9j5rzsgxnlxJiBnHzEEec1or6NxcQ
RIhDwZlZD8u9utR32C4xq835hy/Lkr4r6nUzi9XEGEe18lPZMR+xblVnsqlETuzajnzxHgHhJpL/
Op/9EDD0DD2XFxCOn6jYd5P8H+lyLnYPEU1p3kgHIjCUAqCS+WDW9CK/sPqM63b1FAljCSJC40Bk
l+E0sUKwLA+CYVpmnPYHxnZNe8afDLXGF+Qy9LZYz0pkP4f6i5oO4RoyYmHbRllrjrZ54MpR+NOl
zY0jVkyhcEWvjU3K+ncGrfToQM40GntLc667dXdJhFcp6tZldObrHVcwNaSg75fg4X1a53Frvn8Z
pVTMEU3pqypL5eDoqGZXvkmH9wAc65Xm8LziOeXzgEY+ksI8frQ5fGLTqCSe8MD7zUcBmz2EowYv
uyK4BT43ylvU+6NUpFfO/3hkkphYz2/e3o0YcEb7ob6vWAlDh18NAvmNdzXALNzgWKLEcL8wWpsq
M65Uik6zlrF3Ii+AU7DLdFgyYxz2aotgH8sM3V+KRTLlWwtOBpJWGFD4bwyXQTwhtG1wzlVVevTc
1Qjz31UH2vzyUJnN9pov1z73xm3sDMMI404hbc2+9guSZ3AupnZYGU9DjfD0/PZEmx7lkWTeVMYH
gnfmf+FIf8RtAXyPT0URMiRcK/5XrDRSQ+E4x4BOH2n1bfD4LBW6OX4FdtF5mh95s9JwlYYykt3j
7EXfwA7mThPg/Xt+FtIjNkMJB3ERig7vaahF220LSCZU3mskXjGQt+4C2XE57eyt8ThB2BMJtiue
vU0Wog0tzE+84OmZLI5wgiqkNd6J1Tjt15xa7l8lQDPVxcZM9wtVI7LlHUrsTpmf9b5hXPQIpArq
YQ7+u88C8IV1Qfjbcmx6z/v+wNx9J0ra2iVO0LiL1rWTc6ilZmUabZs7r2cOi387GmSvA3tXUNSt
14Fo0nui2qgWqPEZYv4PxhFgyuzkMANVgFeTnZKr4Kw6zSoLYJuQLzt1PE72OxRKZpsGiutF3/FN
YLtkxI+mjnAbSwaLArPxK5Cn7txqz68HizNLIwzgf2FIZ9iuuh03KUIeA325FtyOBAADRLrXtLhw
USV3gqsAFz9p25mKZsDqxi4HnUvXAYAKHl1HAGYawXp8nqUCltxQrHmMRm0vDEQyc8dlkMf7lPQI
CZUFgRZuNVz6+s6Pko+NPTPUSpdQhvBNltDJUsoE3zB8bUzjxDS80x5mSUMRlSCVi+AtOSfY3bFp
eMpd+x+zfnGgm5CG4hU8UHsEiL/yPb00ujeCqPgVXUxsIWsUn1k/+2K+kzZ3kUF1/amlV3szlXun
wJoudX7jJtpqKWnPLJsT2JtMiKuJo49hvkGLNgUUNxhiaaEbkedVraSBgiq0+0/JZ0IICx4dXx2r
6kBYPcSgca69x6V1/ePfQ/5oWsUL5npIFvAqrag3Ch2IvTuzcGkJUYyOjCJjeYw4pK3CRKbscT8a
1vAGpc5TyhThCtyb7mnUr67TztkJyrVkEP5ta+nr67dUa/1sxgfacCBQBa8eHjVqZT37zAE1NbYB
fUaKX1LLfDqrZM2OEfJloB/BMYfPOZDM2DT8xvIOr1Whq0eZezpiKFsBug9CD/7MWPRVwAPY8a/h
XiP3xqnlr42t7bTdVKIqbuQBBwI3CjwESRP5U6+XjB+l9ay/RwXeYht6PNFRTU085QXuaVmvq7ik
46YawPcSgRn4W8YvTEBhcmbuXcEStiN+f/oaPYBzK1J00eRgcj4Atl+0m+hyNZCNExUC1iDcHiJH
XZwB7QPHRDIuRHX4J/UZKhqsfsLz53OS5WbNgHVw8zShhGbud/fxgb0fhuZlLyC61kye61yYAued
Gwi0IX8sEh7aU90mxX4njLe1Sdmu50uM4JzIrBybOeReth4hvhgaCkRiBMHQ5ja81ciEYAm0ohZt
tNNiXApaMpNUAmPFhYh0lYqwkCuliGqsCh4dodZevh4Tyd569pGrEnPvZM0LWy9cugNJt38dbvFR
MxObxb+CamfD1GcOKQlfeU0uX7g9WFoL5hDcJwlXIZlWplKZ8Gb91JE5KTfAM5qpAXlSKo0FqSBZ
5o33uyT2C4BMZH7vYOK5cRfQ2xoHQM6bs6T6t6MdlLSyPsxf4rGHz8vb2g3fpTV5ZUSSy7vqE61j
idB+dXIDMUy7X//o0XK7if7s+y9e7AEGr9s6at5Ifeh4rTGdjlh05BZg6vSj3IYmHNE+ZR0M953Q
bctzqjOH1qDH8/esLlu5G8Wln4LlCKjXFYGcNsGUS9TxSIld4MugiDnkMwE4sPByF0T6adfeKH9i
e8zA/GqYBCvEiaCVEd7K+DT2Y0LHpv5EsapzKQm3UmgbR4tJAe+9shYwYguy+Mc0MnauS6l3ARDj
xei6/F58vUzCu7IrNQj+/UB1B5oiBOFxYwvEp0ZxYV6Hf9Ad9b9DKkf8GNweI9J599zC8gHG0YMa
oiR3NgtK9KH8nUMwWpr6/5JwMns1YoOJWbWkTh3pr2/0qHbVqywHmdDMo3Z7CrcWYO7btD0UDFDM
gx7ZGOx3SDNLp3/xi2en6kJymNyS7YnDj0gdZ7+ibxGY3BOlwIPe+xhY83K/ESFFLprlezV+VuSB
rCJ/mR01FjmK97PzQzzVpKO4iKo3TKIUGbM82X40cc6NDKrVHETlQvz2oT4CSLETevXR6LNGZ4E5
Crz7qb56ejK0sArUzgKSnqiESdsdotd0DyWI2G07oFiVuhhUec5MYWQWY0mITQbsijZ1la5oHyl9
MW/TYUmmVvZzjAlNfC4Vqm8X/KozMlu9LXezibWBF1m7dkSlC2ziHDRf30m2Bd5OWd2Lya1eY3Ng
7SQ+7wl/6SAz6iJ6LEzEUrDYeeW3b1VuSAjrNICUbYsHRv3DqHzEV5/gr05cMHFqNV6z7ynt7P+4
TgR0Mfjgi0x85JgBA0T9NLtDdssgZuRuELtIYNOmVLqo8p6XxJTinmi2Pn62GQBlTMzxMukoZnEb
nXvZtUHmZ1Vbs07eaPVozDVOp6i1cW4xyu1KWm/y9mVixLrj+2o8CpnvLPurmFtEny2ogVk2mBlW
edmD6XRfXahyEaUaPEfiNpK1Z//neV2CFlk6tzxfsSzBzi7Yn8DrrGV1ngrlLvbm/kSY5yUWLEw8
jK+IcNbfqijKiTg3DOdT9wIKxxQp+LgSKCoqtmh8qAZZsGwkWuoySht2kG6+t/JKI4bJIpXyiDj0
6TZ7ewg+2RnzgNrGJ67tdoBB/i5pGrO8w3CAXMP77frerh2I6Vc9+xmRnHnW25JHxAmy1S4rG2mu
w/pC40ShNSLX8nbwEYqp0Izg5IE5+hnxipwW4Ercmzxb+ixMjU8lzbH9VgosoPRqgDqDrNgRwNsN
mCN347ijobGw+W4vogmQ0Dp3q7+pyf99cnA4YOaFrILfHs6XMZ1SPt0nJe2pSvybBqMnlTf5fMqu
whcSAHnC8s0Cq53TxA6Lg3SYKQ7EdGlz8ml2cl6oJq3V0tiD6qGgRhNPAttgOMx2XDFOZcRZUEal
snnQOKxULobwMo12bd+ldigNCMCJeGwClGeZhUBeqxS7nmLho8KD1DhTqB7b7nxOSq36O14wqSyF
Kb80ZcOoNGH/rVIIrmetogmmKnCWdHq06z9ANZVVBRDEGZ5kdHPrxL0HswiN03xR1NYJDzyyMjSo
iTh5WgkfWejs1StWqdNu7N5K1wsSrlPdD0bZlifONIUpm5QnGOvv8hdULjulTapbozVdvtYfUYdW
pIgDL3D/9TgDIPCcWraGT08dXn1TE4Po9nVGIJfo/Rkr+DfRvzquujc0sYyJKwoMkTgA2vkadyCE
Ghs1VkM+S2FSKFJGL5B9ne9DNHmYpdKrtDUI4cMCmn6iRySOV4t7bXcgrvRqloe8WEKhbGvJdxjb
Km20XsxK1TkLkARs7MW6uZTWl7q75ic7iTocUJDs72ePA9KZ2JQjVupx0kMCWTiRQMocUk/s2sh8
OzpOytIHHNEDdiywHXHYRl9ExvRiWPwaibYruB4gf4NYHYQ5t3Ti6KCUYI5c0KwXLIwXBfjRuJjk
IXVyt39HpxeRC/s6tBYOh89Xsu4Blykg7ofSCIn6cXxvcdyI+ROM7A/3JFbYzL0hhrcsFKQP4eC9
PH9mQSeGxva1sCQNkfK70cv+WUKufsmT/2YR9wp782N1KuhRFmIpn+0WJzs9HsHwv5D4zZAVD9oo
Nblr31Anoo5bCzxjGXsyX28PFLoXtpI7krUcB0hL6xBf1mObxzU1twzIUi8tlVm+P/CMrM9s8ZO8
0Fi3zccvRmnJIozWljtIsckin9qXtGnEU1uKE8jp9zoHgq6YQqZfShM7QIDaY9iSIfSEGCgLOsJ6
hBHj5l9jFGkTbDCFgPlkT07ufK7bJdu7/Wrw9TR/0QQMgT1qziy2Vx+85mclTUYVgo4aBnPkzVuk
rJlWF8kzLVGz+YDiPfka+BKqFevLkbACKBACXFdOXOfTNOMFUw3gEfXXSVy5MeJAnjLAmbG8xj2f
D2zw9kyNFST5nreKDhdUi1F3dNnwiqFldOebKPyy3x9ItnLZbkRutopgAwXAA5qCYeOauYcL2L/8
+TPnmShZZcLsx67/8ByaKl3Jzl6JPwKvZYJ4FVAVePU/qfM7jPqSqF90B6eJ3XViAGuCU/vdpxzv
H7+MyirsaxmR50hPmFd1zy5epPIlWFnzYgkWU915HSp6ionBugGlBMMgiM1PC3zdmSrcqo6D9g5r
T5T93SHResEb/Lhl1q5DEjAvidDq6KZcli8S0xyxZCcs71pIPCXX9K0qSXaxTkfsjaFT81vFgd0U
IRX0zNu5vlSXNgsqiZ+CcjhCT7K1Kruj8iF64eRJ22rnB5MXpsmpbakEUw3KxnlHD5zPdOdNEWFF
ldraXi9VhPN/8584pzaKrpcFWYxx2cg5dV5v1gEFiBv/5MqL3GYEqJRdWn6W669NOyFwtGHL2xau
Z1SRScVHGppQpLcEB58tFaL8QCoy6P94bR/c5dpngFxpqM1nngn0cREhFdP7gr1gL2XBkUFGzPUp
sXJq2TDMw0qhxjgKxYD/CMWaZDbEQUnLKHyYWGxu8J+hWPVz2JTkxIncfqoV+2vlFUrg0OjNZ7xY
zYYpLv0Wn+4krKqPM3DSoCOt5CFMfQvemwXCCFEzKHYhwfo5YZtTUxTOGAFhyF+sgcXuSjvNvN9y
eqhr6zDivSWl8nEqb8oluRT9Mq6YFxbtIm+sHrV9KZsyMkztQOrM/DWtE1IvipAqeHzJV88djASq
xlD6Inkde8fXgdXUmmswx5cyh8fKbO/YhsWWIZqPlIT/ae0nBd0QBWbjpGad0xr4nvcRlGfFKihp
d5hbabMoCylZFuQnO7GazvzeX9fVUfpMgSf4rbDZBwxBKqnPY8S5EFLkf3rieeBKC+LctJxC9+2Z
mmL9KEKXkv174GmqyrrNfjMsyTiTmYqxT47fiJMyHL3iuawelb3pCjDTIGVuMTfiGXyAilQUmrIH
M8+d4S3pYLfmL/PEVQQdkDPI/gtuUetCd96QWBb1RQgV9e5bzZTy9YIh4ugw7AwebKKPLy8sfmvo
jAe7ic4LQ5ZylzLa4OYF8qDmUfBjCg9Xf93KFio/vuG2z0n32r14v4wZmnifHxP4ohGuPAChSVCL
MDBLWCnU3SAHo8p1J4EKZFGjw4dbSko5sib//tLFosgJsXwdNgfXm/XqjvlZ9/uCsEONHreqX1+v
7ibKfsTqWP9DQzIiuNvAAlk3rQmZO03J/cCs/cvGYdq5k4FgFcre915WWKc3JCuwuJK7Li3TFsTi
ok3FPc9f4rxZHQjOoUO4LtN9lXfMOftb1u73YOEaHuXz9/qVIkBzwjIO5Fg3vbVphL0BxH/X//wR
tbtgBSyQPd0GrLlFuFpFwhU+fC17jiN8VosD2VlFTPifEB/BmE9zF2KaBKEpfzk22Q73MGz4re4B
Xzd3ZTj3HicHMfRM8JyAi55W+aj2jkIj2YLAEGSGRj6F/J2IJOW+mrMNSBaASebhArCyG558GeUe
D8Lfr862NtQl87dbUu6FuZUY09TcTsYKezm6m9ohE2jn/xoeRPrB/15ui1LsBfSWTCE9p8+9YRi+
cvlNzjcq+u1yo9yRAj0D+q6BkgaexKXiJtxNmytxi+O+uMOt12ytzofQM/th3RF6S+2Jfucun4cA
it2uXXdi2EB9HadXzz+xix5MivSFbjzcFGq2T1frswhhFLOW7WTmbHdKJoDYlIzHs9vxILPurYR4
iES3H/Py2QJE/07ZErMxTpXnlSy2JQpMfA8d+3vR9rnOEqbQnxNT0JF6O8FN2cDViZR9Ize0NHzi
TNQhqa82NpVv9snZNM9Z+ka8a9sQYZmTSzJr9ApIdoxUkOhYOBesSZ2XL8OV47ACdqo+2FKC72Wd
Xp4vwMx1Tx8kiQIbdHkrMQ5WeKow8+qZo6CFX/Aly6zlw/aP7hwEOngZT2cLgyVc2Rj4bNzZfDdX
sY7upzKc1U3YAyXUaWLSdWGNuc1WeqmS6edxYeYdhkIi3w5XOqEl/HMUsPQ7RyRvMZebqhq2Fa1Y
Lhbkr0y2Jp5GpcrLC7CS+HKN+DDXMe8+YOJkw1qt2m8X01glgcg3Z4fKIi569d3vTDDk9Ts/ljAX
yQuw0XLcKOFMdXffMI7qw9gWMhH1H30hyRWvY4gZNQN2Cy4EfMqd82sghgkL7Yxx5FAszizanOXs
s4AlpXoPJ1Rq7KI5Uew55NzwrY++MAHu5+ajoBEcsFHXX7O8eCvhjKIKs2totfM4tzYcUob8+O8K
MrpFKKEvNlAepN4Sb2IG0c27MHManv6V9mImB6iJ0c9gfb7+08E0CTyUTrpu67mA1DLrqF+DQBob
JAN3zoN282XDXZcx/DFghJyBgopMUyU5T2rS6IxWtGOuPSd77xVlmkv5iX07PExeCUOYZr9gh+wi
fzu4VF9nJQ8pLg/MwVXUdmtVx1RXA43ezj4zHXCsyj8i1qa2LoL13EgdFVKtzUJx7fBL7+ZLnVTO
99x1736Q0yWu52+D9eAtRoVNTJssb2Yy/Yjxp2T1aGAiW6NCOtGef84O3Sq6jmyPRTlPr6HAv/Sp
cUnAaTBet0mg7PnCtYtenuGLizAYRj6AASK+cE9vVk9dfIt+CrOo5DSeqo1MLsO/Z2fYtr8im49m
EeA5+mRPXoRogku2wr96f6+9MKeCWy54ZRE/U8hvEXv6QN71dLDbfUuopvLX1IBBkk9PTw4tHPhD
CPgl0iclV60eM8gW9cl904CMkvjXZ+0aal7soHhKcNB2E17gPDOI3ofNjHA7nmGXukWYY47AbdPu
5JKO2YciIaF+dGBmuxAWcKqMrSKLD7p70gbRWPCzPtfzj/hxw/cLh+Dbp9CVhdOYjIFKAJq/pzr0
92uz5YAmTSIEhIdq6Nql3E13GnHKpLoOReGAoVYkMgLsBouUZmOpZgtLb4xSm712ValY34cRoAd4
CLjJGvwKoRKFpM+DjHJJwb4/rpUZLphxrITp2J4FWaeGIPMeKi6P8gJESTsZcafkbZMeCAzOch3/
6nr+BQAMHSILUU7XIZ1V84C1Vikr+kUIO4TC3Ng9XkrdlzVzwpogrQ4Y1nCaTmFWB2zKdVTGzBH8
8VgFh85JC5GLU7U23noedJjDTgYDz3oEY7K7xlRYDg1xU1R6dTJAhYbY2O5SEJrYVfX3KdytX6cw
rrbGX+8aF/db+5YtpY/2xl9Rb9XUv2edXvgE9kqb2mBF7Vi3P4DIwqyxE4Rv4Ivahad3Wh9ocK9P
1jz/BVgVC4CXXisSXj5gkgXLL8Z9eJIKQEBIcJsNui8XxwgK2VXoeo4O5PZwFFto8lmKgYYLrBRW
4X67xNep1PL7RJEDmM1eoaWABwzU+KLHAKKNMeXXAcIx7CPy4ZMT60oaCyW8arDfjmbtOzZjFUjd
9kWLdUpA/jpu2xaQzAVJskk7I6mcq92D87D7szgMDOPSgfY85w4ciMbUJ07DRqrVAb5nqI8qoM/W
kLCXtozI4ykqiAJetKJ6NupMhIXpsrIMBOM9qKDSlsuYtSAP8cAp6NbsAtGwZGKryqGy1f89H13a
5Aw2FRzPKrGTRscyjOMYrJxUp9VYLjmVk9d95GNaC3yAVAWu+or+yvYYBpNllxhsuXPQpiQmWC0h
VMccXwfrrXU+8ftCWIfQ8rWy/ZFnQhlOzK7rkXFHn+lFJ2R5QdY2gm+hUCm4uusv+qgdsLKOgkcJ
cTkiDfW410rj54PAM4Q6WlNrUuoNKh4FWXo1PBYyxY9oNAXtMyScHnFdXLtSGjGl2dgw8o/1fsWq
VtIgjb1YTkQEa0XyCQiWYZl4c3RtoBzUdGIbzvqktSkk6JRwjqlxg+kLi2AaAGfA964mbuOU4l1N
PmrFcBwO2myNCUir60EBgZhMQHyLAPIFmsRpbfZqXf0N+hnR8OBQgOUFZvLWfTpZBhBagzp5eqnv
tY6nvXNehJktp5zaHPXJZrTepMv8smoZv80oN1IGgw5nxWxSHzMyoxMFLjoUCl4CprO4eyc9CUGV
INpk5SZtYMC0TCCW+im3OH0PaxBNiKcmcUpkucU5dDQmaKH3kKJNmSNX/CqaIX0ENt+PMt92Y+LB
NXFwkpSrnUH+s+zJ/eCYf/kmFi4HfNgoVamKnkmzUHeeneWMTHEyadCTAKDwMFWKjzVhf8VJFHXZ
A1ApxJylE+TW7KBm+hAuBx2KQGgbIHrBBhwn2gzDsD8bZx/rPljNZCQAUIV1ZRqjYXojXZ8hsS+M
n1+456T334jORhHVePZjw8GlqPiIS0n6HYKN75rHy5xSMhgJkI81e4/GILLmsmAKSTpjhXCRoKvJ
q8BjLsNKViAwH4AwlCjFTsOaHqE0DJz9DPGP4zpfSHyJ1OWIviQyRJ+RbzpaHsL5uJ4Bf8cArMDH
A7K7FUv0ZUykv7dvmLzpZIIs41b1LCW51t2t+o7PMSi9uxO+0woHPYElM1iIYagAbPUQOmEKkQGx
+OSfpXTAU4Wk6NamZcfojMiP26Oamd2Hoodbev36qkmUf8tt3Szdbl+bk2GEILlqyobgHWRPJUy2
La5dikblp6yE0bOLfifNqd+0MdTXKrw2cT1sjTCE5SPz87so09j85/odLXBp3MenNRXZFqMbEARy
Spa88fSX3j8bvbmZGiqMOJRF/hZ7KJXVxZbMavPYI5SRzK006P+7KkymG5XlCcGXPmN6PX8ZMyfZ
oHRDXilEFdBhNwI4awPCSD0usI1Vy45KH9iL9vNPUGAVmWA31X/ElBXM6QzjAta70ePM+M4tm0YW
zfahuILQ+ayjGKaIWBQf0QgOczO4kOwJCkVC83wvAHPMYECopTwb+Rb+M0cbqby8+V322IN7QN7B
wmIUvP2EbIy84fel1DIfuRKjk9Io6cb8B0/U/yZ6VLNH9DFfd057o5lC8YGKbHk/oWuwWs4SMdVf
2bJdLMsInpnkcxBkbkKJwOguYFHRN6/5QZQaI2eD5nGWBUFqtWwc1eW9JCBjtyGs0vS9Hlks04q3
VaXiNhdiKgU4Pp4h/aTkhiyVfsrQiYxkLyZNFnerV2dXTWLvrPsVAQeIpBuBb3M/76u9kkIQwptM
9rmarR0isx0eKDoYaYxzJnrFQ4bFLez3UT3MyUN9zLoIOmfyrWYQs4QDt313dnbD3pkENpVlzYtT
yLyqpKpbFoeM27IqtY5IZMS2jD7vTiPVl9dJVHCFpUHeyim/C69SAVl07azDVN2wLbRvANGsLiLW
2aai0xnTMKzbjGRTyn/qZD168ZNbzTDRclPLySfCU/heZ746dJE/gB+y6Ixvm6ydKNY8X5XdOwPV
G4lmDfwrMSmGXW1HfJ29srKHrtYed70irtbnO2Ex6uJuriJy6tzx7VPOvTSl5SdCl3msTtvDnN+H
eqZkmvcp3IbF/lY13Z8C2upQwqFefQzq78RANUahTLyBCuOTbTAmukbeEWBzPqs/MbjgddA1HH3l
u2+pVGel3qtaqfPNxwMi6HH+cOBXzVomYbAgG2toospAtvw/JaKG55j/uVDA+0UUmSndCw97cCTm
1N25qFaBF7kwRewMWLbzCufPnB5l190SOHn0xwfOn9JJOjGX493kTPcbHPS0AyDECfrTKVDkyVhr
A2YcfEizuiSzv3kJ6TXc4/04FvfMEpNtMncXq9asdypnLRNCP0UWAj7zIBmaklDBinm83B96CQ7r
V+1YrLUYK37T2lgJZpt479qXgX+e8GsfrdArF7/s/xUky5wLRap491bMpoPg+eC3Kc9Cni0gAn+i
TzMZA1aNZMsrPy/VUaLg16WBHGR5iGsITmtHHKSZF6CclwY2dGtqqM7ynl9YrF/OaaaOd6+UgMoc
O47QdbqPiddVfnVnXCTpFnXlFVqLgHQi5NnOanE7na+LAKAT/rJ2x4WwxnzrVk1lmdeOemdCp7Ty
YmuCLtuySwzMAq0TuLJMv5pBbj/JEhMDlbAjy8LM5/Webb3HfixrG7ILgGSlZ83rV04jsEgDA4Md
AZNdiOhFyQ9uH0qenGNNSm/VfEe+wPA6K6Hq8rWpLdTMQe424+h3Skajbv1SbgGKDFThZMj7Zgu5
xxRje8ypnOd6PNpsiIm+8tYjPVkT9+4zkLLgmyU7hdLPBIMJ0StWIVlb3kUW2yXo3+b4uhX/zgyq
wDm2B9RWDWmDg4gHzS9h97QRdzOUp4TLe2WZt+/2gnBFtZntpGEOJdqpHt+gNyV5D58oggeM4T4e
9m6kPvUTvF0QbdJGzPXv+wtSgjOV52NtRQRKt54ykJxTjJbPB7EX2CzPf3vMd4XoGWXV/CCim/5y
+AXoUXPGQm+4z5tBam9ZpJwPhUV8P6T0SfPb7fIDdl2+hLxHeR7TRGQAwFyLoN9CERT83Zdar8pc
FtrObbHiQ3CXG25LXUnoDVhvo7Q3R/JIemrlLReTxBcYRSKKb1ah4sBUM94KaoVO3tp4JwFCHNU0
HPkmYm+EbNYngw9Mc2SqlPlHc0A8gvx9DhA6mhykHYQ+xSShbfxAxKXN4sJVb78DtgfmDtz9s2qc
ILoNEDjdYX8M1qQKzgwB74XpGXkVyTBTEu81yfgc+aIAF8H+pXfQR074ED65BtVpmuCmLPxfwomN
7f0i+TIEjfcXPG64ai3ExjgMo5VZ8k5uOCo2nRTpscm3mwmNbGiS9974F1lpshhErM6+8IlLq7V8
hmCrRJpDh0ysfQhAlfpf5WdsDuKywVWkc64L2NsZHKDwq3FeDnZnJdL1l/E/QZ2zZPI7nk8jOhgq
9oqtym/iJOR/4GVm1/JIIWAfTJsKboaNtRpwseerKyfejsL6dclXmHX4m0ohcw0tvbJui7QsgbHe
WAtl1RGujJBlGGC25QEpo6J9kBB0OTFyBc5PwjBBlKwG/IxnOIedE4x2rbGdnNhQNwJRq5hmxAnz
0T6I+oxzIwWr6O6jwevfat6fugSWph/AkUAssJ3476hoHYUWdMQL1mrTgpj0oQxEBBvb28XM/KWr
hsne/53SEa58FX5soxQR1qa/PNfHGZLvXcwB+/l5bVwlN2AKNc5Ntg6cEr2bk9EI2IXaW0tH3ilc
FErpVCZrDts4DIvieKBlMXEvukBVhH+7LtBqxFr/sDtDky3Z2qD4Ib/l3O4UBo+waptCDhU0pb5N
gt1IP7u/L4ba43aC06dk3UmrFYqKjuHx7zuPupSK/dveVygZ3u7sMUQLZjftMcQYJpm2Ww7XTCtK
y+0Ff8ZJtgSxpDzoVsbw8FcpZoOfkNOq/lu231zGtxWzBmNuBXb2dWdN/UQ5R3Vf3x/lpZOhoHnm
tnTmtX2HsewB7EPiue2p7+D0sQzfVP6ggoZckjN7vZpHS2BajMXK/hvNGFTuWdKoZDVTy6+Bn0GU
I9FAUDk3ulgiWYuErVL6lcBiPO0MIKqNotrnPXrKpGShPBgGYCXWUe3Z5R9ZmB+hjvxOhOWH7nCe
HC1GsyOGc08YKTQnFFbhGfnB9FLlRBIKX9ODyzKAgHfEjc7Nmfh+vuxelEtv66BVyQ+jTlCfymRP
qCywNcKiQ6L4ImJ49ASB3P2/VGGJW6HiR2YKtza4JWuOEtU/lnQt+lYQWDZlDIRdBlGDfmgN74za
PjUFXMbRmq9+ij71RM9VfcQS1PkoM2cjMXs9+Gqff73hsKkRFsxWX4dA6s/E15HCJdHbNDYZ92g8
ZnCMvuqtmUgaHUOSgXdOFBOVt9pdOC1DYQJjMuKv31z1vam4S2j3cGip4UaABkQqZNWCtBmUjo1h
oiCK1ijRDfIFgOe+GKY2dNYBIwAbQDgUq4p8RWDaejHXXdZpNnxVLyP2cZ4qcj0xSQUxZCARl2Oz
97iBD0XipJlJWHFQN5bVv3qKjofceqnmiBy6yd+VL6Sfx+j1TUM4hppydFFg8X05bys8OH2f/tZ2
dqPthmC0DmYcR2iMkyxjDoB9Ukz7Dm6tR+Urw7ivyofa+9WYbadnT7MUzBNhsKUEkBh937zyrGIH
HjMFEXQ2N28boGCw/XWaIc/3IJmmJRCDGPcBKfpoST/Q/0+SoJs5kHCRqo9jybLUtqahr3THR3ZP
NNYOCBhejWsNxBYsD3JJw+qkiyHwq7FYWFn6Tku98gDIBYEE61aMJBISIsAiNp6KY75e8AjyDXoO
P7l+LgWmkpTn2Hda4ArkLtY8ar0A2zB5veYy7S/enIEgnbJnEw7JYRCrtualLRZxGtq3S8rPwuec
+BhEPWybolq7Wuizt0X7Nl+lSdvKiAiX7ZopbGNXdKpJ6uYVM9yyPUgHEQt07rGJos6kZivZxp+y
WvshwiWrsO4HUT54MX+1mR+u6JmHLzHaIbaBs+mazui7qIxuIFmLljI3TAg/0PMY9HcrGpmxiHJV
x8mV7uULt7x7pR/fE/YBL3W1i9RDkrCemmuH0gj9ahT8k0EXZxf/Jj4snNoT0IqETEi57FturBaT
L3bUKYPwy8RRSxBrtieyyoTgPQwiSUeQjauLRf5uK7n5fV321Gpeob+Te1B/I/LevO3FFmvnPntv
OUb9z+o8vj7eByvp0xdP4L6AfHJu4GV0fDCeLivqpvyqhJvO5Ewqtg6HdA5y7SvJ+cMc2UQ7m/3z
zY7uuUYmDnfRN3JanzN4qyWCHluJ5xn6AUfwgyfOznhjwaGHlFyXKHXDkn0RTT0eHmVvh6kGNZ+X
ECCmrejsZE74F4ZpMqYCL60iTe01zihiMhXL69gEyREN8sOffGR+aP5CAOb/eruSNXWirte1HLAT
ijv+0cL1YJryAnqTDW6TUKs8QUhBAwo19njhQwpD1dLHU6kN0C9ahPcER74SsiqSzYtEJ6HJ07NK
d3OWCJ5tZovWnQdZ+Z6Cx/nnzqPP5KbL3lVG1hYS2xc0lsjloEIOP5PdHp7ruZNucTW8DeUqBFsA
0TNPJjj+63LvXGXUWtF3Ys+2FsEOvacRpP2BijgKf76E9AQADY1qXT22ry+wjtqsz7PvpPOxhaJK
qyaXpqklprm9vxh7MSeHZTSm67iPkYqlE9eNvgQLzOwHM2ftcrjQ2BRf0EOYCRE89P6CKDXOzPeK
eICJtHL+c5xw0bUBclEnzpkX5BOAYKsCAtBXRl1AmCpLPk58QwFBE2Op9BdrIaCPpU14JepM0Int
fSVCwMBwUSuEui4BF4TimbqMuzIFgwiYNSjUIvvH15TkzhcEtvAjo47irOMtBjVBX4xuGXYMsA1D
08IOxJ4WCf+hecaH2XTHsDh4O3AdtfW+6DGm+YjRNLX3bcYaN4oSxe7jXzJkXun1C+V6quyKhJij
yz6KU/j18bDegOyBGIV7tYWKCUswOMKZ1mockrIpXO4fsRK8PiieipRnD71W+ITaXAWajw+ldz5g
e4s2SRBxD1eHdnOiWQMWbmfroegy3jZzjdJoV6MvU6z9KdTYBwmBJJg8jlwMlNzSod6RLvSb4wqJ
NAI1GdRWu1YOzJGYTVvhhAPkVwLrueF5NLhnvsqJXZtDAH03EW8d3Xle1stgZuIhHRvLlUpeQSgz
jjyMTA/Ql8jOUSiH/VxPUxMaVUAVH1qeYeWlCxDpkI8LnxWOJWngZIYLUXrGsHu8PoN3NxuxJYWR
euX2IRaOQ9pRrLj+lvwpjCt9hC2WrTNiyckBrUOwWyggkAF4Ynp6Bkc2zG5x6x7DL2+XSDIWt7Ve
7bVscSPfTAn2vE64GSae8bGoYGZ9FfkbsxXTJcMCcaxLb5mMl+Blw6eARO1OHz+Oz1OmK4Ccn1lk
D3OT9nHThDW1qSkEA4LvhUqzzfY1SrFOT0D43YCuz5xCRp979oM/Hs6ppmelOuyHr15ZujMekV+i
OHP9nTWCcex3LHKoYyg+kmAdeU0Fxx6hcRBWxUsJtfh/QYiFWLiDAXjkhrr1bYZMBZNCygAQzM+P
zbdt2R5QoEln5QyUWSlhsKrFcLjP4XkX9taZAyiuDDREO7e1ALJDzDvv5GeKqa07p5ms/TbNmKNm
wTrlzvOc9wyJuU3nqoA8OuJqU4IV0MiRx3TZNXjCCwbyCGozmw9fYxEj0dZyX1fXLx2dZWaK+/do
fMK97qofYgUyUY70U6R/mh4yMunbQOb8BKd3LSE7i8wCHAGeYU6CY7WXQxdiftMRcS+n7agrrC2G
75BzDPXRvd2zYWQcV1q2GmhnxugaO0rVyzrspGLIcafM14946YobEtEHRDOPydQ7QB06oLmFvF/a
73ferTYT4aS+wA626uCdZid6c7sSm1w77rVbWf3wUgJ/64qy+ieZ0aFbTC5TOX3XXDdmxd5I/3R3
67WxsYnxyKNkBz4CJY1eH3zbMeWMY5v15uLCMXFDmQZR3HmQvgTqF22OvM/r422m1CLGCTQ86ywE
Dmm5lXHabtkMbhOxhQ2AP7rAfx5XrDtIY27kd12KewlfLAV0PkCCMPBcKJPpYLmjI32bYlGoTAiK
6Bzb/yKZyo+RtF4eMAQNUs3omB95oD6bb1MkaGwV1Ra10ffBW7TVDvKcSAR3gyOYUAS8V0ZNBWuD
lCbLH2NiOO36tnXGFjbQe2VGRYLPCMCmWJoSmKoWGHI4wy5uFtZHfe+XHKLf5NmjIS/HRDWNMEfa
UFXy0V+a1QDbVKIsYzFVXMYqMe/stUaa1HGFIKBBBj5SW65gW08VTTdzsJdeUJ/kYfjURw6Wx1qR
4Z4vlb/b23s7rJ6xHrFGS6SMUqfjs42bcFu2G23HOxoEve3y7nYYGq2mjt13yHGEwIE++tiw0L4e
Pih1+HJkLa56Tbq1+wy2M352loWgSv956WqS7G989AoigjT7fYrvXvtZ5PQ8iZVB9VLpwXyWbQSw
hQYHBylbH8IY3uvxUHTxCdmRzc1yq0uQw9dAN6XHHEycWz5f7ZzxW8dC/LD4QktLSmKI+euCmu6p
DaMhEwiGeHb6eA573A7Bc8TmVfcTEPILHu8ErfnNDtaj06bPla70we9XQE3JPJUAP5wS8q18RaPM
mBjxnnavPxzNssRS3Y4VCDsqeeWipM2gZZ4xPyc67USHAhCNmK910ZesKh8Xd2CF0vbqof3RaeA3
xnJExEdn21QvKJ59AZ1K8I7tMt9PCkeoAacIsJMtRBfKiXhbNFHZOWU0PvGJQHTAUBscnSO1SDJ+
jXSI46ab+joZExL2jVr4bCtegDVfKlt3mCjAuuqfgDQpI9xno6DFDn4YiidtWsrD7cae9nK9eOao
qCtu5UJheCt+liVGD7OjHJpQfizRFL+7Pj4AR0x7AoCgrSL6xFmlQt4fO8psHLSuYPfU4yvFLLQU
FaefSqS4dX+t6SDrhqVmYyW3gRla+JIDHLon7YWzmekaeufhOL63fBkNvek29eGgIyb/8dFc+LvG
wnfoptwx8LRT7ej3HM+mK2sV9SXZ7lkAuK+rtF56JLCsg+2v5Fq9ndAQNSduXiKSpcKlEWCv3hNp
3XzvtIxqX4XIb0d+7611XSGd0xUnL1bIQjQ2BpHSiqa/kl21HirTCerkwEGnhOsqOyELGqgfmoBF
56wFOiAJ7U9k5M4mdAsI8f+V4Zs+t18EMsutx0t1DMm+duC2dx+eBiYQPXyjJMoOTMUCBZuRjj5Y
vLfFPN1Z3FfzNJYEnOuJF5g5YZHrwr8kfNCcamEx5yHCz2lk+ap7Awr+Q0DhFImoD/Xzznt8YVYJ
/b5LhPfpYK/GbPNu7X/Wi8UQmH7vk1lFxLQ+vClYhJ62TxhBkPK726CmRuTUBykjS1/xmzYPvzH1
sgk5RKQV8Ax3lL2Uo9xn0iQjWKl3V03QI/HuT4gKblLJ4Yst0Txj/0u668F8PwRrdlr7lO+5+fmv
+EJPPDPb+8bAEspU+CC9IU6njeFvbZncdXzaQR6CLIrZjOXvoziyVMVJtFc72SvXUDR11plNPBqc
k9L+9mIxGZn+Dpqxy2mAiNmqx7KnWe7ZbwUckcGM0jwEZVgOk4BCpG6jo72l5sWk7+P0z6uZHwIj
FvaWY1KDgCupuIUS5G4kzfNi+Erk5139Aj45Qh1gVxHejLlUmp+eakgVIQhRLpb2wgFE0Lv4XeFm
9i+WQ652KGf+ZbsnHMvYFjpgBAdpTqMTZ6agyxWCPuu0RaDLlmKtS4HIZ3Mi/na5+EJKgQjKMMve
wTqFuUcHc/ipm4wmvgMuaivnriuJpijD4/ljSJxHS34UQkbzIIq7x6syf8Sw4uNAUm/bophoE8hW
X5V82nrmSXbcy9hlPZoXAdsgpa6Lqh1SSJkbh/pXFegSnud7m0qhpmNNOZY+kMi9zkryxohRe4TW
bRlc4WdYnZXJ8t7+inUAGlph4C86c8i3k2ooIYfG19+HbAwjECD1O6FwCiqAlcB+VSlfIULNeXUT
Cr1Z3L1FbjKnC76Ci4rI+CFBTpoGyb+G0GC77EmuPYyLy9JM3QQbafsnrbksBxsqsACPrNOWywih
l3/rDPL28TBQgBy4UmvkmY0OCJyrsIbkCrDOUJTKuxnuJw3k/aNHZRnGRlf5uiovwCOMdBQ9QfMh
USIW6FUU3p4RkMj+nrPC2rP2bbJRUwv8c7BfVOIUs8PhOv7Uvkdwz/23JL3hA7wi3bTV3Qatuaw7
icMCpsRWkP3XEgqER/GzX/Cpy8zdcwIiZw+pdnOvcvQrVe83LiLFa3hNQhokvQy3rpUIU6xU/rpW
rqOX/SYW9dx7vwXnu2+BdEdWO+cmeMThxwkNnOJLvV4BWtBSVo7auxRfKD0ZTnB6j2Ig6c7bJuqg
kfC11vvJzyzLQJz/RTKRTlpPDPEAjsx+udo48hRK/DpbIFXzhcvWnblA6ekECvqvy7vbc4BkftDB
vMnfTpxKMzUdLlz7iITmEhLEdwVz3OmdY0Vk6ZcvS/cqDSOS0U21cOK7LIc6+wx4ry2IsIrx361k
r/7p6hIe0TuqZHbWniJBFAdsCzE7higV2sk7chg9Tx9Eh5fgG8TJ84UWma0T2sQQR7kYhjbpf5x7
9rxwVFTDPlzuol5gO8NR1mp1BCgzQSo4GlRjSh8VlkhsPoxuvmriWwK4DO+edZYaQWNutx2HhLMX
3xpSWolsQEV/c9T2k+KgHCujKQ1claJg2IOiKjvDFltkzEVWAF/yvC5blZPtVCZi9sEl+YHjyFtR
WGNfZ39Xzf/uvKdQn2PzNPuCsMTqd3X3AOfDHWghqOXEyfB/DWKToDVJmSrANMeSuQOAL9k+jTAf
H1urLsq77Mer0SekNARE29QcApOSn6aCozR/uXi2yGw2gQsRWFP3L/6xDlH4tukYjb3WUknT+83x
OiBgegTE2TG9i1CxAg+8fdzICkEUyt+blRD8BtAKXcBz7HMZsWYP7qglmy4wjOHVWAeJhYJaU22v
0NLTFtJRwm4/jF8Ib3PmMmzp18ZaLhRg0VhMevwH0o1BIHJlleVPiwqB2GdCwkSu4dZAGTfm0EZY
F95F+6uyULjHdgnLIxvgBClXyZ0ThyjoHsEIud8CyaNSRxzr//lWnuCDjsunh1FNWZB23d8IxJPf
MT/T1wdu2qDftVrG3nDqjCq3oJari2IvyVfoKEzKxwK7xfR1jx09Fd251vmJDt+W0Lq1mEfe+M7a
ksXsJX0apPVfLrFQ1CXgj3L1JzmaKmANIPAwdQ7ie0dV281/TTi9vs8AMp+81wuYWCTkzqCaivss
8AXTVdrBK/uB0Z8K6Q3m42iyjlPC4p1/pETHHyxcO4a3yiYvz52U8kgzOj4LwjFBMM0h66Y52Rtg
JdW6C2s9qDvjTuGixkhb6xtdJ+TQ2uFe+odODHHXWVLAWnnZx6IpPw0ZhDFvUXtJHx6YUlt0G9Fo
LnmiZJR/gEU4JzJ/rwLPxgLWl0fhrLuHvOowk8cwmvGk6SKjc1IWUs4dzZG7tCjp6R/qMq3pBoIa
T2+hmTP4rRhzM0+B/fre2BLS1NNPnM2ndkxsKRoNOSq1kEwL2Nv2jT1irIhqlchXlsuumLxCkTQj
KxI3HDE5b1TSes3wNTeaIIrrB6DIZ0Xoc9EqkRp7H5qayiJtVrGRwpRMSXo5wQlSQuyZgGKxmv0W
j0GZzDFtoSZiufop2lK7jW0xARiS7rcjDFXAD2bL79LKjpyY091wby17HsRzr8UMAeZRj6d4VT5a
+vNqcaYs1pIeWlN4ZAIixVWmph0nFZ7mWmV5zDfsjpVHz5gsYag1JHN/Bf3PL08n6hZwlkW84OJw
cJzMdEFXhePocHkErdU3diNlwdeMAzPV+D4HjTUN65197CoI5r+6JviyO+AlWUHv8bTU0mDplQg2
yHN/kbTnf2fWD6rqAGhxHt8oDS4l4dQlXm8+CN3maqSG4fk5vxvICFFdZYyPSXOSTVYTK4HPGFz9
X+zzmu0YuqhODH9i8NUUvCcJdyQ1dZWbQfCfEnbItZMOx144eJh9EWIF9tPKfn4T28w7U+sFV3K9
/c1druQl9E/y5Z4Wu2iD7nb96V+EAUrXoibTgsIgtL/ihVJo70qT9Dw4Kjsl0kkTz+kXMUkxfhOR
TiYKJRhenR1YAiKOAP1wWm4AGawHVHGKxwMr2YUC2FvBdKvoRcg+FDmWyaf4HFV0fJ5LnJKpxfXl
vXNi+TNdP9VeyCKUUWHlhZhexRVwXYmY70vAXOgwdnOom+qMfZCX0myZudc7I8MjZTNTYEQggy++
0ROgmXjbJwYlklrqeDKgv5pjJJAPbbNEU8LICJIuQecCrKZK/1Penz/CBw/cVeCmPk9n0cMLOLKa
JZowkFhc9cmSOLQKawt+oZ0n0o2i1MUgQXB/kCWTKYA/ZARvAs5L+datKxwMukmkeQ8is9l3RJ/g
ZkqeAM7YTHjluzpc0bq/XrWTpUWr83rss54fBITFErF3QkIfgebh4lbQwacEnDRGDEx7Ivis17Lo
aFYEz32H1A6VtSAAYULlXJkXhQXqvfK/7SpIJL7iZ5arZBzychHQjDfNipWcF5I0GTizoQolRR6j
7FqVq2T3gtM3dKIV8KocI7WMuqm5gxzn10MeDvJZYmSfrBNzZlg+4MCNGeSbVPWn4zUdNJ8vxdzD
3UPpxGPCHXJfB81UW7wnd0IDq1ndD5EuKAGJuOiugAl3GS15/8wDaBMKtSEAIk6kXGYEzeWrf/7x
4kJV6uFrLCi3LdvzbP3NOQFxziTD67I/Fwx/ma1gZrH8dPbOUBQFfAJ7O4YBCKt1/NQcrHBaUp7v
usN1RXwNQgk0vr2nwCUTjoJ3Y0JibtiK8kWeYWgYoVTFsXrcrDshaErPghvlBFwEsLbOz+u4ywR2
tWC0AlESfb4j+GsIdxocRjrr2rgkt1bxxmrhemVFgQ2+JRsITsMYSZCPd3Q+5rE4NpNBO5ktFYA0
wCA0ldAx3NomJP2Oe+R05cKwVzZm6AbdVFEw8zNsXsdns05z+LSOT/5ZczxXVpzn8t4XXUPHeDt+
WJZ2r8/mWtOi2QpjD3F5Jabo/Jh0GhyCF3z7hGApsdf+TbzGwWo6OpiTVpWm/EOs3y3mj0uGij4g
0LF7zBjw6TiDb+S9TfVAIn2TU48rgA3IWYLarZklUqloKz3Hk+u8YOzpB28h5lAyfdRvjrhEeuVV
8jx6Z0QxLCO3UXVnmoO6q+op3FDI49xKP3dR6R5zt7ULqG5SEZs2mpZrM5aG1mVG0/q7dOwnBCy0
6pCLvGWOtooLEztZ3Qyg4IZ12fVfAD4WwHtqbtBBi2PCGleTSFq9GDe6pBS6X/IpQzozU7hGfk7w
Tt6AXem7RMDxyFyNM1/0m9FTNViArQtwjGDsRbcPLt95+Znpugoh7HoLTRCk2SCX4QT7gQsEH0PP
G/AjYjake05e5yoQZdThtCEUA8KiTVpkajgdOc0Eqgb4AhkmmPy+dqzDS4yeuFLD9aI1VL3Ycu8Y
Q/A011sGWzOXWfjYnrIuNSdRQf5u0B+wL9OV/e6yzazWnq1RJU7+nfTvMW9w/VZ99kr1V9GoNSp1
kxZH9SpsgpQyYYkTzqqcQZCaD4sfRMaV9p02kfg0a6oKAL1Q7s0MUYl4hImC5MICyOHwFWrGQY2f
XwzQi/PJokXHHEfe7U2tBDYfEWlAcQlv7rLe12msB6qZhGBJqs7CCcf1SwHz0oo0ZfyG9cttigK0
/aiMLR7pI2EWZKyH7hvTDwMfaqpImMRSCYI9MZd2YB4sfGE37fgNC/7/rGk/0Qjd8KZcnqkNmB6g
U9D1gnYb0sVLM5IM5DeJ+qup11UyM2C52uZndguzDQOwjBWbH95s/PPJsQoKATLH6Ss2oyA7P50J
EKJHIXa8nUAv9zYTJwYSsGVdm0gFuKMh3InIvtxMhg6Jm7up3zRF/Erwk2DwzcHrigWtskBsZpPN
gdweYVP9rB3rCq0uTUJk5fFsv2eTwkGNOGtYkyZyukNTQQJ2hkdXGpetZssZ3TvT4xf7zHjy67+o
2twLwXx7rULGtN+vuoRJGacc7o/IXoJB4NJ9E17nugRKOsVemKQHvsRlowQVTtCKprTL5VRLUQnX
HuBm3FqVI8iZjkq3I/o99W5V2Qzu60+c+KAwmv8cFclopDAQ0T9AHx5/z7xXC/8VjFSFfA+Ijjsz
iHmiENCkFuNekG7DAqwBa/VlHHtiwW6b5JWw0b3+tsKo87+MZVlUntUj3LZxQGauqGauDwscnk/P
tvKfZlyH2R9HkvRjTuPrAB6eiKhlDRFLc/TdtukPIIn9qeoAbsWDUmnje7Ja/Wy7X2BzRLKwSZx3
xJcONBXJA05x+0lJfitMLfinekONW+8k/i6xJBBon+QtAFH2AeqCcjMTF0pWcrmeWwkALpzcmjFi
c4cYJF3eYxitsUO97uNm60ZltrpIDixV5daW8g1FASDGzvCT0810lsnVZG/cdqem0gxppar07SBa
SX5RMFbp9IAQK6ilanTVafIXqbmxl61SABH7PjQ/TgqBrak6vp82/RHajObss7FBy6iL2Zi22lv4
GqgvjEIL1vQoWnGn5kuNCPfrTczpb2oCeFMCEcUiT07xm1twBkCcW0J+DtV5AQhlR/FbKnzORqTw
8vMTqoRFt70xM09hYofbEIi7m9D/TsM7kZyBtGRrtltBkMwF4FZmmx0MMpg/cF5sbR3ta1Hfpije
zGSAo0fQMzac5yKMyjAUv4G7tQYBtQ81w/BFOMQP8Xh61TYjDP7lheyGUL7QG0qOgcOhgtL+AdcG
4EZms9IwW450JtWLQVP9DXr8rRmbLU+g4dIK/tvFvARwW0YmxpYUIfZhZgz8LXH1Ag20Tmo6VhAr
5jc8c4ScTXaWNuHKBAJjZeo8rJNb9FUBBctIYcZxsC7dKYMrWhR+t3jGjaQCm0cVHkr7eP5rLs8n
Goi+PGfn+1tilR49+HcpLmMXOQf/9tI68SpSiUtcLLSeInKkdskZ0ZtE+TY6SCF2lJmCaJMpM8my
yu5ms3PAbTwHTFRmtZZJUkxQ7lUylyFCVDXgZQ5xSogesmxfsbFDzeVALSM9eycWj60PAL23aekY
CGMVfLNL5rWLx5UlEBH2GjQb3Vi5X3x8DDx7LvZwhAXvFW/X+lNyxa4Jz6PQSWD7JdWQqmgH5DFp
U0U1Aic27y+H25QqTCXjx753ERXwE++t4ocFxb9QZYAIrnUSa63I9txQcg9JDpVJgTEW2V2t5SnQ
SJlUr8ZyId4iIVpOwUFl4Ti9YDu/pkM1swjMkAp3JRYDm4Ql06NF+4S+pZ97uHnUbIBSbLY2nBtN
xe6JT1GGXflNip1qk1AObdAjYpeEU0Ysy+b7ssxOgBRaYji+/GVtnzfv/LioX0U64Izxff7xAg/j
Rygq0sA531z4Nu+Imh7uKEwt/NyseCsfgeRll3vQI5JIXY75YWbvVyaoFA3nRV7SfQR7fM5hi1R8
UWlt1po3Z/EsRNEb9jMBCqpMkn8ZDqmz8tlDMcZp1/tX8GoKyvkcZkEe75JYQytASzftquj8iSnA
3j0m73/2c+ISEkfixRJboSViaIFacUG7I2wlZYVtCvq6KC9coEV0+P0iO58rPhI4FNQ/9TV4w94W
BSkjkLJK1sunyCSVA7wf0oLgxp7qROxXuQV70g8CmfMQKs/iaEQT9yucDVNImRK7dM4v2EfuKD/+
PyQSfxMD++A14ioJ8nqiy0zNYKAIIWIjviIArtEk4GViZtTgH4Ggxo8B6yrHjuMP1170Zk/Qom7T
rkAGWY7nnTjJC6uQzv623r2Ye/DD1kdzOPkqUqgmI1+leY6+wtmxHRytd+/mFmxgBFXMYN4pGmaK
5xfI+47HnPYznEvF0iKT9H9N/VlKST9Mkwi9SWdV+y5OQAerkIJprE8/HwBBgSlSBgCtTiQmLRMt
Eb78HfZr2QAL+BBuK6ZeYOLXt+tiwjthkiA0R/wmPTtYiW1NrBnZDJisl2yNQB8sY4wpDFfk0ifd
QzYfylZuEUYY1/kpOzH9wuyy2E/WS2rUjbWhIaeW7dm+4ATl15HqG4E32QKsmrysqamaU2M5YFY4
KTARGMAF+aoAob4C3w8PQ/V4N9tfF+LqTlEMQXNynCjtK9mtFK8JY1atGRjj0ie9S9Ei89vwFOQr
m2pPER+KUoKJ3QdNR/xeCd/0X/R5lS9M7is0mTAmHEr6+o/Ui2lO+jdZJvkoFby0yD8YdtcnkwA6
Yw+q9Z48b13smMhQDm1/YedvVyVqsPA8A1A24hBfejYhwhfL10qu+0qATe0tRjzsV1k1yKY8yr2h
Q50QVxj3YkJZ3/jrT4a0S4etXu9rH30bT/+CStBVDq3Cxwl7OHGD0P/JaIkevLsoMW8hxGVP606I
P/yz/01fZ2fmxWob5BoKn9kXgIlYrEt0HAAkue1E8MUgWhWFf17gv/KWcydlaIOk7UCrA3zTaJbq
LM18faQQII9XW4a5AEPSf51hhg0UT1UQLfM6VcFjoEXCFLZ9rl6d/69o/tLkQOZ9Iupmlr3YUonq
Tm+iDnZ7vkU6zfAXDLdBV+R/goIIJ8XSf8qVx08Et4y+448pF1MHIBs5+gv/qZMtT4nZF9bdOIUU
ZtpIOQmg65fKDYgxOEaTZeMp//YT9vosIB9uz+OovsfJGJxxHEEccyBhxkV3fNnF/UD10cHrOSfy
E1EXUKbUOxuFgbT/6AAIjZ+gLVVGdt1TcE5MUro/b++paurToAhbU2gnknDaqi78yKaxg9Yn5yWP
0vgYIo122SDU44ZnMnmpwD7vPCm8fsMZSY3a949XCSVBXbGRBDmki1KOe2+v0ekg2NXiLhybgKSz
q4c4A9PfrByDnIdlr0iEQc4TNniPMPw6sOyBuKhbQilvQFnPAvOj2E92UJn9OpGyLPHTZxyfIK+J
LzVWJTw8Lf100xgxqUKEtmIVvU85B1p/hQ5TjvIGLupwk5jEi7VlMPa1nJ8hB2IzcErI8zWpDS9G
A6FH+9BQqqqUQ4qomofBWS3ubCN8ityZVUv3yc0WiB7dQrNr3nQ0cBT7twBNQTWriPkkRdaZ9pnx
W7c2HeFq3uEl2OFIEo/Q4atQOmyVoqer/EhRapmD6WfKbhBlzi0thE2CKvxOsq3Y23ft9dROL0Ke
giQRoOb68PQhjQp5QV8Jcae9HbuVv88R6v0NRE2JoiCa3BD54MIzZ+LOPXoLqIeX8ko8SscOP3yR
9eEtJg36kRNanOb/Re5blitu6bq2IIHB3ZFhW2pFjtUSuPQREmugk8j9Kt3b1HD0p2iAGUqEGzxa
5eb4jxqYNsdKqfnN0XlpFU60lmK4+nHzkC9r3qM9eXv5NazC7JqcE6fhr/U32O2ojFrtOggcTmr+
csZf6mzwdQHp+Y4pN/rWNlSodHhcnnqcYgQZq+6rUE+ajvpUSWY6rQ7EwGcDZW0Qe/a1M/R5edO9
lxHMmcgzN9GJGNBCQwjkaQfpTN96kppZ9G0pJ5PAoaHkVzW0JYb/5Y5zCyXJjZdY+sVHLya3LB34
McZqHvUH+IbkQejoQtFmCc1rL1YL6opvCsxkR6dhxMGGO4K7s2LULcxH07EP2ZyvNsAbCB/Gcxkx
U8vhVGIjwcIHcGjBpK8m5+naSNZxMBkZxwju98VaLTGez8hn3wuLzOUhj2bl3GrNKI0+t0AMybRa
QHR/AIc7WpQr/fACzolDJdXwkS51Pn/1n0ANnevuHrEEdH46qj8Q8mnm121CPB0/jNtNrgdaybnG
sYDzr1wmQ6W4szlb4n1ENRGkS+ex1heYh733jLPhe4Nt4C8Th9MfVzO9x59RnSKsDzC3c1sV6g41
MB3pT73sj06rpwlskMqpfAz3mtYg2PiGbfvB9VO5ghOnOcQ5Elc5zKtw77ZzviQQHlj9h2wI0vNw
nefxs15txFRx/ASGiTl3Lf/xk0ktwXro2A/yyM6OIgxXLy6I5v/MurkpRJQ+LUPkddzsSF/eJsR+
hr1YtTQxCoPHZO00FeKntTPnpy7nh6YZylNWo4Hs22b3o4D+7bpwdMUztvGUUSI+JCPuv2FSbQvm
u18sbXLCohhLtEivyT7o+smTyblFFKPJsVYKv+S7deOKd3mRvFBenEjsKs3Ou4+SE9ovbqVsv40V
7WYdMirsmflQPNZqq5Wt8IbSnlzzCWGvQzVyPAfOkS8gPI8Bf+70S20OpJ438OUXlOmfghkTglau
MY/Pvq5SlNGd/mvMt3EbPFTSXjgJoX+9BFv21sbghaMtzOtP7XqtH28aTwOcIVVZCourf5Gjjzy4
Ll3tMWh8L47yzj6cZpqf5HK1fA5QeT5yupRmiU9z3gzl/zzO9SGFMyELADZnG7OqMugOTQEvbH66
ute5gnSC4+OT3Ht5fFIk5Ru4DHHfjPgejG3ft2NbgNGZ6T942jESTHtoRTEBRcVVutObKBiYPWld
z3kXolueVcoAj0M06EkdZwMdtBrOqnzJY5w8NCI2T7f1TjHp1krY3YKgtWjqwDMs8b0g23qpBUNI
TYpAYHS0/jJSwIAaEpDObELdAGz183PTTtr1jVp9KO51gMv4exuNNyLtl5p9ZChtf2qx90rLwYlY
C9D21GgVadTqP3HVWRrnxB2OWYjpzwA10o6Ri+6uRx6FCDTT52dglCZc8PiCHE8wccqCRPC60Ipo
i8zP2oKwcseHMfXTO0tg9oPgto0WwqWHDx3a8aY/Ahlwc47uSa3XXAkGsIcUtpnD0ZHswTHPW+Ed
u0jWFZCn+VHlIvm3+whaHD33hSiz7vjuv2eC3QXdcoyakvuT3BvywKdrdYXJi4P443NjyVVfSop3
O2u7S84Jd5x+psRmIdBpuCpR2mQpPPkgIeDdYXx+gjzLCUyIdj9tcYpCRUuCvedJslA4yu34ped7
n8XafjRxzsZiUb2KLiCaBYGHPikboK4bpatf3Q7kLxxRLh6Y8ocJgZpKZNf8IlOwRV5wvydfuJBN
vWD+2YPIXQfVg9g76zyTgQ+PLbaVEKK3SFpsk63v3HYIJr/IuOLRT++KPHTuf36S7qYZQfjZWwf4
kS4FChHj8f1bMIIiegGcggYDjtEWAJRFNrpMM9QBt606ZPIm1tAwr3I0tQSNCFzlaIAuFarK6L/6
Zruj/Hq+To3OfcRysZjWUzkosumvWmT8KWuTClmGG5rO+6hg0rQka52rQsw4/QYzswvQk2oZ2Kq3
XSchk3dlxxbMTftHAzee8orMBMMJx6dn5mpTLe/d3bmQBUde1x1COM1dKXUGQzQal9EY+Ft1d/2Z
kOvyoFj0MxLbEeruApHbGGTgj6t0JpnR9w5iakLFxffX7QpPgBkbjm0v58zE2XXN2FFirwNByTlv
916eWx5Mow2DtMP14UHHFUScg1BjFNOtUgt/a1mnpleRZknVpzErChLG1ACY1wPnIHERX9+7Ry6Y
gDUYUcPaDxAruxrKwpg9tqelehKP7nZXt32++VyQThJ0aY/O3TbLqfb+/4bs2+7J3Q675joXgfl4
FLrH8nriLD0hfyC+5wxcaoQC1qhLL+zU8xe6VaCNviWJarspySLgwjPUoB0nwzPMKmwkSmciq+ZZ
XDse9MQxEGKAMq4HqkGmlPGlqq3nidMZc0H1ABJsI7tJD13hKTxy0jK0jz3gU6Pbz52Ypkj2b3/Q
QreMVE1qstHFdrAPhmqyVjBHLqLKpgvKYUKMKTICUW9QbvlHmsmFTzaH97+rvbIWfutN57JgixME
eLphxSO3Eqx/P6dgPXOJxT8C8T7CVxTBRN7Kb50IMBnyf4gPE+hTmOJPChobqX0vmb0M1+vJe36g
H2c9dRGHcso0QHV/7jYcphrkeeU3OCN9dLuyAz3Lk0imBHDViLDgryzmflZ7wj2eTc0NF9DVkoOt
oohshlF8kwQnVrxx90GOdDs/gLndqujXDh67hQkVYhOA1gRtlG6azRzbBbF1lvsgwiGZZkGkc4js
VNfiuCEOiQzFzTwFR/+nMEEEmC6r/8u/jVGl1rHu9pwtSIiobprjqEQwIlswQvuUnDBn1ZVtvXgZ
rTrA9wBAtoU9CU5Jk4CQvH0/v81ROzc+Y9bLmUEf4S9aTkyIsQEbs4gSp+hm1Vv0gx0l0i4lHjNu
nBt0AftpjMThq3nrIbNAG61b/U8BPRLxTLVbKWAZttyELeHuhwT5mRsgwFTO9dHVFhJ9yEzQALTQ
I+JXlDCdRu/w6D1yxdtNELMnyjahRaJIrgqAdmyKbVEYETBRJzpO4UYRE2xtUkdEAgeT7a4Jcu1X
veerbw4JKd44vspjR8AKoQUCymA4qjyzLKahFsbvnCxGLUypn8MiG10w9J47MDW6idk+ede4psW9
8N1DCrh5Escx6h5DTUSLcomMMUIzh9dLx0JdLzAxZrwL1IczW7yVlt6CHO0aeBCMy/vcWP9tGmUQ
aJ/234uSkHLpKclYwh0BhT8zRnWo9GkZyWIv1q4h+1gmSJGtn9NelrPYCNlNs4x/v9yLWsWq3wdJ
Vw+DmfFpsddrfAyj3asK533wALzKlbFIvCWqpsOU06ygo/392rcwX5kouh9e9dtSGKvw1JSn2IBo
KFC+VskLdwksws3hTLTCNsffsh7EvWQIMhT3zX+Eq+S6rkNQsCtkfKuJywPWc9TKM05tkjolP0NO
2RbQd2Kha1ITLJ9j04w5TR9ACEEiC1PkE+RdxpdL/JXuq6srcCoScZzsoT1+0I3EDpRv9gDg4J81
hjM8D6GIiWR7WNrAC4okfhkj1tdlFCcQ6t/BGzsrgF5xeRLkaiq2NZMaNy6OLT4A8icJd1VJztgr
YLpWDtvoYj1waywUe4BbH/sT6Z6O3Ev7PACWNyQVvTiycSaE0caKiWvsUPSjkewZ/JEQhyGuhbtO
RGg5XLCRAvp0tm8OSA0LUqgMloWaPSrYDmwuI94S6x3Aw4S9h1NTkzp6d9qjGOxpOgLDJiV3um5G
awAEZtEsRSkucH6P9UeEM7MqxaRsFGw0qUkIphCwVc/UQ7YCqNMh3vaViL03G5IswhvWT55tJSia
qjmsNCPHd6j0TgasL9R8zfC7QkZ97a4fYhxss9mR0TBkUQnaccoT8/3CO05FqHVsB5vYwj7pfVml
D4mtA9CAgUEVib+BgKwNHSt78sXFjYYKDkh7CI/oOVuSCMybb0gGm3KFUIvU8A/rO2Gdmzc7H0QJ
zVwAdd3i55ZSmVMnMxYWO9f/02fYNQXu7X29R3GcnDCKeo6/HHITOCOQkiOS+dd8vVY4gaeZZ/3Z
23e6tcqTZ3xUpi7RzKUgwl0VOcFNsmnyX56eeX4HjQbpBg5yozmu/bPmG03n4e1ILh4ErbAklOtD
mZqjNG5TnnNtRy/2AiwKxEOflabG6wZI87XtMoUZrkPU/fC+9pgtpB5Npfuc1ux5F2dnnkmSXWdS
/Mz4c/wAlC6d0kNfvxRBDkar2JqQ1SW3YFN74TgOg5mFytVjIICIalU9wnxGOcY2N/8EhyBDlZsd
qrGqCFuEFSyaj0Qb6mLfo8q3XwghlYud0N37ItlWmRxUNkTQZuCSk81hOybr/h8IPre3yvldu8kq
HKWvKR7DiQ87G5NY7ZePVwBrN6r6Ws4GJwUHcmgcCdEpM8l9UFYHZ2Cp7dAABXzLY/2sDI2WJKts
pJrv9ulWLgIyWnIYF3eGIPeBkMHCq9/5OS5w6hx8ySPXQLqlB2wTQcRQMYscOIat/geO0OYnNnyz
GME83i/CcpNhnl1wdR25rytmiOBAFWOiGb4bLirWmKoLjOV0iKCBTiLlWTw56YVh2Sp/AcX5rvL8
r+iovcU0VvHRxh/draFy9LbmI/EFW4KRdaqoMMWjlQwsxy28coDK+TexUGrZll22AMMe0k6dUvXV
xs+CEPm0B4/EhwUxgfF842I1brJ3JvfSUP7Qhb99AuX7mt3syKZmpCfb/XurE4lmx6otYe/6qvof
GGVlPiFWmeHUpEDeItWRrzMOhZctwVJTxRq7uGZmw12XYizPxWAmMoNRUw40ITF9QYiOkiXVnJsO
bx5hvxW3bXhzFNbofdHDwGYAygx/Mk68+3eqHPLCzTYtVWvtqxvglM1jSUsK/6+MF3fxiBGsPnzE
2cjDOR8Q26SmpCbs+h3vzZ8TChzOkC3uIpckxtRtovp/DFsKwNzTCde0P8QVBcwXPGHlS2eLaE3s
+x5iqMMa6KTm57Iw90DBVB8fxMEjV4y19tw7FWDz9Tn8rDxsKf5eDyi5oRn+tqInsHOQOXCC/8FN
wypT5Jk9fDlDR1FNrjYtvce+HWu71Nhh2qAGv0Un4bTmm8Ofluw9moGJUEup3A/XZTfdo1zO8FAc
2I+Btge7TpirOWbathh0fuEviU9kiiKDwlAFDMgbZfJpeQxVgF7YgFhvZbrpnHAdY5PMyQFIV9bC
hgSmNlgQQ6/b5heGBE1ZIqUQObaFDTRbDp2TgqR8wvL62wQYpkYD+xxku8A76puM61/2tDWzRaIC
2qP3y6tx7gHt3daiHyo0yICuDyXj9pkPtcP4RPlZNkih/5FibTw5IvThViXXEXQ5YBneljWdF3cW
+CGme4Ac4JAi1CezpxxBKETT0LjoZLT/x+7j871G1lcLsvOBVm5UhbgMu6/3XcYqWxpWMVOh1Ac8
K/87P/xOn/nLskL0t8XFitc7wj2b9Prjn2WgiYVDhg2pPjSeaUtNVWIE+9ABgaZqSlJ4RYVqWxgG
9+2KTC0bR2sYZ4dV/7uKrfVc6sCm3l9rzbmQgm7gygBDLY3dxxQaYmFumvoVSfQLMNBq0xA8Usa8
EtLRLTyv9zXQmb2VAmN5xBlIKdb/jvjmSGOnEYNNfqQvk2xYSO6g1D+md0FQL9KqwnDQhbmjolJQ
DjaVRGYwN7N1K/XoEHUyZYTiEU5KB/pX4lM0V4retPIoGebqLLnmG8YNKMU4ffkJEzXRJm5pm4EG
VstVPTHdL+PpzcnPWkbAdld7XSrFVfiiIKixifQWgl1dXwUuLk0oo4k00d/IVnA4C2HmTxuOCJe2
QRhq6TztOa9E+r0vxAzcBgpbrognsa9Y+KbivJ+E2uEEBM3z5g4/dd+xsfZVTWfAJkp9/4ePmj6L
9lKNzDj5crw0uqpnYQa48CaKXXsvnU3vhYxmpwb46B3kE4CLPZApvWzERwbr2x0DoRppKlMAtU31
9P0zWkS8kU/8BSHqkIUHMwMjFcFdb7Q+l6IvV0dP4d/GLXbHMNCW13cHeGdaSnaLmdzFH4xa4AvO
6Ja4qju+CaXvihFy0wSfjS337rf2j822XJ0uXL/hjZ1BSufeFDJ29dPvwlQLH500LvTomOP9y+6X
1H5eVON4R0RH/pZjY+ytqMrekLK401n2Doq2MhFU5aqUn0HtuKTVjnrHD7dyxv6WZBwYln9HWPyd
SPi37V05cp7IZ8l7JYPNIp5UFHfeL8SpacVO/T24qD9e036AX0iT/vNDNhY9A1PfnJ50xbdm3I73
NoOrasJ/MpyyGNDrD3G01ncmhFShh16ZF45m37tTrQLoFTlvtr6MqD8ESnYm7+6LQQxv3KlaegSL
nemSOarx7+JEAl+aCu1XA/GLx5mMo9ar8GU2rvrmUmn90eDZXs8/GbqL956X0br2oyBAabt/JB15
1jDqJ2iUyb3fs3WFI6BkWp5q48iMSEgxvNm+IRJpVGo99R8rfvKiKKqBxcRXqBe+cnTc4GtUrnPR
rpvzHxytQPh8IovHkRrUNFUN5n31iRGgh3B0GeWwtaoPdCkQa223wK9YXFM+y/onkBjVSkWEobq7
NVnhRp4rsKW1GWAcjT0acW2lNYf5UWWuQhL8MEuC2sICLRFR4p+kV7P4wbFFVo/HaARyuIlUKqHU
DlWRTv260xEkVabu40EROwJsRVGiaiKhOVdgZ+psQ3QD7RfQPLDLlNbg+8BW/aOWTdxuK5Q4dZP1
F3xz7oTxvIvn2NCRmTX2UuuiNR3zgG1wFEMxOeNUycncawZh4XUO4Gl7AmgXe/8vkTVAo59RVOt8
4E5QEOQeiAxKfeMNbmzYEj3OT1djWPXXoKfnG5l7ltuBMgFpL3zS3fxrytqy4w5xPQub92Q99QD0
2dyZ9gLKJ+vfIe9DZCAwgYOut73MWpfBDnJgFXuAqCv+XjXpSxVkoWU0kPIB0iHJbiOn901WjB7j
oOjtwnTazSYZ012Dukk+64035zhz0UR/8lTR0CuWDRVTGDJUIuf/NDzgwK9Qr5iWKqLJlGhNt4Ww
AQJY2yv+yoYCg/MSPsERZvPVq35imGUY/44z8+bQfGqRmMr77C2EWw0MHnMvhjzF60AcW2WiCWPL
uvOB1X2280dI0TVPMY1y2hRj0JQmEsYC19J+rIp7TfOHgGTeJ9EKO7DC4abhCPxbWyfe5+HZAoH2
d9D0Ha2dFz76skybgCNRDJpoOwzINigSfuJdnUcmTmmMCShQCVecqTqe+Cscmg328mLe7VC36Pwg
DW9ptVo8ck2a7NFhIVPjh4/OvAuipQbSa5JlAMuuuu9AAj/fuoINJ69jJEgoJcjeWNB1jz4YDfz+
VPrKTlHrui1cOI5WT6kLrgr9prPoMObDG9I2tARSN+9TpozaLNYzaAueybB6XExWWclHOy78cgX+
oTIQ3Gqddb9mPtOd4VLPbYurDJWjVOmIEpfOlImiNKPv2X0a1QNloY6ZSx6El2iEoLXd0gIihdGH
CqPilOhq6ykrQCjB44nuHewkA7kd6GEWBPKNWxbL1pu7hxWNygNtUpHlqaq+B62bH89RdM73xGt3
EkOGDLDy7tn1bQvU38rbdS0NXaqzBw3NbN16Akr2yjknOxC/NgSJYjIcuDbE1YKHzjg9v5TrBnH6
X1pB8LikGKmfkwuOp2UzEIpzzlOBjx8IVMsHu2zhArONkWNxmO8wP+Aj7MqOhvgQpgMsDsi8OJax
VDqxF+KWVcXkm5VXuJ7lXmZ3PCOMdy2IhIy2iIwdtFWsqj6z2eiK1NCvOoXjXd3xhtA1IzalKIlB
qca3mBJBd7E/GgptpUH+AAFbvwh/7C4uM5s8l4HbkXrJU5EbSVMIpQZ9OenFjiSapFACC25zwlMW
DXHeKYGwjXx+jPpxEr83yiaTwTxvxvddfDTle30GvjhU7HdA/3+47zK5qXpBaW96Tz/ZdAtFU1X3
mzPgSL6Q+teyVqgpttjRiMC0alyEbNSDOO/EhakWPtp4CR2rPIlm7i1NjSkmD4HwOOFDD5BYAwOh
SaxE2bIYqUPQEDxTepIvSxpMVbKdhtI+xw8XpAsNLz6QpDsxuYmLpWxdrdne+T9+E43xMRWSOjLN
+n4odUn3VO2u8ddgtbd6j2S3XKcc0J6X9RNu/ttgJATFNZu7UwHHAdxIQSoQaU8CErpMl6CGhgq6
MFKSe/JY+A7KMQhfVLnt42iUlfA/N0dVJw2ZJL2Xag+u3myD0RaJdJatUfRgEL0LWHf15g6is10g
B61dz8nKVIMZ/dU3YHZiOPaAGhB/H4KH3cmreuhxs2jJyH47dIjmopYQrTkTAtehEiitwW+5Ii+Z
fiJvd3X7ddaJscbBQCXKcIJAtGvpPxwJM8PEW5CvhEjk6f+hnM1W5BhZJMGd1Qn/SwCM2fIR9Y0t
6ZP6EBPifGFLM+v++rG1bPc0/FsFzO6uxnpn2UdejBhOWGK2F/alF00BiM+FatTzUYov7swyhM7k
qEal2VXBwj2pquDqHr0Ysh3MQXz2+a356AJipKaP03rbuT8ktqCa2PGpl+QWXTtZXg8AIMGDJP0N
wM28qzWT3PdzavUHLxdFvg05FuB1HDWxC5SgBCZfkh4fJ82wl34FRGQp60ToouquJfBOFp3zFMoY
T4huqu4B81fI/onh0gqZchBhNilbt9cqHZRhMvTgevK7E4G50DFzkdqtKTks5FxXjQGsrejFNDH4
u2k5MLfbqi8B8OhQlD/KaZB2WbS83VV79zBsuo3m8OqtGlNuwtc5mdv9UN/V96EdSZpix3HS0xvy
ESdIChK93221BTgw4B8CdJgd5lfeEReAsHqwt5t9IyG/Sitnw20+/75jnDvcvQGjycYCiZsUGqkB
4/BRL8INPJeWM23QeISQ3ao50qqoRtpaTS4XtuHgKdJXh5UK/hu8eLjL1Uhb6kPYfrl897fzVn71
+u2Exr65zF1pfxirhwYLvoMhshf2WE5FWiv/8zZdPpZ3k4q1yoGB/ULwkSuVwbt8PBlOHE2jeLGk
aEKVSxP6NhJqpeTdJrMjoHCA/eAubaflMXSCcadIUKwA073jtnx3UFTS8wtL/ckiv8BP24VXDy17
JjTbIuyUL0n5jCrfhyxa3m0Nnj0KgVm+Jgv5NAwT0Gg2/Vj0+eDLd94VIg8ywWCfC2VA2EVI+3kN
pg+ACniXP1W4/a4fhuJIFrjfskOSqGoClAMnFEVGIV0+QKPrASeLySQn8jRGUKH5RHRNp2d1HLh8
2RmMErKNXVmhwSdkHQWyyfZRNBslB3Rx8HjwR1NAWGeGOBABPYp3JjU/FRhS8dx38duIRIZ0hDGC
b2PHEHRkK3MmqELSoXqWVQFqA4x3gO3XmQ6IoQ5V/0l4DR8v4czOySoT6WGnx1BSwQI/nfELZ3sj
gjKzHfKMjUaemoBdfMbsx8tLEFkhT1TfD1qap2lwtC3PvcnGxd5w9+Kft9rGl/uZkj7m6scaKInS
WjEUlxQynbBQ7VAnpAA+OaPk8aFCrtzD3kIz49MORS85OlysUFX3PNVRlBprg6TwJ2s9L/8PXroH
q4NYwJyqKM1oi5osL7DVeAT/2IsmnMYeYyPa4ztl0WR4qrBXpr0R3KK5D4LIWL2ug4+SH0akCrpG
FTDKzukfEOMApeNZCKoDm9g82RRWGgxyjYU6V/HV/iwMW0viM8T4CzqSf6lPuzSlvafCL0uX01/9
pfDf9nqGZn6xjnIIkQ8PjH3M2mm+td6TjRsQ4Fh258i2UkZtkogi/RryDYIIw3H3gx+c+O37zmOb
FE27pLfYxqo+SGonQ1S689SGwdEr3BJ3vz/G78LcwRBmgYXsusR/Y0+9ow7vqzuFqanTDLvQak12
NMOIz4Fi5d/1uYI/umEVkXbfO+mYn+O6hEtSk5n3kzxYMf+FFSdOtYslJ0fsN6LUJQcT4lCwW5QI
EU55G84v478LSkXOs9XTGz7OrktbeYTOnZ66AopE/e4H22scCy4R+9C4+IXXfqS6GQLmFOc2RLhq
AyaOiQ+9U+gObGrHz01yfOTpcpFYPUT5v2yzBDXEMPzreidaVtBLO5OhYvWrYmrcbaoQvDiCbvu/
d8Xz+H7CGwnWW6DICC3Gyt5vlOyHv5bsZhAbCm/3YVj1ELoeCs23tyn44xljB05ih0QNWvlRPFM/
xMxL3F7CKYFYNIPD2khayKBe5F0WRgM17M3waXBrIbAET7PqG6VBIJF3NxnLBJJ6iD69PCTx2Mur
0wDQy0QTLuk2rNtjKWQ9c5N+wWEA90BhbCX3beV0f0yFeQ1SDiVhunh+z0mBN35LKBp2LBy8rxa/
3kx6UPpcJ1GE3oh8H2Ig3ERG14VXeSIpfR9dU79O6QUIKzVmbzqu3lyoUWuUgY6PdUb4Yo456PYh
WsVi+SSIreDV1lxwu5bwft477EJvZfiIUH3GrGODs7S3btr2tBIajZ20+tDjFW1lbyIhNe9oQ9wb
GW4gzqaVF2nfjFELOUjPdRLZ7rOlw3kIycgKaaH7kiUcfN9ls3TiKRPDIgIQA5dJK+6MQlGMagIb
tZWkxAI/hP6/2Ocb3NQvLzcOJimeO4Xtg+KCtBPjIlZrsos5SSYs4bZRXqiDvOu78pGAwKcSm9xg
BwW4XbIqNhS8BtmypLeW92Bsyi1HVkhHY351ekXAPpUf2YeQTgg0PLUseRwOr88xRWWZ0uRT3diO
/0QkZY77iIN24bcLmHqQtbe2RqWcWH/k949HjtjBG2vR2uaX0ICbNZhnsRyAq+IMqtlGTVCHsrsk
yyvniKeoDA0d0ckTk5zHxIGU2+PIeQIu0QqJWaHtIy0ZDZlZs4/b2gmkTjKI7qco6t51i79+wzZY
70PFLjNmbUWRox/ZPj3mAClW1VeeKbf4Ra1wvDX8m4EmDnC66Ow+C7b1qOclshWLFCupy46Gde6Q
1km4y8JfhGyw5WlOqjhibpxxtQNnTs0A2Z141IcrXWgJVze4aPtQt3vq4Dy/LcJ89bYTLRBrUQWz
lVbJFafn1vjvCc7V7Mo4hvIwVdiJUxKU4Y7JBf0Vpn5k7Noyh+ZOxEs/NNAJLfYuKKD8iCpCnPXQ
A3FZBBP5DNVvL3rbX0M/RSsBQYLFvNX7vAjUjXll3hyfYFKsRziU5W5IRKby4+G8XRzBWOM2VKoc
uxM/wLrcwpPeobH/ka5jCAuO6iyeXXCrfQj0Qft/E8+eYH2TlGp/X4l3i6Fkhq3qsntD7cISrYJr
NzdPpqzqVBfsMx2/xukzINhNZxPaRxyxoIYbK9tDbaLFhDsFyszncCMiQQJHcfNyLZr2N+V4siNq
NrPMvnD0As5FdWLrbLsboU02EBc0S1ardPvv3IDXXYmZr7e7BI52xqOWoSXst1V49q4rWWc0y38G
OKvlGmjjZtDVRd/7HlfavECPq0E/f41aRWhQN6IE44JG7QZ3U1ceYS79fR4dPzDOGgofZOzGumYa
vr9Op2rHub5KiL4gBIO5ckwJKFH3LnCRZp1yqOqcygijvc8ctV8/BP4qogufsbIPWdVbnUWZ5oU3
whCk4ZrB46qL9rN2caMJP3eXYB/v4MtbBCzIgzlLH+DQI2AxOOzgZefLsNKMO7N0cjUWUz2T0pxB
+1t93scG0GMJZZYEqp2aIJg92CFp+HHL7KvsJqO61tpwiTsFchxQ+t9bPdDvEhQzchAEdiGazUUK
74W/qPEPvIiCB8YTguZENAgjMDz9MR068IXfR7sdQrHawnXaoPjq8wVdqgJsftadSUSL97epi3Uh
GvLMt8gyDCMBKD+4MF8caiQDvit5brOZ8f0kDzR3LIBWKlG5+pBKh6SYKRwkSfaYPZXXwhjOa4cf
bURhuidibsRdUkaQ/o97MlxUOIzDGcZ8hVxQALxJO5YTXiVRvbfH7HhnISKYTniX2thycWOZ4+Cz
Kx92gm2YuotUxAGPk/7T9WeM0V9pIkmow5RYDPyzF7hT5ym/ydGXtwuJD1rpVXLlR07vgEfPLHpU
9+MTlhxfK5uruovMsZF2eFicTI5uANC/vBp75l1Aan3QBDBHTay43hAqg/5x6n3pfn4IipMsRh0J
43t48UuuW+uBMJ+c2M60d2TuzDvFsCIpcEB9Ts/8P8ockVcs/9/ij/6X4u3/bOAJr3E0ODj2DU1s
1IIJbbNd0Xb/2ByqYO8yKYDtoxorwxsOsqQdSyJrhKGr1BFLQUVH1p9nzIygH2z0nZlwQwHudvTI
flrvlT2EX56D2ITiMdn8hOW4Vf9fT3VYA0DWwkF761ih02XKct/SS32WH5IWbin5DxzQTAmYc2mF
gTqL/v2MXKKrlB6yiMga8ynaMnvaruXwPGJ6202U06IPMiyMGKNnFllgeK+WJuoRx0VW+44n/745
JCl1IzyanqA6AaaseLg6pXH+fUIWhFILAwlQbe5UGEsaXmrdHJZUhOHRoKSBmFzAC+bZXjJtA7Oh
tdBAEyBTnTLLExkDy53+jH3SpIbB5fgDHqAOLwJGGauANcDmlIyn6vwgR4Jx+JpWBDQXRdQI4N++
+rwnnLnXiB7gMLAx9CPb+V0sSiv5w1+xSD+j22ahGRmxo5wIEecQdDKqFjHDchBRGpVMkhGKa/V2
ZsczzLTaF2307iRr2B257w5/oTcjlVRHpsbdMODxgfuuztsO0tlwBC+8k1XiC97iLgY97Cf65R8J
mmWzhYA+S4dPvgcsYWho0PiuO8Los84Dr0AEeNyVw2zt4Lz/PWLYS+TKyuk5560byRYj4faC7Xuy
f5mqm/9M7aPmN3irfevhNbxW6wvTzDsfCa0fvO7Lo+g0M2n/OPgx69NYN14uZjT6XO/OL8YfdQsX
+32/cBAXPCJ4oISS8EaOSCtRWg/YHEYp8wV3yuH9Fs93dOrOy8TciwiYZK2TKu0yKKhZGhD+8bqs
t8Ip9qK8zH2KWPSgla/i9snTuP/ERsYDYiFO+S3DE2EdXPTseo1BDoQyrbqGJCrAjNvgh5SYuIVL
8zC8KQ/PY0AQQbxM/bYGPDEVwxy/KOqIsc7ZMqCfi6ZEWd0LP/vGOrcw8v6JUVQEExXd8GRWfOEz
Mnt5zEOyElg5G21zwXk5gh/sv6d4c+5yXCS8T+yUefjRljZ/0Nr8woT3KNbGM6EFYXWq0L9hxRc8
+rUQ4sML5UAIDicwREEyJ14OwxeWDzxnkih/iO/YcPo/V9JCXbzeEKaqmVJK7kYphKQkGl64uVUe
a8vTy4GTgXPulbtAF1vQjdfRb+EI/7jvcjvtKW9FLC5aQRTm/Q3oJJy3IzDd6+TGyEXNjL3XNRer
zRpE5E+EDl01uweTQHehSmeWEvmettG7D7PC5vFFyy3Pqe4rzv5NUYzpCwuWM2rV0SowZvlvvA1R
3amR0rK0yWbVuoBst1nEiuvIwaPGsSpQq1Oxvf20xdAqDpYrgJn7eiCQWe28Nr8txuqYf1Y4/Z2p
rT6PrFhyrlDh/96kbPidJWaSGv90O2Ou68GRKL7FPnjGXEkoYnt99oJEO5AnFTJB6tPbduGmnLrZ
SzuEmg9ILUz/p4TSSEdHz9hQBzwt8TVmyOqF2FN14OJx4EVL2dqyZ6JhVJXosj+j9WcjbKR7LAzV
RxowUy8dM1+5XlZ1pPfRUfZmBZcyKHqXuzsTKvXzuCWotZCmI4N5zzhyFNQpuMXPRm9pFJBwMP6O
EPRrPvaXtyqb/3uSg6BUj9XzzfnZpjetcSI7VKwCWcaXNqueHeOVYwbr3wJco6TXy6LWuRrFH+Zn
Se/h7+dx1CMiif5cv/WBQ+gIvI90hAnsbrRGcLpeNBDterTDxGReTG6Bq3c+UjXQ1u3nzKdKp4ro
EExMcZCU9nVNgZ3t6Zrs7aeEwxQyUzp2ovLqmhir8csweFI7q4IxQ846Nbc0EuAoEXUlyLTYEL1B
/8qN5DNCvN1cIJvHLFDeHMaqh+kmhvLkeqrmSikVtWubdE8CRHlGmmQGTa69JGniBJ5U0YEdjDMD
svtAou5mSw1VwStwGwdQNQ8f94nMKo/3bbkHFCOS4AE0NugJKRNMKDe7kWxFSbGIKLW+q2FKM2O+
tGhyltduyL3IiCOAgY64Q9Phb/iU8VT+0NHeSnaOJP5db2xtdkhL6/UqiHeW3+g19qeGgjNuUs1o
hjONSI8JDI1K5uPmbsIW4G3Nh3jcXtPq1abQbtUy45couHIz7ThmOL+Jk+M9Sxofw7TAb6yvI/dE
9KmHob2KS1zoA5uOuFWgJs7fEBvgONfw+msSzwanafCgGm5DpJzOVKxGVYYRNjfiC+ZK6RdHl/LU
mx0dCtP8e0TK52uVmFsNyFJuJ9g9JrXvEiT3sOIv5Wa3qkGyKYNOWxHkTJgXWmXjg884UIJJ9dyj
Kh3Fvv4UfmgTr3TC+gnxaGwVcC3NG8xxkqcgx2HyZ+l7Ct9TbtsCniDqCaT5pQ/5OOol7WASu/z8
9Nv4hyRNwAbxItDDAqmK5PAbFXjvxNAc52R6PJm71e1mAqfQBVpgIFwcvhGMV/SZ75mt7uB24bVA
oWsdP//jlZybpuL2tFX6poU1uQ/A340+msX3EC/8dg89bTGutT1BHqwgquOwgvMYEYZKf4scOiR/
2AoQ/OsDlJiKhibhYcMe0/KC4fz0+DyCVrXtA8oNkzmnm7bIyY62MDIkjfuKq++UfkWauyhjZZDE
7D+rWfzzaUt8GIIpozCyEnA2ujAibBbb3G1ApzRg3JkcNrT0C91voortCyCZkB2ezs/epIt31NKj
muxH9iuXVgXaSECnWk4KTKdSv9CMdWq6PLAJX5wBGq6ZjL7rXwCZNmHobGUlxd2MLcNCFWwrXWMu
KhBkxxNT4saTSZWl9Y8bdjLNNRolmp5NDIgZXVuZ8ORC7aWr8aZyDUa93P+OA4sPvbKSVX2FG1Db
GUnYZGht9jBXmRpbdiXkjio9E8akTY6G0f7vWT1mmudPfgn2jlCOtTA3wyTnQ+DOM0n4VSsXCw6R
dEFqYzGSSUuHyST8vyG38Wq3s/c7yqu2Ffj3oTW3TbI0zIrfBRXrexKM932DcjTg1wWJyeYSVqpq
AgZxLR8RSWE1dsUHgo6x6BXearRLoZiyAjoOdlrb+lvkYejWmyPv3bP8iiGTypXVRocKu98QVUDi
R/pcjq8PFRW0Hh5YQ/NlP7nU5xVaIKPKcHGECdqaD24Q89fXmDkaE+o4Hl2P4EyneT31bRbYoYp1
aFJ+lhqGbCZjc8G9NCLM54GH25Al8Btn3/5R7N9R7RJozlypbRFql5c6otpO/40lg+unpAlC6J+b
N1PKtEev99nhho7mCHQAg/gNQ0Zu0qT+hmh/Y8iMkdRzh+tvyzp+j+SVSv+8lRWZxyeliQF0Nw/f
u9S2xITTdJOFcqtv1vpQ1IYLz5wp9KUi0MkuvtXKvEDT2c0YjSob8QKHUaimHDw1QtbaOKDWGXsa
mWlaVTOg1hJI7FI1gH6gGv/NPFAa1+ztuTmXy6I5XTK5qFYpPkB9MeiQfMNj+j5pwiwBTATcpm7m
Mh9RrYCh5mgRp3Rr44KlvcJlXTmLVQB93NYag+BBHbpO5GHqMyhXTv3Pdhrq4qo7nlTv8XJNhjBX
g2AQAcmimyHLLmBB7LQLuDtdvVDVZlFhAhUF2ytHvdtvpBz0rH2h1tHXbx9RW12Y7FUaRXgw53L7
lrF51VYe2GayujW1t50RkOpJ9FuA8+buHaH2XDO5ReoO9PN/EzX5Bp7WDNtJUyaGfXiX9RMKs18b
C7PZXCxai08UNb209VRZjRW7RqhU8r8i6ZLsJBsDOu55Xi5KlgnbYbDA/84o7Pa4Gi8hZZThAvKC
QV9dhWqUI8rvcXIdTdiGI4sIJ9zE1TLs+Tk2RA5d+tZw5Tot1nwe/wtCKPDM853Jrf51PnNh0DK2
VT8/p+9vjdVcigZad6KjgkgqbyrcYCweuhdcxMOlxaVVRHbSKcsvBFzTY0JHqLMWjfqM4oMfx/pN
IN/M0pWh3GGaOXn1RunU53EaHT9uSy8poxnl2KjEQgOsMpyav6o4QhOb5wvgRIMTyQeQWDHfNdCC
qA2LnNOvh9o5+IvF1n6w0OeDQywQIK6plLxEJkMIeXfmECqGS4SvZKs5nzK7RkObAZGzlD+RmtHY
Z87chQ0+KjZtFSFNFM2/tHexI4pTcNj/MiZTR41QB6mFqEZjegcvibDvJRupQNHUN3cRUq5iN6l/
tIoCRkGpi0qra4EFdqqvvBK8H/ixZW6GZ3PrkmudK4kf9k/EGRmwDkp7IdKgnCzXyPY/h6tBc9Lc
d+GckobSRt14UwpNp0vr9kb3BbhVbknXlmKp4/OYdsdl7Ol+AW1k9ayteWJS8qEVpROBCaCtu2jv
EY0dhH4UhLazzlNUAwpMHkoRd5MOBhGGw2C3s0Eq9qau2VT6IVb2js+pwlH5YKB9sPKJZxiJ9yx0
jhvjHkrdb8LrqyPZakEUmYCFjjdAcQ6/LIz+hUr2SHNusFa3NkYRX3Uq+R/x8mU6PWLBm7BV559A
zRFc+NrV4reBf3OBKU9CN79/XQg35ieGNhSOtqlAyREFk1FVLhzpLRECY31n2AJqQhEQisnmYJGa
SOxt+nA+kkiv4AKemkwrOIbOXlK0tzOmE9Pv/xOW6j559WFti9UVDhJh+6kvblol6dDmY5Kdn/XH
fJ4umBpGDaWBiY5ijFoQNRUi1YuubqawP/dw5GRkjVEN/DCV8PT7K4F71Fx9VD+kD2Wx0Wkt8bRP
AsRQ1yKAOLyN7tmMengFomLmU8YL4999cbeRSQHVQCJxFdgcO9uNYbeRd2HzKHVwhxQJBIyjZLmy
ryUKt9XagP11XYeLywqhTG8fHEZqcAK7ImN+qZqaMWviIaos9wuwVAnB35W/ycPoeBAf34sB4cnR
34HhVci31YLOfUSifGC3AA8tZLiPY1WNh+JJ/gI3JYnhcqSshav1Uiii3mF1ubnevkzl0nFJWLoo
NH9isC4RSpeta2s3upkPp6x3NjYU/cFWalKZ5VS/HnYEqQDcv3DEPCNvJOGyADb45KJyN1F4j0+O
395WdCeVUnTVWKS7KvhGaUiqIrakfdGTj+Sx0C803VDIL2bUAaLcX+xgJQ7oGnKJyK+PNHd1u0BZ
FOyiJIUi9lZce8RfBXH7a12RMow22hvr1xT4MQ+K5qEkszgTUDBR2VngLvOoBLn4jTPIEDlI7IoB
AUGrDW3rnp3Duxpu/CGTWzcZ0p8671CpdNVpRFa4cLkgzUydfwuthHVae9TzNv6lXkqU1LPg0tbr
PbDXziVmn/eKp7N5bc2o2wnFl5ka3WuJacg6A0uKrxZLmWfBIYcLeMVoU7xlgsjbKNdguAXs/2Ac
7l29xGf4lsR3bCYMOchexGXyoHSv1Yj9rMzXfYTsoL7jbKNKk+EiPI7EUBSxiBSRS5IUvO71c4jg
PZAVJHKm6rbGr+4SnrVXSvhUo+lf60AfyoOdhL/sB5SqXE49xN4RAT8ayPedLqtKG752NMp3LCNj
5MBOwNcFkKm7j7cR1ubR/d5exZrUrpemBHuEYNpSruYAoftxRqybM3ppvi4n1Ppi0NkqOCuLxW+R
xxHI7ChHdr5VDQHFvxxVezdShd6UzdWfCl7t+zjaqjP+/dSFhKRh2NyLgL0n+WVefZRMPCJj+5eF
2Ta/4rKlQYWohnsYd3LRih2CfIx5R3bUHkRChNpsmVcMpic1dvo+z2fWuiBp013NU3yd6uvc0vcK
1d4bYBiaXEOZ3hXXEU2Krf9wWX9dyL5vZcpL8Pm/OQRA2l6ARaDMLDX1LJDZIsz0j/WoRVS8VXVc
l7dvWtQChqeFOGDMKq8mkkLw/kBT7jmo9M/LHyviMLbgQbCUoGyAjW3TAWUCkOpDNnnBc6xGO0do
WDmNzS6X8kUQkLFC++mtrTtTLwMEpA0DpxYVe25qRxRm8rTwZTJQN2G5F5XG0Pma0x/Jr5l+32YD
Vm7KC2diUd+nbmxDqw9CMYeWiheXo9eOp9FURoopZDNGb+m2dZqiK4npIoL/n7gHcbPEy8ebGErT
Jzkuht1ixYfr2M/oiKW9rzdhsvhPvt3Rjn7aEGkgDm45qMR6prQgGhFYxFfnaVc7Alyctx5yJqUr
AEbt/Bc0scRVOUTAv3HWZBx2szyFokuYeDWJ67x4zuWBzqwTDjLEJb0dOrlqb07KPL23zfxY92wo
gMLp4lPNSwExV5j3ckXMIhc2bF9Hc4lUCa54lCckdkHNedS2JbQ0ipx+9gM+AntoWT+URIV0WKc0
1RVa6iqqRywLNfXwgVCQB+gEPuUyZLaO4J9//i+TQRmgAnefrVhoxVYshtKarVq2FoHSfYvn3EVT
WyTEFXiN+SwiKcmozHfQY1f+RTbMcXA/ndwdsH0sliB31X4J4OsVeKFjpgRWcWPhU/wCF5Z+bhIY
bLMi9FJgpVVxyb2kAq/jc+gbB6bb90e8i9ECQoEWRl/0p/fAk5RYLuOJDHPCFY4buTmaFSWd7Gcz
exGG/A6tDmpVl8ipBaL0QwH3h05gtH7gqOF+LyNS5KSecN8/zCvU1BsgHijMmNsNSMnv1zy08BRe
5fRNd97UpgsNrNUxCkVD89xGfuiMJUNpLefJa7B2Q5AXMDohDd7XNPYDTui57VQ1yE72AW8H8C5e
kVipFITWpKO0RBFUa9PE5qHFvrSFlJOwu7YYNLmtzmvFFn/HCKNuxWDSmsYjSxgb78LeidLaKMrD
TQRHRJz4IGBDrR7uzKn8yO9Q0ZTXzVm2sdqLQfzjRdiPtlDoT6n0X/TD9GGa1JVywOTW42CJzaY/
OEH7CdOcYly6NCxKl6ZqS12NRnreW7PzM0/oKN3hVgCGcpIciaTmX5V6HNti9U3HbLCKSx4POiBT
ZCmHc7H7w9EMuejM2vPY9jUvE+7HmQKbmeNgpyIKpH9RzigksekTWRKCWnsz59wir6IRad/XTWCK
OqBjct6LDeukBjwyzMx3949rzlhdsVneSmC7b2D9/FCUYYx31d0qlG8Ms1mq/5MZpiTOx9KBY4eX
Trg3In+vsZMUt0FPN3MozGwtmSHnuMyo/Oazuib3pDDW9HNMYNOI8xs6cQjouGRBm5heMDDrOa5c
9UXN2HtxucB/oQRXd6otbZIPNebs0S7aEaveMxLjAtC05ybrcQ6NaQZ2sBLwrapYn7nBJWW3kJci
tGQ3PUO/7DdxTWBC3bAlXuEaWIJ2erj0d7tuPiQ2b7rkzrCXnexk+b5vYRrPOxu+7yJtCZ+Ai3ou
K/nOIfWznBe4gItrzQK0tISextcF0QBe17Y8VS3oI5zYcPB3kYywqSsRqdd/kvkGXYbIp0ZaZY9m
ClpsYMOJ5/ZigH5xUPircIqlAQVhQ6r/SoTwNRCve4QQ+hJGwa2aLQCCHywcXpOckpZX+e13qL0N
DFwGoNx4mZW6pvZUBCYCx074jMEp1J/CzoMYe5tz24Id3qqSee9VTl6jlfv6MqfRuhsaBlUy9rV2
p/vpzehFJf6cQQMCEoi28I0WbX4XRbMUeGAvJlNXS89JQpqRf4SZaWB3dscqx644IHM1gvDeKVwD
5RmdzD/SkHojJBzz96943OB/pcsCDPYnAmhEHy7BZ1CV5xwGQ57tJ4/Wf61C+aHKyBTKeL1XMTWn
aEz40PGHnMdtmw7o4Q5LP9Q7eH3ZymGjSdIhKtWwRYix6Ax0Ui7qLJL29G9+m5OvJQBxyLUODffH
a8uO0Mk7fvjtbQHgbA/+ojkUDyDAIY4YDPzyxAT5qAmF9C+pOrw3P6liSwWKT4ieXOLCZ2UI4NTe
MNyEWbEtrx79ShGgGCcO49KJ4JdCfacAWRjhUh53u2Z/CtCDUr7B/VAS+/j79hU6jn/5KEyxwJ3D
XLa5/dEx1gSxEGRr9JwZxkYlvgmASwVkCJkKcoEP3SSmU8yD66N2mYDpkCIIUYh36cE+guPsvs0v
Z+v+iA0S9cloV3YyHqaWQ+DtOtypevVQWv2L8W3BN3L0YDUUMOnSyTBW+8uxliJTqeaCjJ/8xM8i
6oEbZ2rZ0fNsYjZLVMk0ZaORIeecVqVbjXKkJ0EjBCDlZXjn/FF1/BHn29J5yWRNI0SiLoBr8P7C
4xTTWtpcZCUQY8cNB1d0aycxn8nlQHByH+jFaQb2AD8PphqSohyIzimrNcnjulJ6VFXk72lYVfqp
5H27wV6DNBJ4OAKLEwoL4eOtPg7LvdajuX1lW9sSslMH7FwXD5pV+sV6kLuc11dW1u/zRgH3TEDk
7RY+TtFTuJRSXC0jOdcYNoF/3IfSMxc3owFXG07jxQxaf0dOo2LvfSoHghrzKG2mbkEJOIZSGbLM
E/ahG/YpLwxm0lpf8caTKUlMyKFXajV7rwZ4fWR8WIke6NEX0AbW3EAC0PUM6v3LKmTas/vBJN1A
0ANY/tqqhXyVwSg3bAb6crPaIEFDaAksl5JlF/CuISBabkzbrkupmzvtg5ZGq2JNK0vpTrB6ZbIe
rr7gFe8Eycqb0wk5u6OHU033A9kjJAK6k6RxkDpXfpehmh4ph1IPf98Tbqp4hsFHCOxoA9JxpMSX
AYXFnT9q5dxtnvHNC6c4YSfs06wLNlaGL+rILwngssdQZ7Rfj0LdSGn1FrS8EzaUu98qHAL/7sXK
ewpSaXyShhUPQ2J6yByAMifQKSAqLtbCWVg2kAoeekqn1yI913H/SB/6BBRcNJK4r40UdL5a4anG
Y+Dg4dzKV1IRwOcNOmiUvhTlPJ1+4I3cIJQYn/OKfZR9dNYsTcD0QIMe5VcW5m52hT2Xnw2JFPit
U5GaQzuvNVXi1LRZ61S3KeZfU+ICSMUVR2GyQ4w3qGmgWbxtpWyRPC7dBh4Lqm8xR/dAQyGbPsOh
qwAEfv0EK6Weaj/ZE7nKjBujNcUGpCv1kwt1hOXfv4rJClKPzz6t97iK2t9eB+/pOCbVBtEoOwxr
NcJ109umyA2xjoR1JvVVkljNivDsHpzQT+lR3URGmbayhOKFMRiMzE4x4ZRUQ5K2aXj47DBmTbNw
WSRpmypY/9lc3t8Iq3Pp/7zXwi4UmeD1u7l20PEbuKghi6zaR35mcAHzuKE/scZNjnJmN1+rquYZ
A9g3qw0TqeR7PEjXDYAP+BrLcZNyzYTvcp5DULS5WbYqNctODdgsbvlrJyWQRmEnZ8kVWGdcdL//
IpeNOhxSxQL5sJiK/RwlHX0g/AdxsRAEoEr2mTX5UCv1l0O3Gd6rS8khNFveP8g4YXCbB80rvmKW
uJKGfpENPhgZd4rydmtDeezo51ov0a2vEkiBkfi9+fE1pOW8LaZcO1hVgpPtO89YAlC5tUqMLzdN
jqQtd+mD3IHcGG7aALOGacvEfT+osXQbKCcgJ+LFZYEWyO3tP6gTgNLHAty6E2BwURUYfLGZYuh7
CIRMuZoC94AL/PXaMM3X5jZeNiWoQZpvfKhZAdx2+GZ50wam0G0g1JFbNADGuM5SCeU45J1af8Bb
cqG0p211MuIoujvL6Tx/db31wvLHRGEOMOEc6zzwqVHuP0LoTMml0apZHsIpkIOUF/X6n4Z7oMv6
KUTWLxoVhlyGywPYSXt6oHIW55celH2WZ6cOM4JCVPtS5ocZZyE5t8wHEh7h8v63fSblm+ra/1np
xKIL6rznLEkRYcXHtQ1b3aplWV0NL+cXxAoGghkoz0wM75DpYOPXKhPIJ3N1nvyKD0qXd+3PiIq7
EDv+GrnlnNENhwz6YwHGa8eYuODz54wcTeSZbdtv+5R5ML1efvaRuErP4R6boEFLTsH+jkV7N/F/
K0BnCOpEQO5XN5stozHmpWOLFsHun03cP7Md4nuaEMQTHlO51o2/NBxBsSDJXCqiJUFHUYcSGpfe
p4b4eFokqSS6ekpSgMIYDMyxTA++tJOFPbZH2a7BOCMiP67aDUwnFU9nZuvkkw8WaQiOvaRu3uUL
u5BMt7RN+cd6hOxZOCAO7SEpZ3CzUU3E8pxNJQAGEyGOYFLm1aKibPXwxMiMlDJ+mXPQTKJ+YZSg
x71oIVelAQXWve9A1JADi+qpBdWqdzQ1Lf2/JMByE+qaisLWctSHoHyhtLU6YFaCMTKPJyhg9nl7
WHFBQm27VmfCXUleiLkDwIS0CYTtmLlCWAH3UWOtPoe/KQ6uCFpK7NuGvRljVyf5BakQTcnwM+BO
fTzzkleTS8RT5Qbm2B1dwz1+EB2TsJMzf0r2ZtwgH8aUbcvALQqJGUYhEk9Zl/6cNb+JivHLFQF1
viUQQ14qPJH0kmuVwT65o55UOzv/Kuu9NlwQpHHuvQWiKy8bdehGHqSLPCY5wvbwQrwnpkwAZgpS
190fyRBTkd8Kl5B09gQWxDRmmL/6N4qxD4a4QuOXNneosYUCWyfhqxAvqoQ3zgJSvYZ50owNP+j7
Liia/p6S6EVbeUZci0xum6568FNxz/1Fro4ZPIXKd6BWecJWZ03fQBF4+XbfBSPicSjYjOnw8wEE
qAgD8evgTq3vwlf4h+mqohKv8GcpDgDaxRciWitqiRMOTcVI6W4yYXwUUqKBv9KaOjdPuvSI3DPx
vBao4qLTJqRN4FBv3oHJ6AK83+B6Li//6aWvl5/JfeUo+l/HOnoyIVdHXSMd5uHJiKEEqiUXTA8I
3PxDqhJ1mGGjW+UHTfckQJ5pfXP9RqBoZvfNrApgN8T03PQ7nqxYTlUYHyMrPJMpbRbn8Am6zWqz
278hdQDJ8fHtOaAhWORqQlRQXbIctJAhWkL/9K0b896VQFTK6BJi6VmGW/HvoZObyQtNExvUUqlW
HjjLmDT4tahqqWEEKQKwuqPGBIhE9DfJvS5mOY2P3Ue7WcoA0PnmQ83OBpb39+rdY/V70RRl7H26
DnqHVTaOSYZ5s2sOcGUlO7YJ0bFSlGdxUz6zmkH4iqRhEalyn5WVyOz2tWHccQ7NvVp+DIgBpl92
g3hSVvzyN/Aw5JOIViL1IqueU3edMTgLYNKtDC3TPVKb2Xr0eNSv96ZSUIbhyxWSsXp368wkn31m
KPErBqICWjFkxDnMqLH9ow8Qye1NkLiPf5oc7Jf9oyal2mhxKSIi7m28FKIu9z9uJvOi4RyQ+cuJ
vH48jCbWmTQ4DLK+9pRSDsDnZduEmqcxlZZLpPSWQ5+eUfawR3yBZvNgO3zZ7cvG7DoDyQTROGsT
nQdIrsTQLPdpd2OFDttyRMJayuAxTB/q7BAme+dSehR54Ahe5GI3CEcR+ATPr5ypNmLCvLwJ/uqD
TCHYun66L0HPRqRtRQEctkqlfczxGLm1cBP8dIbNqD5yFjCWvUbuB8Oi03tWdyFzeyDQhA2/AsXi
lL0CEswNe+zjDTEdns5Bt3Dd3vsjjTrGKyQdl88C/XqEfJ2xLc8ogMcRJFK4pPqJY6uNRKdPuea/
wVZ8unVb3GwLeKQ1OAd1B5Oyt9F8fRaGJJ1wSYO3EO0OVMOyJjgqf+oCefIvY3uZ+QrpxXiKnQDl
nPCNcPNNTPNlv6InoE76conFmyN94xKUKdwkmKPcmuI00H0/nYDCIFVTAhFlA7WF5ZtWUH8/Z1fW
EE35DL0tR4oPgZhTBZin9YC1cHJR1Cey6KbwBjEvkgF3rjmuOXg8PLv788oectau9TC1ccXoQDxe
M6z71//K/OWNuDVpEUJbY9+5Poe3tnCVNVT9wMTc3H5tJCq0lFIQos/q7xYCMXSw73KjVvl1a91j
eY4yM3bEXLdjJSd1s3xUqLNEdydvOH+3v37LZDnk8HJXd2FcJY/rcU6uw2ABJx62+3CnX46M/nkz
7voM81zeRqIB5O4CLkSMtZMTgn/QmBa+GiglZ14qKODBkVuRHFQHZqlFI9reP/zJlobqHRh3HxGS
BFDUQoPmHZfSSCTX+NG6Sd870LWoioQWK8qsK+y/aJJCfVm2bC+3QhXbTopLv2WxTHEpuM8cLMU+
qsQXFLwp9ts2pM6Pzsfu4FZ6p1azVYSBNjUYwIt4oQ0pqAi9ikFW35RT70PFQcU8k0IdlCC1hzY/
NH6+KZlhL/RR/0CXD5x/SKnu+y1bSllsVKO77dB/2i7F6gk9L7v+qRRkDNMLng+ZP3CoK73pkpzI
L8VWE5W5KTYHjqGc6u+4fUdS5NgDRGOdzg3kuL/zXvjoZuBaxakdz8n79/5NDq2Ptblag/LfGVLH
lx4sGTzIn/FfxUdUKELDrbpYhuu5bJ68Zex6ZpXEn3IFXiSAfrpuXiYPHdCP+7Nog6OH2NUyEJqw
U50oGGy21CBOMw7QHxMvw13bFmP9jA6+r1/GvNl28jikwzINlP2Br8LnPAWrUKRhF4lxl5mwBlos
ablmGvOrDDGu+/1t6sVWtmSGMoq3xyni51bD6zjDAmmwp9DlBEKNIiwvu5GuRuMYSWvHFPiyon8N
qPT+3Nqvd0e0SW1BNsNB1QAhRmxmeH1bD6yP92PLEy4tLa2AwZvycWlnycWh1LzAw34Wu8LNjlic
/FN6la4fPvHha9nbyDwArafeqqmrYdcDl8RP7KTytOo3mq7s4ebypyZsTDFkTHtKtaWmfGU9julc
NZzT1Z3QfFtNuB+Uxt51N+RVqR3RS480SuExGM7kgRYuQGvXFR8mx6GJTy1sbqUwq8qzeC/CHZEM
G6eurnT79MwaFhfp0ypwA01p8Xn0oCs2lmCEJ9CbrdMO0MvLg7NTRZwsy/qJRQinemkguyroPPng
pzOMxnjHMPZDlngL1F4zzuhLMV6pmJJjIM9f+Zi2nMfdCllCB2nA+kizpyZOF23osTaqarxzp5kk
O1Q/92QishiCv6LPBbpUSiJVcE6AAkmlnkWSVTwUCJbiWCht52ijoM+6pak3ONb7zWbYkx01HcEQ
t0Lnwa0MFPKtYA5R3zDZgnP+YyhU5NMLj51sOdn3cEyLgaVeTtTMko/gKqm5B4HSiy73TTx9Zxqt
1imFEdYHUw/qszas4uTivqbCrk3O5DWZ+DGbkkEEE9mvvpIdAhNWI5FI8TS3fiu5g6vQy4yzDwlD
1a1VpbyJzjmnIfygACJKzWaibwxvBeZ8kOx0xLXAPQNtDlV7AC0bIylLY4p9XhnnkY8h9b96o6Mf
b/YSHcaGpe62OFyI7eaF9RGh1jzcfcKEkTp1+0kyfRTjhjHfsXHUjXBdY9/Cia7ZI4UNtC0+s+UL
kLtdPaq4+SO1JOf/i3tdVVMo2wYw/5QCEVGxwPJa00b3uOOgDkbGAOPEearrtx8+re+AwViQAuGi
zMYupuiBUAzGNGEO/e8yTQb7nHQYnAyRlK/NHvrBf/R5Kar0R5IiPB4xdNvXpG15EOb/JmVWyAj3
iSoGoVVvi6JyyUZbOtsQZPA0Vfdg6tspQh9rynjFU0aHY8PKWrFPaXf8vGJ4WUey6Dl7sEvJYmtA
0yTREcvePmzWBExOORiW/mClc9gwnd+SBqN5DcCcv2OB64rof04a1NEo0gAgUkpARWRJ0ysF6BAY
mkZGpxBAW0Hu2OG7kh/ChDU1k7x6CjFtS9MvtFJgVySPaEtiz1zquJcSZS7XrkGqR2uMpnJAktnv
H1jCT6houjerVTLCi8mEdXrOIBJXHp4cUItJX4vI5itovtJqkHkl2d4KQNjCSzMb1RlhSFxbP0+A
lz3Ia4MMFavcLKjYCg4Bb5lLOFqxWGg5GUXsm8AihZMumG5kFo4/Z/xSQpYtvaKm3PI5EY/hR7Gd
CM3BMCY6Lp65jEuwa800Bhl2Ln0VTNdgo1dfshrVpM7OniYuJlTMahMq6SbTwFRwRzXef7KvJTUC
JP2mpM5z0pTo7o1sxLEK4aMUb1et4MxCQkiw+BDzCEcrf2LRyx/HEBtb2XbdyvIBJMzYliu8WcS2
QsR1H9GssOSecP+8UTQ+E9xEF04+rCYCFbR4w0fiGOrvnPewN9ChaFqGXNwRpRdvzwATy856Iz17
DX3X7TytlrwIYUZwTicJ8aBbqr4mBODISb27P3nlCLGZoKUJnB5ZZKMxtkYhkunsN7ufEqWHdcB8
JJM1qPwccD+8vFStcyxaI+Qrc1i+VG+LKTOsZDT5n6XcjVICbpenTVEnPH1uP1uRNHqJiGcbTh/K
tuC28vX9HE5cKL99puT9bSditmiiNBJsN/WdSocyNVQ2/AWKdONy4iWd+T1Wk9y0BVdlcFSeH9pO
tadEkO/4cF0YxgRt/1UMMB/ZehK4RsJyACOJWXFbEdViUoxRNcdtvFzzEFNpvBdvaryZIOa6SItb
CPyYw7nrCUX0UCX7fM/IGvbbfhasckqlPtYqMtS5ap9zjnmJSuv+7UBv6EEFR/u6Tx0SaTW2YLqI
+fW3oQlSPSXrDg8eq1rJbF+MGnwO1VsNZ+Apgj2rERclM3+bhxoeKGR8hKyt4a/qCg12zPE8Ohzc
ma5MZ1sxCzCaXlytgnwXQtTlwf1coU8N4591Typa3E1TQPoSbCDerStT3dcB3B0gfqyaJOEnbSJ3
YAUiTWAwAdcl2MTJGscbvWqkIPo3D8sT7unc2DwU+Q+UftIrw2+bIFPPBl2aiKvSNX9HqYAl8L95
M2r+NGwdCjA6pP4ZnghIugrFde4jxEzdO3uT+wkSlVkhy11Jt9rm/Dq63bC6Ed39a5qukVitUvem
Sd0kjxypaAyIBAYrwEhu/g0h83GyDFsGvrl7XEsk5hRWeBMtnfp0Az0Lf5pz87H5TFKeL3Fv1f33
ea8/pgjBrgBrG8Al9YQawtQnu/hwyVGho/lEkgcWtdGgCYBXSs5C9YygERPzUABoGZpi590/cbrf
8IM4i4xdkn6tasId/o5nhRir/wm1uaq0r8Nvlal1Ce+1edtcZrCcPb7ZrTneFJCl1hXSREvCFiLW
HhI/MiYKWcG6WnrvPKdl4TRfaB3asLK+hupDy+gRE09+72dXKjJP9xB0AdJk5fpuLAO3hbc4uPJ4
VvL8wp1qxuwBQqDTOjWd3PUURC1ksHkbNvNXyddp34cv4LYyE0gPIAW8yrru0nM9PwNJfrkFEWkX
dIL6kdV2WBusV+vgjKXrzfRhU8oXyIHmk6iGIUF0DfC94qqgbDFRijIWmO4q/3lX0nlXDwaA9BOx
2GY8rVmifcNN9XYlRNRDtkniXz5mWlYTDliKPS58hsbSY6aU4334/AL3DdGPQ2b/gUMeY6XnMeGi
qOFSEfFQqJibU3UlsAm/+Uh+2cu5SFUy4N8/fBlL2m3StVg7jH6eGxRUt7y8ffIYhMwiJ8zEgG+r
phzEDQwX2th5UkRgHLEd5v0Ru61mGzzj4IiurC9qPCzMl+7Y3cqg+IrBhBnMMKjSWf5eYeWEjn9y
+vyI39ampBf85jOrLEvj+uIqrdltqYtrsYJWp8WupYNzXOoIE6nJCv2HNj7qCnz5f2jYyum3O8gM
wGUcX6tWasVYz0lprBMn52urLexv1Vl5p0zpZc3s5qmjlwralHYycKDHZPB3g8LfFbIvNyLB7YhN
D3p88mjawvLjsWPhmGLVekU/4ZaZZBST5Ce7JCV0oAC3wEQ2DXfgfh+f6i65GL/Ywu7SReZjuLdB
zSIQjnyHoo88NzHfHyNp5g+LD4z9THEy3txEiYwg2DgEpsxpzLtjNKcA2zkZk3V1XFCyKPlZiU2m
7u8q71jXizxja7x8Gjiful87xk0S1zoK5s67LJ4K+sPkEBm7m6AQcTg7ve1CKLiHAwkRc9ICNJRr
Oz/k6ntJ5NrbYVJDZhOfygtZHjTZHidI4QeJHYzsBF0EqW8ADSg794b7yMmJHwhA+6N0o+ipnBaI
eie2doYU1mCWCJ0uZba5/IZ30Sl7tEXKjp9d/IQlVPpPwCQyjOc5+DqKJw9S57tEErqbk0xdlsYH
l7eXKpF1Srt/rBVdOuKyydwSB+L4u8Of261Q6Ea7wu6v4HoWlWdNqNmoLUvP/HGGuBo5YuXOQsGv
oTUNhlyJBZzJpZrFIM5xNYSq+o4tkiDxC29uiynzUc4DkSBL6k5TNl7YLHX5mVkla2xuyza2Fc58
79ViXscCEdj8Og6UOLDOtzq9mgiL5MPJGEHIPvP14DN/vhfycc8fn6R0DS4IX4WymAXn5dSj7Yw2
i7juaYh7bTrqVtRCwI3InR8Okgt86vyiAaSNIKm0bX832cp03C8SnHRWv2nM0+s6ggN0I9xNcBap
aqXg7zmt//odwPB4orzyqNzdUINHGmeb7nNp5FLTxOHmorWMemtUm9iGKy9PN6wOiFGppYq5PdCk
pMhY6vmeQogB1Xan5htkYIpnf9VXk3JbZoHjkK3zop/Zx7g3SmcshVl5dFK9158eDVceYvoRdt/r
MHWH8Iq9trkYvhHk837uBJ4bUyetaNCVwF5JUH2YTdrlOMBnEtsyOSmpkFiQep9+bM2JrLONo00Q
sqtEFR0xev0Bzol23R+xvHJw0ITUhF0E7nfGzQduKBcQHw8/0ljjMsOJaIEPvX2PHV/Qv4BRdDKC
CTh1ZoHW/o0cIWT9GIiunFNPmKC39gxqi5K3brNXbgGcHlG7Ow5AoXcYKT4s0fq43UszsLX0dyM4
FickNUJRzIKd0Z9evBMzr7p5gPXRQjnPhhKHFXhh0t0Lcmop3zXVp06xXNMbLHjAd1o/pQEKvz8n
ahn5FjFUK5IUpF9Mm19R95EEwoTqI54KZzYmYK86vC0f8PnQ4Old2InGDkpTc8xqBzoqa5HB0CmG
qFUwpiFcOi9DDiAQB8G/AKbUzQKpvgmXAlKPrBY/pWf9C1CiHY3ldxkASFKAYuFp+yn1/RpfA7Sp
fLSqezB7mGe5nnVJt67zIxD+b+g3JuLutY61VqdjPPJ2qerx5vffGh40MDBTgefWlzLVTr0mRzlj
R3eYC8XMqU95Q9lB98sssc3zlLMgh4L7zaXLe0CB5y0qjAiQpNCBM2p+sTZvvVRl0g75P8foTKeP
AKyqr3aTJdM6t5yIOKvm9CFiDUTuVftBdn5z7CgHdE3qPUGbyuDOmixfJPGdU6sKMIm6UJL1lwQS
urMtFUq51NUqVO9s+jUHF/0Xz60srXc6q/eDifa8NrogGQCYWpEvxJpUVrnEKul1BBrUvME79bb5
XpLqyGtTD2RKNo8b1CzyF9gcSx7F+dVSTDRHBkV9D8CTZQzyX6cArbgp7+OzmsZvrCCD2xkfCr5F
QCNZ/WP2Rj3lnhR5YoJwXfQEOkXCMARGpCmfaLgmgCQh3o0o5D2WbfKiOOjX9FxzalD9D6tauSal
l8WZPr844ZwTsz/aGnMk21Tk/ezNOw0bSjW4H/VRt4X5HCRqbdriqgQ5ao5nCMp6Wn5iaEt7QiuM
CMw5a6xEdJE2h5UhVsU/DhCEoMiMwBCH1MfHrEqjT7mwnhpOp2mTXlc/pR6jykOh33bPdn0e2c1S
VWbtR60MKAnZUgqeGEYDJDacbV6D4cNiD3dWn8O82s54edcPRgX6YRHxXPjQ+1FSkDEhLVe+B7Fc
PVFt/r3AxjTDgO74vwlc1TWjbrMIA/1eC3g4JGLDVHdPioLGA4d2IE0Wp7KcXNQEuUtCaVpvEFPS
Ig37/Rkzk8udQOLvKpZdp6FuW8dDhFI4G6VPstWN/SuOHEuwfdLo1ls0qBtfjzLjzaEeaQU4aokz
f1N2yAFjRGODRjIUvLrQ8tlqYgY79rjYFOlEcKz1yCwF4/nDysgFL7/QgYiwtvP5ieBjAvfvIhtr
kCnduZk2bIvN6dupp2T/wgwOUiMDHcBiFYw5LlPX8DArAjS4b8ppop7xb3xG7rDCGon22+GOD+EI
ai12biRZu/FD//mfQM6FbowTfor6oRd8FAC7FuVIkHcOhdJKgs59gI1sGk8v/Uw8iCShtNj+T5Ki
DuUMvBXG5VEhGsKBTFa7j3v3+5GFWfmlzgqZ98IW5s39tA265z32Vch/7+FvDwo9qWSHSDnFwn3/
8ZKSlEIbvc8LDu1Pdep42dp+5+xP2q//CnqgrhJ3ANZYEbKHRVb9ZVQIzm7ktopUFfe+xkaKq3fW
1kD4CMSoZ9Ap9xoqtLw/gRLgBYx3uDl/pCuPoqqFZiovuenXkrJIYNmE3+gvjR87AYhwZhQiZ4YD
7UpH1KlIkpxRYAbuR4pnHVTez0Ppe/2jE+mkOd4NXpbVsCvUCea9o6BMRCZkh6aSat1fPpl6hy+N
g0iJ3Zvhp6avZ/i05X5/+7CQZwWzAVV+c1VH7v3l//ok6chR6w+H6dlhrHNZsiTwwNs1RzrqobBG
fsK4rcqJ+Rgv22a4Luo54Ul2XvwayJpvLkbbrkeBjrS7XT4FFluORd1J0EH2wg9rPyMNvRi8GZ5M
Mcq9/qT5J1Sq79Z3I1CPumFdJts2c1IsJWsicUCyshguVQNmdofwSDvyD89ssA96Q7yRpB3DRRj7
6c+KjCS3/kcP1S1AVAuCA+MHAqBxgYmZJxY//3hXI8xjDX8f0RfY/6Hl9Ur6tjcq8Jqxo5utRvV/
EeWI3qwXBC3oIZ6VtqgTDpbpzcy6rhQHcz8S48P+S3Qa8HrlllzuVm0ybx9LKjuBzlBqfxdWfE+K
f5pMNO5a2x3p2m0lQaqHBFU4uT6JV98tWNL1+3/GK+5QXVaceBFlN/TY/muXLiPH47M1Ym54ls0W
wBPYBZc04iBJVn2/2AjlFq+dXNcICV60jnc7SKt2OU6Wl04SuQki8mihM4BsS9Ic4SUwiIa4SU09
PRhYilCD5sTdie8FCppdvISrwrGrkpEeNyl7RpYWqwEgLxn7/o0G3WQ3/npEEgWVHA8/JJZCB5/l
zEnk8JrS+uukXJlx0gcYGTCAo2GS+6hicAknb0RjsR0gG07uhaCQy3CxtGnBOx6ZZxVcYxgveCPY
9zVCVHzQ7s2brt5KMt8lAoixQCRgrfJASSxISDKK2DEFeIS1SuTi6qncYKYvjdbK5uYJme7vfou0
gmR35EMz6qQb6aeE/r576X5YM0tXYxDglu5COhvhfx403j6ZcH9duxDITDzITvvj4gi/n2Sx6xrE
C3YmRjqy2uggxnzN46iNX9X+fqjkM3+ZErXyVaH15XKYGUxH+hUfEfVfVt6eqPCBICEpuvDfe4j4
D4CMmjGwHMLdYO2E7xnZ7ksBD6YUrN28x+EUnNjrZY2ndQj5cXbFvkfjOY3LaBeLDe2HkO/Yf2GB
aispI6kV4ubYKu600NAbLyoOfOKo5Um4zo+ETLJojuoZsKzC5HEhfPXGsQtpCCXYn7Fv43cb6PIc
aYZjR4jhD5lPb5pJ7vHDEc/NbYPMcwfTQoxZAm6Vz8BgnrSuYnXCBnrlbMNzOo3bKxqScoNBWTU2
QbxXr8bLaBW7y2DCMpcYfhgrOorNwxSEnRjbbXC28RfMsg8GUsbzjhKlf5U/1aRYr37voUa8JvB0
kvCvYkgeCl6lTjWCB6ADyVlYFmChUBP6aYhejMzzO1ONqlPXeNqc89poayyHf+mUDGXIghBCbxK+
2YFD/04v19C9lNvR7OLyDHTYoz3rgo4uYTskWyJJmqUdIOY+o3oZXbMLx5X5jntScin0Iyv2/WEW
i1MPE17AS7+HNXh/l6CyIBKEnF4+HhhiwE/Jb2GmgK+EzsfqhK+213VrJuNx67tiZpQ061Oib+8k
1GrLZ6hw+vGSmKp9R+3ZPzOTRtf6omr5jaLd5Qgxy0hPGzQ8Xy3rv/1+/vTk7Kyinvoax+qwXZ0G
H4W5JYmxbQyuhzQzZpz5LdFPoBJKLyTWuu0l0NO7r5SOoKXVeXRIBbERzfUJbpHiO8getT43UdHE
maL8chwpOLZbV5OZRKJp/9MldKmUXD6RiYGR+IdCCb+Jc7jarJT+1CLf6fFAxRLyDyiFm2+7OV6G
gcpS897A7+QmBBzWiErrlSajoBrnKylLjD7LW9BIccGty1BJu9CmV/d9XYRW2D6NV0eSEpnUh2mX
t0itcnI7FuU5ah7o2CDThZfnpd5xQo6uKraQp9BmXaJza+DN0t2YddWWCTrqVIwakiWTOMQJyRCe
BnV8AU7/e1jegO7Clm4dmisvtrkQOkUINy3f0QgIwF9/c2zGWnyvi3oWMg1cuwol9muPRgFZeEe9
EYABmfkcYniRFVdRPnyLFTjriHeT6GkTv0GYsTba97HvrFTIAGfhqr14xVrpGQIdpBcVmxYQjcsZ
v5nH+YiH1uGLwYrSmeBpHCS3nAv4QAq19O76HMBpv2E7EF1Yoz0vFnZ52diaO1QV4mpIXuIdAYh8
BmGycT31cPLed86FRP5VUqO0eBFUfMqoua4eoVSN8Vcn6rrDu61J2tHdVWrsQH3TZy/cJ+VO0eQ+
TMDoU/HV50SdBZixBBAfQdDg/V2+6FvxQGP6Gkepq5UNmce0Cfd++nZSaJ7Gs1D9CyeGLGjSTm8s
C+pYsZzKNuf3l1TWl3tIs1rumLgyRZdD5k4OTebB1WhLTOZ0QCZlN24KFC8SYqrFXQgaSIqglOMF
uhqddJEEND0Nl1nQeLDkEawLu4qA3shSxbEunhXjUJnTGhSizjEvwOjItIET6qh5aNKP45L/bLgv
6kVzTFWdT2jOX2AEtRGO0FRLx6C85dc4SkAeV7gXTkUp3EnoHWetrdvWYcd8nIHWuto4CeVa1Rat
aYlDnE9I289PPujpfBwDM3V+ofggvxeWT80HKxKS/rPFEtqzyp9OdlUA261qaj3IXcWGr+QLxPof
wo1zAN4YKsttria7dgOFospgFJ6ZRvozv+FdCo6TKi6thC9Ib2aMfuY4IaBiqM+kykhh2WY+53C1
kfgfhW3i1Ojk0u4NeWGRCJbVYj/JYRzuIk8vX21m6NBrg9KFYor4XgWJSTg0FV9D2y90hkK8uPTl
Tel9lN/eGK5hu2dA62WES370p7p+lmTmiAVTIKeYK1wDef/0nDpzmPpsVriMl1wpYoM5yLH7yTPS
XNBkEiAwv5e7nGQZYF+3mlXjouacMxsGO6G5juZrIwYCbQFAiIELYoJhPtC5T4GDWaVIGWhJlJLr
2ppXhLHeLYsqogdpsHg1FOXcErRQcE9gnLCLwW8htTuuV39aMvGaAwoD0EPd2aOpHMIOFJf6srIs
mAOsS4IVk7HkSGftOrHM2jRRUZykCGP5L9T9SwS79XdRu8n7S9uHIwD8e+MBL0gcdAWlFj9HitdH
AubcU4WmAShSau36cFmVpjZAChopykY7kMLF6B3/uJbzR+RxTHG3CafsrRBxdeH0RHLUMHY8MzZi
SI7jWdaJZMs6Hw6hS7mrz6sh6c7x91/Ljh433UzfHZ1VmAwxXeKZ+v4PPjJm28R7jL8GeTWurZ+K
yBZwkGRqFsL1FO9QVS64jTit82L2nBLE7lZu5jqitVAcWtgpmYRGNgPTSG4TFO2QhQXuSB9QJawI
Mp/0/NN5GQHqWbfx3xtHWMSLT7JJTL67DvxWmwoa3V01J0DSZvRAqyBzCJxUm98KkcNjAnRdu/iL
0pXD9H8CoHIync15V+YsA1NzNIsIu1itBrJEN2qy3izrztbYNZB9ePpDplaVhCiu/2f77Yc/USoM
n45+1QbX2mb8hVHTIkNN26YA8ssifj3tNn9FSICTi5ity+IiaMSmM0F5dKn8WNmSiVK1sBsV53KJ
tLzVkcT0cuUCfqEiY85gm8Vef9leGsp3W7xZe07fub+C2CN7yOdS0vC7hFlWtXwtcc+S8CVctepO
Egfz9eC4YecXPvr77U+UnAZWeFwux4QFkYyl+Ui1oayeeqk1MYKf1T2HbkBjSuJ7XJTZuz8CpWmI
uF+f+NREPt7Q7Cic0wZqR71XEA6U0xQBrfFQHhDJpCGo99XDNVDI7avVFzTLyetjgiWtYboQop7d
rkQzfH6qXWpjARoQPgwBEnj6RDqF7NPcFS5EOUY9EWpxA/l47SICzcsuh91B95bowW0BOa+vm+6o
RBh4geSJTQ1e3pavDCv3SFmyldFEfbp/4K8csz2CKDEvOG8DfGvueXGMPdWOBVV4QOLCk7qF11f3
djWqiH22WmVVlxLaph722Wm/cWLILvYKJnsn9UhrwsMeru5kQr8kxXUe42t0WKpOCnuxb+rH6aFp
cuifBnEzTE/G9GYxftlqRU3bilC/1+lCFceNOdc42TGYGIiKZy1cON2A35MH72jwSpOyzh8xEOvq
lnKoPIgcUY31n9cZwi+qt+g1HH5LCB+lEic8ngHxc7Yq1H0So07j1UmIrhA6ahNlR0z/xk9erVE9
ZnDVGoc2Bjorlb1kVjRd/XX3KX63/57eoSwBMWO0KWxcMQmHyxsNTaAZuQk7141KmGt91PyKp+Cy
jZP36BFozIBRkbk0ES1qEMhnk8f4HX+uxyeHOvOuzqjdcK7ocl16uYuwXmbGfAeEH1AHMlT+jN2w
uw5ZPHNYU5Dq4K3DOK+RrH+549hEb0thCZcuE8bw9+BSQMmsCJsqMN57dZnANizeWWrF2sEmN5Hr
cCE9YN+cgmOJzPdBpnBsY77FSXB5cKHJdF8bwAI2ikDKB06tjgkn8EjwR9gSYADJ9FjenFg1NgG8
u+uen06MmUx3U8sF5rmS/mhN77y5lxG65/3cBVX/tD5Cq850mlrVmfdaazvqyngKR10CL/2Fl+Qq
Q7WFWqvWZGhfbbU8TOP/U+HW/oCjQ3oKYMAOp3yFAdcoo/wAjXDvpnmNa57KhdzL7CkHMXvUscRp
kKDgw/M/hbAfk5UXBveW0aaAqJcDDi0H+fD2KXCL0z4UMx+nfcGncsN5oDHUhvSrW0ULqJXYH+Ec
dGR/g29+iVw3ft3CN/eRuVqifswQ5guUFc9jJbAvGmrZAKmlchbBZVopJAHdJ4hk3QbBngdtG/Yw
FTRAKBTh6E0lR8Gjgrx6YF8RodEYDkEXmVXhsbpz0oMAqDJLJVd1nqKBEUDTamjQ/rmmGRO5LpF0
OUkQx6pjNYL/BqkXxopcMPxKYbTNfY6QIo1tR0JgEaY5mfSx5cjn5CX7LEPC+N09JoRPFR8FpQC2
buAsAlAgSdO8mokfMSnGj4PXChi0qIUltNpIkWMPnKEZ/6DH8yyjenUmqjmi28bdEApIhP6fXUmB
W8MB4PhcHScFAsIKqSK/9NVRqoY5xY5nJZmEDq3ng1l4GQXIy3GbIzvjuckRUt8jy/qew7EdqNKc
hhZyYnJpr+lqFVFTb9HQr8rLoy2lQShjKf6c4Mbv4ixVyFOrBV5YJrm+GhbgmFkMYLgod0jtu51p
9VgNt0+DF0pB/F8hpALtvGCy66SfacFU+4iiivF7ARwStERhuGPsCBVUQXP6zgVuk4RhSAQ/udNU
lmOKEcv3ylJb1tPljKqelarDwzSvu51iQ6D/S0S5Va4CHT2vLvta6ITjXaO8dEADHv5IadwqtnwL
nF6qNVvIWYkbhlHeogTVeFm7rLeKIDE6A8nkususaB9KLgGBN6dmUj68waFC9qoypcYeBqVbT2tA
M2m7ywWofUxe1YCoI+HVx4oFCshcaI1TL2GcKQOEcnX05H3t16PTr0dUBrrDO52vY9ZUzUoi7KDb
55BG2NZUYfnpdxhhvi/i5Ff48rHJbZQ7q9zASRXlgUqfUv8YzobVhLrFRYfyRSN4gsbKI4NethKl
CtbHhitimsLseI9G6a7nuvgpK4D8pbEFhA55o9cav+H2wpZKz9Tmz4cCmSjq/rsiTzeHOvQVNXg8
7fSZSIQtPtz7i0tUcbT2lVOV7LbZwN8GSm5dTa40UPyqDJ7+oyky24+xwuSuVHXcsxU10bUAEeJF
ijBwM4NYRIkYoqIeg/kWIgXNmHZvFceki7y6p4zOzVjI3y5RrJebNAuT8P5DLYhFF2M1dSSO0Ivo
/1phibnacXU9bUd4bi1OKonNe9EexU67/jN/Zn/y0tPnVB39K4tBCHr9ZBTP0IG/v2HDVcR2hCNg
pYm0BWsDmYN1MBye6c6bU2jsw5/DHpOMJIEPrJMhpy+1TOjJvk6HomTcT4QEIuLSNdSKUwpe/yRj
Gi/f0FBNyyg5HQ4BYhcBAQ5oGddkVLvB6Q0loQ4w/IJ+7iHto9BJkW2SrZ9wBjpVzP8oCTICzMzt
JpAAooKYTLUd/atqgp2CgjjKDJSYgdzqpXTpuxwj2o/v0nZn/CU1Zrb3pcTv0XCGn6ETmaZqnCGP
vpgpYTtS4MYrsw8LqvAYl8uftr+lVYgObhcZXGaEm2gUAD5Y0yAZzwWbiTXP1shfBBG8wF3kWij0
KD8wmzA87gF6IbAq4l4OeyaI4qmbOBZY+Zoh3JcA3O/duO+QYlwVFXoH29GEo2cTbnx+3XpuM/Sr
knYwo+GOm1Zh8ITlyESB+rhBfvDOF008O33VsTsbFcmgozOQFipGRKxO1f1ELMAlS4oXzBnEO9ud
cEXdGqbQN2zMSkqnbtKOxB3FPyb5NaBD7c4yOJcVA8phmzEcWZB6UFqJzTp2skp1an22zhrik39/
irPF6XJbAmpBN4VZTar4Gf/eVmxHNdHpDKo+XD66Litcfx9Ez91yxSb7LIArTI3U6neuEe/k6UbM
abrF735eBwGN+deECHXOutyB14OAz+e6o9xZ89k+oI6HDooZl2x8O3gcbpjBr+voVWesg+ImZLrL
lNvMKFVSz3zJxn7p2fH3X85ynOPwjoTgPbHfHBzhN2LHTgAcrb63v4608FdGTzvP3F0dpzPFODsv
wI3E7VbSFckIHb7XCNupVFKdxynYnmf56YiwxXYfNNYGab+cPiMDMP0TuLvH3r3WOiEFA867ZB3Q
+68nOLaE6cbzPjD414IF0xATZuH/y+4lWRGyqxiJepo4jFSJOWuxR8pJaquGJcP2IbIl9gaAKDtL
hfTPxnXzliCv2ZDfKFCAfuTd2YwXN2lznWHgZR544UYULblXCWH59dZQwXs15ZQCHMFyrUU9vWGZ
vR4Fd4qEFTMx31W0T5/ES8sA33qezqmhtQtWSi8x7p57jYQzFn4LJPJwCUhs4vMU5xGFafPGIP/e
hTTswwLXjhTHM8TrgCUqv6BCso716lNaZs6PAON9mrYrvUk1NKXaC23hHyp8jDeeSE57r/AsUejm
R5gYTitLqoPLNqnsKBMW78b1LxzYtX4RR7CkzAIyKs1/5oy0ES7ELsulFv3+IET+3urMzMl/JsMC
ugLFg9IZ/PIgm42+eZIhyzkU1dU4qd7/YKRT7tbpZL27xhAyTJ3DLa4MHANCthaqTTHcN8ERNpYt
hwqflnwBEBP12hLH+rrJGrG/jqrxki/evzTo37vYbc7aM3AFTLPhSuitvaryYaatviGCHWLczlhF
Z7gunvt5wJQXQu+IQBcxY9uXZB0YYIKTFYplyJiJMLYZ/WAmlkpKxNMwrJYgBhcP2/UDjWvt043D
/O1zBuliRT/kesgkg2uyCAgG3YUVlxAYMtBd+316QgHkIHR3oKl+909x3QBvzAhEzW7tl+0hu3Of
lHAs459IYpX0VTfoIy6/KZR8A9CsTPj//5A8j9FiZbLonwnVh+PTlj2S6KamM6Vufi9wcT9SU2+q
T8QHl7RXgU17J4bhkQqAUIYuYkRxOi++z2F1B6ZoGzF64ILVD3RvGInun8TI+NP6V2sIHn2xSfWa
LrzEagjLkVbhigzMZWIsr4dEBx2hmEVhjGQhkwEDc6cQj0zIOpRbdlY7QRFFE3nQ4kB7WGJrRLbZ
s4yOG3+JC/Yy6GJ1ZfwarY9qoWrPNc9u+eMY0GhvTzKm1zF+tFoRO7ISljSFKxvm0+bm4w69LXme
G2td1DxK3iWkSPVzPGpeEyI3q7EumlzNtdGFZyROHfUPu1POF3D/PnYyZExklHBFLFaBkibebEO5
81hi8e36rBEdtQSqip9mAbJCegxSVn99Uv8AadzU1CJfrmPMazzBUKEqHBrkqtk2ocZngJE6tQ3O
/QiWt0z+jQP8dGQp9o7+pFFoWQSgL6GAODAcmFwQ3/CYxDkOMgX7AWTlYUzpKMAF8L70rtrIqblA
eRyG5xwOGe9/yArLgsyRPYMR+BSM2Kq1OxRi/AVaIA2ilWgxXSUWiD6CCURKCsp3Q6/I9WMleujk
YtzEwqush0wbKvWpf2iCEGmzzESs8aKWBAd8uJAvPzo5bcvtpL2mgm7TRmZh1XLAd8rzxE3IRyEz
o7P1EKNkn6V82nmneUk2oyi3b5fC7+0UBtzLAkocKp9Po223GVymC1OWf+SGUvkdxkBmeT3iluV4
3SXqnZJMcx6WzU+ErYOlLTvu9iN9x6sKPG+ZhQcaMjay8kuYBpr0f2+4MZ0zyiQbtSzrWE1QG8XU
GwnwaB6Gck5Lamo/yBzU4veqCnkY4HH9HxDDZruo4BmfuA1qdfFK07GAqLwjzCTqcZFHIEWB1IoB
OvhltpzbXvOBO70mbXU5Xvw0C8vn3ACe/bF817S3hKG76T33jrotD2Oz8bbYLia4I7JoNCJZmOtH
2YPoZe56FwnYeMz91yaYZkof51MCcouwEjXB9zxSalIx6C0lIAtoD2qYiNrLIE4Ow9/PPbIkp/6g
axSAVh3moqVEhvVxkGWG8JRxpkjmcMZ4eBO+utjQiUbny19422dOo1dIE1wBlXi33mYM7HsHMTwZ
C1OLaEHVRQM0+T5V5/hAvshGBeNPEvdG7kvS3IiMD3EVJ8BthZxDxXoUTbuHAWt5d4TpAUkW5xo5
I+5c1smysBDaZzt3Wg5GFZq1zgXprducfEqQUCAI4m+4eivwBrUhl/iHzVVhdXHJd26L8EmWj0ZY
nptBZYqCGFzNnhm0nrDTsVQEqJZLfqf3+ndMUaCo12lnOe9s2POFyQMlAYNiGmuLTsiW4Vzr2lwI
DcsR2TXB//VW9gMPv9Ck7L7eJ8udX1/f3YmvEYMP5n/mEM5esjVLPB/RuiUzmms3Xn4MwiRrhfLI
+rxfkkcYhDEtXZUgmzi7/Q9T7gEktYS1U1o64B+dhDdqOxG/O5qCE+0LukqCzOlMAwDMCEsQSgvw
OUMoUwaWy8LJLMvQK5PRDIBjuIVLon9ua+vNa6AUrt0kuFKiQ7ssBVvLo4e+J40FVTqq35pBvEkp
aJlGgR1WIbnz2AZ6I0O7D+ciQI0qG7VAVVZdy7XrZITXsg3P8ttn4GAe2wHEBb3QW2p62YdGcFog
wp01aq0lwjd862R8i1etXJR+feY4lSWohGOzKgN6EAdgvTH768PGnzOb9UDqd7+J1rmiLggKaiS4
WMokpfXDu2fYYHi8dRkqaanngPDluy42wCsehNLL2gAhbMooYCidL5uKXDKojms7luwnbsyX+Jgl
XZusq6jRgCSN7hsjMUAU5SdWecVl5dSR5vlwKnQKZ0PAnKxT6By6okVmv0JSn+BPg0Q/bz9YBlxU
t5xH7mL9mkj9OXweiYFaR2mr2I1ADceKekbYtCks4kXcgkKBuCoU6+ksIXUl9MKzcefs8SjW9eaO
4vOYRHm3O5DD7peZSOsdEEvbZwvouvi06/4o+HBcoBaxlUY4IglccDIWwGJTMY6f0SuO79vizNJX
oDaf/1WG21XxpPtHHkLTaeLjPyvhbTeYHloFDT3RSJEsrIv9jy/wKwrPCiojPIfE470r5IM/e5RR
kYVxKW9C/NdZaazrMp4WJgPrl95Yrir6dh14jGyG3SQQtv8sle5K8HVB+wZ3dHyKVexNYrEXLFuV
89UKq0GzdKr1ZwwtfmyFPioEnzuigEwtsMQ9HhTVDUcNJr6JjF0R9V4oST2sLjYZYIJntCHPwael
k1hQzlfvJQaUMjS1fx0+dNeHs7bx/i1/I1acCK8YXtTgB010TosatIQaWG5gOz0+0HeVBUZXcsOu
tWyasbt+nWMjzgmfrtSWPsDaZbYcl083IP+VRmXkh4vADeIcKT6pYhkBWk0F74GFQeBZU+aZcmHZ
v3833mr3F9ABDRvUFcG1H3YZUu86a4SHkHzVRiotIVo91JWXTHxe1roDlp2WzQtvuP55X3cMl+jB
E4U4bqPiSwrDL1Cxn3fUbyNjceBykfR1lZY7PNUA0FNuxdNqLpIV/OH9WPHqe3Axg/ViM2MX/KSG
XYZdavmPAJs+iAXIofo2NAZKCfdcFlmM1q2jSDhaGFAhC1AU1XvPQ2nTeBtebj7CucL7sb0K8HVj
aq+kQqctBN5Ed2R3iJQQ8u7EJI9sra+kd7ic4Pwpw7dB95h222W57nNkr/SzRM9w8j0bTDa0rB1o
kdVtUgEX51XHLPk1IdycTklm2HV4m1OqZ0+555wSziEgDWTZyGQ7ao2xgROlAoe57AQ739cm0Ib+
QczWGck6+6JYgGXxhAUxFJord4wJ7huV0FLCH/nu8EIMzb2cA+I3lf3mysXgxjkEQrqk1e5I0Xzc
ES4gjdbcCgkYLHSUX7oYZ1qFXU0ARiAQ7eaIfp94cwbakdIE6dzIbaihtjmGq1c9bCl5K2XHPLWO
6RdMTynAphx7Sw+s8XkNz09x5bxJ1FbCo/fa+wKyacy5cCszAcKrnYQgv7m4hq8ePxH1a+l/P5yl
MhBxDxeQyVMzWOT/zz50aIxjiZjYQH61YX7XPTyQsEsIHVw8gi7wIJF+L5njCEi4IMCn9WKpTu0m
hnmx6EDneg3SSgRP9gTomO7pr02IHCiPwevOlxqEyKr96g96LffOBXbWkufVaigpRC08k/739If1
Vv1V7urgafVqKtBWZy0IX5ocGP3nMIfRJxge4se+IlBwzjP0Y3M05BsFRYk07EsV5klg7NUQi11t
/I83705WmXZqbAe3wv5opuhAd/+Zize4PXZUEsSW0ozPDO1qJl5hf2uvIZtp55hOS/OcTcaf91Ga
ZkuTE8JcnU4NVRclfigq+qk0wbYkZryo5QG+ygDhArIlPbduwmB5Et3gaGQtR3Dx/k0FHe91UByQ
5/BCYccJUb0xvXEKR++eOvQLc2GAevNGBjqCERZkvuKvyf4XVbYKTKon65G96bkPlpgnsoVNgiTf
1bxIl18yeytlz+1jgIiWIjcZyUKnGYHWFusNSzmLNa5hO27XCdo8DlmHf0QUJPV8TUU9Vw7Wph/k
Nla3B9rTdi2QtUj9k+w0qp1L+KzWNLgOkiiTXEOczQ7MpFUOFKovVqpgJUrTJcfBXdJyUBXdWWOH
Q8aX7gLxzGpmO9bGq9DMwRua0Gn8zCfk39MfoNh6wzJ2Pf+xy7xgAvBaVGjlFdt9/FiKe59lPmDV
50ojLVPp+9IHVml3KnET6IG8hwz2WrgS8Nlws/HrLxrBdFaNL2KOTRiRTSpZJhLYlJtDSeBi4U27
Uqz2j3RdrbjYsdeYw8CcKvr8SMh3nPr0cvNwC6oTo53ANWUGq5y8341/32m8aHRL7PpOLHv1xux5
OH/Q3bdY13N12lxTg8dQXfsExFb9sufmOL+znOWAybBYLjsSFThBcSn4SDqLUVTG4WqhuSoj+xcl
pxGpOZWfscAPWx9/fp1AjPB9cHIjancd/inJKOEDCCp0lzjmFzFu1d2ROkjTF4amX5opZnVvhcU7
GZ3x/JJCYbxl8x9Gj4+c5bm/OahWzJxOLNsxVdnsVNIAkXdDfzGGI4S9LnOqPgyZRj4V5hjel+/V
avnn1T5l0UFvB+vmDNqGyT9TZln3ueukM6EsgTwKgDjfH5mEtv3+Kd0s5sZa+VYVRr1fxVK4BW3p
kuT6n7oyWHw86qwWp6W/cE9tFHeF+1BCH0t8zkZscpptKjx0M2MN3rqDiRb2zlSRz9btk/A99ueQ
D/PZXXoaLqvrnnZxVccpNruuj1olze/KV7CMTxM66WmEamEVzqkwto+RWaAwRRR2I/t3wcUhC4PA
GuLmyr1p6sQaM1S6Na0aGJs1wMDvrt1dLFAuJj4w+wXP+RxL2XjVbgTA6YUfiEHDa4/Hm6i+An8D
7MXq3l//l5AbMpLC35byJwaOtYQDVtIUkyURnSE0mh1WfFaSw77zwAZ9kOP7nBH/Y7iQVBsuOLvq
TtlY/i1H9pRPWz+Rw3PX8waZpq01i8Q6TIJ0s3aA055Zv+UKTVQkfqjgUvViX8PZH/F8XxCz3usS
49grjxw4NF5xy2PPSdmRBdDk7Iwg+gkKpK0//Bpk6LuASP6tLKLsPjVMdOQ/iE7EPgXteZNHeuR9
AiVAnjgi6TxZKSUOcT0FAxp/Oi5CAtDL98IvJWqXZ+HhOJKY+sNIqhH+l1mdQHEglPmLAT2yb/5x
4uBZC5cBRRBlW01mnMegM4ya6Wc5hTaWmjMXBEnI66eQ3MW1nDcptITmq2B6shGOC5alXKw7S5Hz
QsezmyW0SZNe7PU/eDmF/zRutm4Qfc5XjHOniDxE/0cPmEsHgnq/zt/fzp9P+WzCNtSjfbp9+Ckc
QBQ5EzRqLfOnXH5EN0CbG6+8MMPDjQw2r4Pne8WA+XxmGEU8l0EKU7Id3kjEfRF/My+YVFxEsKeN
+hqAl9mNxX+dLeVkZ8zxJFyacs8QN1mc/QbDVpScOXteDTJUtruzfsOkH+G1Xza+LGC+sBB2WF8s
BzEnn3C0GhdREluodTeyoLmN1sioPf7zuNb5iSbA96H98FafxXHbhiKlqxsUPWeig5dtQ0phNbkX
UNa1772LETFj44jmB9iDzqqt/0WgMYgL62VSh1Oufz2ATJVGT2f4xAifPnOK6hIxSLIo9WWS7Aym
isDLFWSI8CpwO5QWBmAac1Yo3G9svn11/RzuwYSrGoqzls0R1DJOwiOfxP6IhNsYl6h7PDzF0c0N
54DaMuPdVAp0O75SWNj02YnWKxxk4UOZ4xeYvcxS2v3a8uZb1Trqxj4D0jlVy1myWsQdq8UHMSWU
z/9BGb66lafzYgRf7qvBMWcNl5jTUk5SMJn51IHHPyxdwn0mLaKuJKGHv72u3PrJQ3AbwjxonJhe
pdu9hZhYbHpAA/kbpdY73yPoe4Ei5OXBriZEcTfnjf8lBCk/NxEZ6mxONgvfBIHMiNOrcYTF6rJc
5s3Rwmc9PFymB8m4hhq6SMnX6BMnDwbDgO6Q5OzGbuHnewQBInwAXFDl6qRkTXfLPgHsBFRDZcod
0oudqaIpSBBFMmNNUNPCsySh1q/M+ALKDeQKlgExHNI6eV38t839ExOnsFn1Tl1B3daQ5CiRCmTN
tM0ZHugVExSn/Eqf0IdMOvMz6ma6DOu0MMd0ZWBKok5qdkQPmXTXFlo6EbiprK58LOOTQh7ZOffG
B9ChoGOGsLV/6Rfups596k2k0CEbfGh9IIFVtWE4x1shkULz7Q9dlAfBu7kvPd+3KQYZNcIJwg0o
It8lNfvD/8AEU8WBjn1cmUcF1cjFdIhTpz9H/+eU7pmVVtK71KnybqR2BWOFpbounmf5LNZcmNIe
aHur+H/ekMFbGSTG3hl1B+XtaTUIDSF3E5efJ2PMl81uyNQafq5nOs+g4aGt3/LYpgZnICLdRsQu
KajX1l0Goe9uRgRWBV4ZoiKWsZf0u6gv86tjNve4m94j7ed47n4h9i6dMBcG7RgmyNk8S/QxB46D
lGRnfFpyWtgs3APn8Qmn2H3MAOAJXN1r/v3GSjBgBI6Vrm6E9aEeC8aUJhQ2ryAk7bK05PnyAG6x
MhGHZFXzUMAgSdAlSs/xzbYWQ5lIdctD3H5zVm1wyHr61pSDnKW6prMlLfK496a5dShM2ZiHQ3UA
PfUh7NcJa64tynNBi2DSxNBjtxUX458Wf5Nixjzn24YEajhBuMpEXfNi7mO1+5lQ2ow+WptjTHkf
l0za/TW2vRbIRofoQpZcPdLETvPechIuTL5pgfkRh+S5KQaketfDF/UhlPI0zDq+KM8QdaRA4Pze
djOlTImU2RYdQnaXjhyBu0cWrcvHiF+lgnFlpSlsXit/6dDCGCGiCtJMOWjrnkNvniyMsCLtdlLZ
r/38issJObnH0hYFEqdfvBlviw8BIIrWPQp1TgBdLXHhWw2RKqhmJ/v+EtElhal/ljUPxiEqSWMo
PvijjutNonSQR42u8fOgxWm+mpEHdIbQ5TlHMXvnsBNxCWaj02a53cYiNxCyA5bJjaEYtqZwRI5H
3wYgqPkA78uFIXwXtwEHHOgHSPDuC/M+8S+ndxgGeLfnjQUTe4T8gHG/Q8whizDSdGqQ4HfR9953
pfTXWVgmsmMxOtCKiutfFKmkxXwdiVFskrTZ6H1S1YGiEESN9s0R5EXHHcvtFaAKzpxuHuC7dlRU
cW2YgkpzCaiYDvLF/hzLaEl0blXWjT7C5Z0uwDYdkoAeSAN+KVHRqQT6yGuBtYaq8bIjpTrZAoHN
smdd+FgpxBGQ+IYJtDnXil3cdLXEIg6pcP7ww8tpU6kwM6bq60iCqT/azOT0FYOPnzXlZaLa+U16
DVC8y1fa0lKd9qnlvXpykFaD0o0s0VSgSEFS3R7fPrFw22mtoouFUS8obNSEzZp2kGu+k64COEi4
UOtrG6K37T0fiORxtQXPTfRG1plvPX7MDVweuhprQjMygiAGv8dkDtFnSkcmRv+2rvln+R4Q16Py
ePuQMAo9nWEgeGfgKQov+egxI6P0CQzLj1eJdFMzd+mejcfD7fPhXTB9yulil41Av6MvpZ1mk1eP
40V0MMcNO2mYCQIslJt8qsXSG7QoHTQoDd3412vCNezX9o2icb8+fx/a7y4uTf02SjH7iooBLu+e
GKVS2V9dh5A6/lw6XrXyryb8Jj2UhVkmZ7ApDoPLS+kDwdYYNBdMpbENJR3ZE5SIP/PdIj7WB6WU
E+8DcuWj7N3tEu3RI3TIJ+IbkUXIQQrl2Ql+eo/mrwZ4IVgaRqeCvlhSrYF0jtBmRP9LTdOuQJaO
T0xw95jNCJ9sOi9nM6H7gx0M3jAvC/2uEByyy38qUcRVbV2+js4u66mpbIH68+wXmdxWWSd+o2lu
zQUsJ1u5fcuG+NS3MSGzzU3Pob/RqfFeUb73FVwCKGF3boRRF1ENk4FlHADxAKd2xn/uWynQNUe4
+qVGVKWobl/bWkvHBTKtfivME62WTF95vF4tjVYCXbQT1iLBDC7POmScDNncGSxfNbSxuirgPpV+
0aeZDASapIArNEN39JMv4FPsFkGzGuTGQPd0guSChulFpBwrLM4JYRmE9FA9sJAQ5s6XzP7P0i59
ZnHPoTUegoAcDPLOmlbUHLLiXtzhkrrMkl7iOE7zo3t7LxuSv22n2XYHecvC/j6BNEgyafa7KxKu
U6bqYY1PZltYTUjZR2oHq4eJV6FM6pA5lJc1QTcWzuuVKpG/Npmv6WAHUOfCO9x4Wtf1w0LqLYFu
AyCmxi4+m/JODQybxB+4uDyMJJXh+S7WgeBExfJh9PivrJQSk50uT37H3WKsChlQJ2V8O0xxxw1+
YBaDuiYuR+RHmLmQlvE1jdPIrlbxhorVwKPsK2q8uMjHXS5YHZxIC+fZjcCGfvoJhIG4uPRHKqgY
cv76lwgXsdkeGF37whyhLsx033Q6rkHzlBxu8wf5mG8rpSF1zyyQUIOO/+uwxFcbROMgow2+OF3J
46+ua8Ey3kDs0Q4xC5AIb0MVLRxgO4a9nSckBDbAToTiea4uAB7wMDwHE/vn0aAL1IzZ5PGr+T68
JfcNBSo+H1F3S6ha7fcX9vihRPmFfkSvV7CRS13wVA7cS3g1he8ztldC9lm8sHSpPgo47DtyF5mM
GR9CEGD+JkcshGt8Hs8GOq9CugHnUHK9c+vtkKR4A+QEbNN7vuo+Ew79ZBbiHB9OPKYyll7/zpgr
7edIn9kOapbqz0XFT3Sj1iA9H5sQ+c4QMN0oFUXHsO/GO6Lmzu/2o6s2Qwqlhug5C38KVDkIjvbo
5UvugUsqj3gZ30pGfVN/0/4n3xX+uV5BJP0qjijNM7pvlFwlV+cwSs+Ha8wtWVwnz6IHTnbtwJrb
1rW4Ap9bU9t8y8Xpyuu65rk/tdWk/gvBjK6q8VedX/dVfnfEqT7mFI6xYDo8+4ECLov7xYcWUpqE
zHGQU1OC2vW5GILm2MdAlvaktliCTn+iegS8HH7zEItbtVUPIMZzqZnI1gv9cDEkhNy2tY4rOp1V
fidBK6o7jkBlV8gXTE3kmq8Cv1U7d64Ds6buhlNG2hGNqrL3CDxKlKD2M2fsRVJ1mO29LUsJKowZ
JX07t/jJ/jD4HidUMlndCGr4UgcrrKeupG99Z3efFpDnufuNaxmC7NoZ46qxQFXTP6twzqC/64gm
K8NxUjAQPEuEgPdMMqIYyEXEHaX0kV3zIXPBdT6nxk4Y4MVmnI9QfNSffGki4ilbghw2mz2AxANl
3VFuO2r6BbWsL4lG/B9xgRYX8gnycNYJsX1GEUiezX38UdvGDHbN2xDRlg48JlE87/6Tn56wVqmv
lH7JsyWxOD3zTlaWfH7y5h+eZlbd3N9RNW+ZJN9np4CnsZjqNoDWVuBMVDdDUpj1OiFvCv2W+1KC
48hwtcKMMNxjwj4YtDdFgGM1nUB3jsE18WgnAxiF7nIuHLkHBGmyjmtvADuevETcsix1982HS1Np
V89/yuE+1dFiYE79Q2xfhk0+HdNH97rxzTFOYIIfmWJOoDRFltpjE/paiVfCGOWjPm5giI5xuBo0
hzR1vsn+944wcft9U67ztV+Zy0mE5Az9g2cZr21QN9uLWnlPDnTBqAEIxqy0FkwGd3TcmiydV+kS
9tU6LYtTnCLa8dz9CSRtQul+55kMppygkoVzp/UWH2+8HA6aPFS3mFfGEY2CgMQoStCfybfZFN3z
LwBud5bKHZa9rXIaTDV0t5TKCglAhrJkCVJ5KSxpDW2Zs2BAmIZxhpV+kFdH5glMUn4jnpBsYb0q
9N0DF/Ez6euUwUSTeht6HOJO1gNIGyOx33kae88x3x9mBsd/JHfFBmPkqrDaR6m24elYvrPj0VGb
V9elyNNUPMoR8VrN1q8w0ukAhp92nWgGSI8ijPlSWm7YYaXG4AX2yQXtt4A83t5+cZ/BUQUxpcGv
/CV/UUhMgqNCCTUeHwR8Phd0yHlkhyH4hEzQCcw7XgNVdfAS+Y6DrUmFwHXY1n0qORy7z5jplXkE
ETDz5YLe4xnp1rR84rQIudn2YmoKNZH/GzbdfJUIw72LGXQRkSBpRGH77Ec7mVF5uGQMd/EBbeTk
hr/j7isJhs04xk7IlPFH8WpZzK/Zi12AvwmDhUrFtr7dZMy9Sk4NbW8cOLSzDpbTu+BPYk6o4b7H
WdyCv8zynm63MrWr6+Zye4dYahcRgNIXyVhpPFRvCefm436rB1rVQ3Odv7t9hJYlQB1WUWoJUKWL
Lu34vz2SxdOg+h3oXnYbxY8osqN65CovrnxYatXYtDNCNNsvXra9PTCCZHVHR9nIQuPAbmQTMWxt
1QFU/sVcjHdtBrbuLVDDLQfiJhNyXBpLvtS1FzGUw+rbVPzuH2wkjURoX3QXFM0vIfkFERbCOTNi
6xsdJcdampI7kQz+ndwiPX0O++6NRH1//+ckBbCiPUnKsMC8UFoAkgeF6ft+6xLyBOsaZF1tK2ZG
57StUBuDQhkKRgmuFlbQhM2GiGAZ3YLJsaAO9TCq0pQqtWU1jD/uxJryPQpsK606acZ74KSQxr8R
iTyq++j9Avm///fIctU615EQ8ie7oxwyBN6aNmA0Nw6KNYtujVGdSZoSIA25YIWpmu8Dr0g35Nqc
vopeZ3dO085FSqmA/PzYChr+Vg1fVnDZyrhncCqXGb7TFjQ1S3QalJQI9SS4EVDBz48YfUuEXjR7
88UvT8URPrPZ7VQw18joowNvIQqtWr0DIAwJuNWUH+z505/nohivf+WzJwNAOGpejjvgiUvL8mkB
OMtm7sg/NoK5/IHAhu253iP8ttUC9LmA21dEXGDEy4O70dRW3VNC8xlOHWYDdemLXVhxD82oEUan
uXoQfVLGdOU+V4XH83DRMDt+PLJ76PE0jFAgKGNVFh9ZKCXkW8qLGP6JLSWJNqfvffDCr3EGiZrY
zFThrVszL/TiudFQ+FbKA+bUNOAf00u6drSr//PjmUErwdjqkycfXwUBehdlpdSpVcZzu/L+zk7s
HVOWF32x0T3WchalN8bRHfHXXv1S4UhEE5n0UVwijf2dagVdde4glz2Bs3p0/dc/wXmLiJ/k1KjS
CWWfKAkNGCZVpyegPikShzZO1fQVb1RMC+Kv6WWgZYjg7y3dfZ2+j9mOvGwkYDAVA8glwKTm0+az
vcADS9z+QLAVKGOSCIfFZVF6KYUpr1mNju6iAlMbVXqphbdTg+FVP01o/KCSDMclrOnDko0lZhcx
0IvlDHbfkYOja+hY8x5K3wzYZn3lU6Gf6Ib9p0Y5WetQwkFZvk/I669IKKYs8sauw3+F+Djcc6rT
acr5CTLOoqNbYn3qiDCDr6oFEiKC8ra4UNj+cgGoYd7w0tL7LXnpOtHKZEM7OWCh3R9kDI84RHsn
r5QgmRI47LAcKhiuETc/Jm31lyRYMgyfjDURXNs2aqeELDo7O5smGHCtmKyFl2B43jB9bu9tZEDJ
rkzJKKazaZFcN4N1AzuTRosdgHGLNxALqQ/ujib18uLMw947QVoTGaKJMMyQ/57e2hLvR/ZI+hj2
OP0S0U5DsrjUbKUWilf7bBZYVl2lvp64J+BTTByL0qa9q/uPvI7aMv415zHYQJ0rk/u6z3f64FHy
4ef1rPm3sx5pNEXTwart1jsyDQzDxV0hP6VJyWrit5hNjaLsNdB1eek/igMid03ynaBRwbzKJeGw
kNm0zkjRciDuQRneYnNJujl1qxrfX8BIx31Sr99cW96rplqPPuZtxaCEkt1nwnm8ihIMfzuMENyB
/tPT9V4Ux+DhlYy43rtyU7wcov2LmJRzPH2PmZuT2w6WKb5Jz7PF/Hxq4DI4B989m+1LdVRHzlMv
w7xj9CZbTi/zuDleZDd0EvUwa/KPx7T07ubsXuJtRuv4LWg07dbmGsDyxyLNIrnCsgbn8g9CdLYR
HOWmhCi1Aivc0Qmb+GJxlL5jbWbe3MF4LqVs+U4+4ioJaRCCmpsirQqKEtoJNkdOjEdeWvKGI5Xb
rIrmgbDMrM6jGhTBnPH9ledbBWM7n1fq1H4XzqGUxNM4OERf/pQAFJ86YbyOKw0FVDcKqSAiDg8x
DARmZ7hUVW3EvbKmdOKnmIFM/KMEQdB8DqCKXwzj47PhD1lhjR7vZSTcEEnl/eTB3M7NCiheHMAg
ZTd3p7KutyslpEHmw7UTSmbtYtoiR94ABdywDED3RurGDE309li20cEROW8c35WjFtOWysWEZvu7
sZemXMM+q/Vei3afVN5BbmBarMjd51aA/pXM2y8jrzuyOzdZ4NGWyFIB2wz7Ewdrtvm6Fvtlb82p
9esP9nU61Pc4TvdpIE4G/Gx4rvUG199qnld+VxM8vvXZkoToKQcxpunZXb7OF1LdbMhp7pblYDl7
lmSpSc/gbqSFwYFqSPouHCbLmj4I8Hq2FHB9RGIleOlog7vmu7yCWRYpTzjMGWWNsx8fBzsg9aEg
/0KWsti5p4wXn7a4eel+VuWt/4/mVbXC/MBz0/x0vTtyTAnjo/mIQucWEX8cUurYAmU36NCct1q/
oeI59d4izj97EHgKUPMIm/IMkrEoEU19sffCPQ5tpw7lNe8ycfkXQiuC2eJg4j7YqoCEXIP3GCue
Gxb4Kk/tMSsZArrtrm3mDvpkBhwW1rAj+DcuTGo2/uKXtEK0m/SXYZKUMnzmom+kfOAKZcRPAK2i
afumIKIZbeZ/IWkkMgTUS8WJqwzv7TRGGpQ+XM2SFKC8D9GQu5lQNF8zORcwdPQJ5Fx9M+6I3GAw
z60PIiglle9Fidt8c2AjKlEs+EQGxa6KK4A1OTqB4VfozCf59EZZ4o8c+VyHzE4jR8pchF7Nv2Cj
HP/3rQesWmXyPn/78qd7vNrQgOd8YPSCtjQfCdeXLa02/oRtrUcsEoCS17UEcvzdhqLOSMSct6nV
uCQbQ4dHD+8dmJM4rDVSb/ABR65sjwMxuiQZwZkQgn0J0Q0dWuXZ/6YBg0LQ8pjRowAlH0LS6rgA
mry0nuecvTTD7VeAlFAQPAAu8WThQnmI7J+hCJV2ZtPIlyBElVYllsK0g9iMXO3RgX4R/RJ7gQ1c
pr58RQ6LWlAv/RSj8taC/NHWAYrFtpxFcgu/87cmDqugr8MNugMLEtspkIDylmo+oDrRE1BL8H6L
aO+pgInEFIGJLFgwQNsdjI29jJ1aTz6FurTkIg83yWp3YZroUl5tG+W37sV7dVSf7MxALgk6gcYI
FNHrTCutRxET9EIZhu0WpR9iK4AfUala7JXvUBWLs5BgpvGPd1Ye6muSDF9T6RtJ2HQS3hQNFrVv
kvnKDXPsWXGpjihCVTPnz055DUACr6GKiTtfmYDjlTn1JgdLDqS+GU01C2VfFl/oBTxPXHipoHOe
1LNXiM5GwmIStp0PCpvyY5619e3PjNUyqOWHTMznxz4FGRoejJhpqgq3Mz9yNQgyNFppN0/mmbTY
MfzhT2a/6SxiX09fAcqPysFrCWu1TRmPZEaPmVTN3nh1WbeIl5tUZBO5M3eC/rreE4jNOChr1+6s
VtdrO3KFInq8LVK5cEDb5kwF26c9U2zT2Pfg9dIp9snBTuNm6QEuArhLpDLiPUxRF52XyaBbHbAe
LVhkxpav/y0Lc9o9dKObymaxQgPe1ziMB5qCNct6YbwU12/3nxQBdgHVehG2Y3l+OAHDmnJ6bb6B
TK4ltnY3RKwwMkWogbP3pBmwU/aptLuiT7UW1sc4fGC0ka7UD7ZGOOWq1NuhHEdkzySd+r//ua6M
Er73NgLl9VREPyAnTtqqJwif3j3jPhlJfbgLyoTTxEoMwUZK/hnpFpiCCdq2xkF2ISx8G19VGNxg
s9hgYdjjpzBP+ANsMxZq6qXS7YUawiSUt8Y5mMKVrnQvC30wjomfWi916kTW4MV3WB1EhBDaym7y
N6tgd4jHKgRNiWbpcmQBFQy3l0f3FJsQ/zhRn8wRPfcVR1bPNd342AkybL1Jr8oko7IfsNUv+qGb
a38hhp0gcfCxC7+GOkBRiCEn5pScqKfk9vktmoMm4U5EKsiDy3BYYMNJXfZ6KBMqTkrEM2CTGP1n
XB2eSkYovr+XRXLQ+WOTsyCsfEtl6fLUUNgLJGzriAtnxqBFVMdVvd1GeIR5scC2vWTysufLg/LB
61QEqCZxH20jJEjZATTQcf7vJywe3pC9tPgjYNr6RKcMrdzS4/7wR0qdj6OpYdfe89JFtnoI4COt
jV+wOheJwoGEehnXVb6F62OQXQ3otmiclCA0nHAiEUAXi5GGY4R1tn8QVXERSTVdn8f2/IMY2OMP
Q+kF1vvA/2lAyp2R117xefCdSzebo+oqRNQgK/rjwc/jSWYrLNITJ7ISlLqjLljD4gW2agU3mq/0
xfF6Z0bJD1hzroQFyQWtAYv8w3gm5/MIWFkINny2mLPjZYdjmCCA1usGsSAeK2B2qkNMQo2Pgvpg
SQL6CuWgfWm658vHE9JxQWHAW2m5OwTup7D6W6bNSN/WCGNoe3X1O6YALhR2vN17nuSYMXFjY/Ob
4HPbaew/yNP8WM0nAyU3FY+oar+89HUG85YPIpFy+Ahol2oOsOb3zQkSqaiQfmgdxn1vqCxTyHdH
2qSe3bbxe06J13BW59QermR6IuAeYqBvqrfKR3DSTpCrzzAO1n+m1iLb5jJtRU9+fPJHk1yKvdQA
jg5x49TnNusBx4mu7k2Z9XdrueiJd48dCvVpdEPr3Y09pB99icJSFJmz6hiVO/em35Fgniikw5VA
7UKnF2iPAbNa/jqERlX3r9sf+TDIzvMtqyhj690Ul/RZyhrnSaoyNY42/iXLpC1u+hRziXocrPVx
YKsAPMKWvHTxHADHgqmh+/aQXEWRaYguoS2PDctZ4xLudS328XmO/GYTN6YisUjeLB8/o2DTdQgW
c9ijlWAhK2Db2LO9PG8nU8uPB9BKmm0n/6fikV0gbH2JpKkopN5IHiPx4xiW1D93Buu35nB0aOWI
EFYELf86kzoLF8MMybvOeopHBPTS5gnTIfPPb/QRDAwxzYKE9ZaQa4mO4N6/GRwH+GdOn0QOeL0R
bKSh+HhcIL2O1QJRzwcMX9ZWrfgZLZCNNG3C/tZb9XKZEqco9KricWG1MSgm/XDh2DWjhSkTeKnO
SiWPbJr3eG1vE/ntrzwXyo2r388fbI4ZVIPWEFEo10mwUEYHWks4RIxncT9ZJ96SZNgQhSy79cno
G7scGNR0E5i8k2gZwvIAvu7LsD3vFC86gN55F7oM6zNeI8KVoWtKNR6ssKfH6tdHowBySSC+T2PG
w6tw1VkMQJBMHs2xGHob8jDi0oxsBqU/O6SwpOg0UWOAZ54ZKp+hM++eS6tAamdz8TKmyMyWS+Xr
6i4ZkG/wF9mktXoUAMxgqKGSBlJpX/KMKaIoMqFnEFnhrRhC5tNovkCXweosGt31/8/R9GjR9vIN
eoWE+4nxrQSY0dpKwD9LZMp40mSH+znOyvLIvSv3K993Bv4I6qd1Lw9QaMW/P7g+IzBObb8QPBa7
Z+JJQSLsvR8iqirq2j3GMMaRMFnIw/OU0dRBAVF61CVwTyrLMVmMIIx4O+nQzwoX2I6DXiuFzZhK
CmAEXXkHeb96SZdgNRC9bKEm4ZAyxXMoFKPfpwtxIeDKzKzU4CK2z00Y798ZYt9wYHN02Lc0OO13
3s/5umVbgkIgP4YnaHIZtWKG8fbCAKa4KL22Zflw0QlE19GX+BJbgnmgr53E5BygkEi9jPGGithm
0GsNIYSqaX+DN/E1TivxESckAGFf4672TIgKOsauJd6+555FThD+wFuRuWDdkGJboPm7dkaH41i1
KdNZHIPYU0TTuTgk07ZCtlrInR2fpsxtLoailPrZJM+d4FLAKdhYKzMRu10bcsrlShUItCsKDSFQ
VeIlKQzLvNELrR0TS+R+P5xgkTCuVzYVm8yPcf3VuIMP0xJIShQt8Fex7v8KPVA3AndtfENjvEun
heeBO3HG5GcJq3C5n2OJplLTx3RnZDWijPrYXvmPv1keIwlJMdrshbHxIF+YbstK8LPd2RRfABYB
kn8g/szyvJ7ujdEwDvs17jGSsKXBXPbWSVPmgW9vavzHP5pVtSYrASYY4yNjwu5JBVW/2xZYK5t0
6YEIJ4VwxnLX5lolNYgDJ8qoYJGcxVNHxNLhK8yVzgrKMqjBbDfpA5+pKMe/wQlyy4ix8We7yrjH
UBzGommb5ZNPGaYn7+t2netKZvqm0SS2kc26kFDm6qFNIg7zgQje9ql/cGAqZ+CKYYBsneN8OTgS
yXRfMRhb3c4ZFOevNkjLM5nno0hpGFN/1OOZ/QSXni913NBzsOHnQ3uNVVT2UqWWupOsGu0STd5w
cPPnlreIcZYfWHqvbuUFXNIpf9Oi0TvFhoGLYbjxOd6zbzB7LaGX00C+dnFkbOQVdlhUwN5oFbnU
lyJdqQ904tG2aTuFfLJyMmj8B2PiWVoOlvRdqKf7B6CE0yRnrJL0pG3IJjzySaehEoa1ae03NZbY
WZP37JaGWkBtyP49xQ41ufWYWsYP72voGZ4lNR+56vkCyum7GHqCXN9rJJxfLbv0+EUESUEOqwOF
cJ3+szZ2Pxl+OXmMpRscJd4EXDUnEZqblFg44vDxh1lF0Q7C5V9HqWajx81nKL6IVe88O0xEDD5V
sGF7uae+KlV7Tuba6WWhYd3/5rkiAvjIxkf+IKA8EdgBiUgGaQEdsLHrqQegdj0ojGV4Wa7q3t/2
9SDM32tBgMq/yBBBalrdhLcDbzs5P6h8/3m+OX3X+WEfXqzJj960D6ZgjinCkzPaHgZO3UaSuAnE
XIAkiO8rt5C3kVqa0JogL793HgCdA/6RgNwbmAyyxSFhvvaBvtSldY8hkM+hjmbt+2ALyG3UQrND
QSvhWNjNLmbadLVdoku2GeYVXADy90rL6SUKyu4ExbKNL/Xz+lHQvHtV8UFI8wnHOdwgZwIan2qh
0fp7ZyEVZlAI4sD+0Lww5eVrGYImLFqmRXskxbnGdvkc6UuqgGxjViwCVf0SfrqaIfWzYRst3PV4
zoL1Nu1Ubey/6sLY0uuzyk1WOjdKRYb+uNBFosmBLB+sJcV6EzKnSl+4XZvb3sXD6xI1/X/yYe5n
1K1+cJkSY0YyTgrv2FeWYG5kbXn7p4RUhG7kfpp3Ih6fKvuv1c2hkPjSGiC67vQeF7fFMC36Nh0n
FdPsSqnR5TiRj8gtf0R1pG/QrU/oU7oSSD1nykAOh9/OwXPLZMsT3+eBgR1/ACeRaeBe/XlWprwp
/75F7iJ9UAUYQCDqxMnl9uM1CTPVLqQqgdQ8THO8DFopLscfMY1KDtG/tt7cJnGsbpWC7gyetm5a
37T4Nn9kqHRjXr1DIjczWq+AtFA5ePbLlZG0RcJdHYwVLoKZhHsSqzApbuomWAPqU8BWMjM2UHtU
I9yJ3c8GYw9eG44t5EbCifjHYFBaMqPuwTS5k1EP24yoStSj5xbDyeOWtbcfsKOXO7MMC6knYkme
0RqN1lYSwh/V+leAejrpLVnSzH2HQiROkotV8Bby0LioidQu3Z1AsidEO3v4yoFpqcmJRzd7oXsY
xas8ijjYRUgwem+ABDwI3KnBiH83TQkYdGNQa421NDi3pwkTldaWb4YUCMhFC+wL6OlfLFicfHks
DiUEMX8tc15bvnAwms+UcqnAfHT0gARIJ2vunrp4z2YSylu/FroGZK14FGpQPmWnHZec6s+1MuCr
7S6dp8kQOKRuTDNAdP24swchdjwzIyVg8JydRE+dzakgZvdnwWE7/xTMPsojMnfAG6JF7J+JdHta
FLObZwO/TMdEWlVDqya3trZfxb2M9ELJXtTgHsMn9lEBxQiBRCBLk8AQqHSUDOa5aXpbjqDpdfPh
W1GeSqbFAL//XCs9NYk1NahjZSvg5n86enlkeMAxI4BPFriaK9ajqaFkVQgkWQOAUxkPH09i/jti
fkWPFzlIOC6cLdzxtgwtYi/i5a/cBWUYXNDeH1Q6IiXHlc9OgezfJM74R3Z4KuR9D51qIAkhcqje
az3UOoCeKq3lNHbuasTMwUQwre9p7FrAQR2x5oPzbme0aHnBwLoOMDY7MAcjqz0gkI6NuIgjjyCj
FyipoqbRCUVyByPYU4gubJ0kNk20OhpWIVF6WgSZee925xJAb6G6SK0mzN109cpOL7rHCjYJhboq
S9HVxobkUsIClNxkCOYDproVRykh5nlMWCWoMMHPXcKcudU8AqOwgY6hemLexhRSHBuSwUWIBhTb
RA2IgatcQikOICYVhzYOYrQ4ONiGFq8N6DjABcCQ2/Lvc/26xEB6ENssiVj7Jw+61X63b1L1kThk
CwtkxcHfuXmRcN9XAE49DRQ9O45JBIs0pPjqqm/OlWjJze85CtZR1INe1mxEkIcsxWXpheNwZjXu
M4ENNHrGZHLtxOqgnpWyYixHY0HT/OCgpguEV7c1TKwxUyryLh+XK+p1nCrDchmVwSyqz8koAAeQ
WP3Ef4cCIhFKZ/gmnAw2VqLnperQ4x6J3fjtETSQ+9s6Pu1uetbV0PnX5BjORDjiDbCjklvdLYxq
JUmSNmJo/y+a/FahGtH1d3wnDVbaAi7jKVgfQhsJzd4Ndl1RKwcAO0wDLFR9rGN6xSPgQCdH1QnM
vTj6NHZrBZfjSecPA1zh02E9mKtkBokp5IgCaTvf6GG2Msi+FYv0/KiT5gJX7z2maXTStaS1vmfu
whGXBkPhEHPYQCTWlKFpB1TtaukeiKGDEJggzLvFuS+Rqz8RIqxQ3CYf42y2a1iOPbX0AuA10VmB
95fbddyfHqj44KPI7xElkgekg9aHFsET7E6IFEgaidowmYlYBvYEm77kpxiThZY8Kc2hXZ1u2QFg
nZwIIrcun8+CQP3yBMkclHQMe/9X14DnJ/A/n9KsM1uARd2875dZPKlCjpXNPGCUx0btTn5D5l60
sg8sShCCDT6KcD/6T7+Rotqw03eNnWPAv7ehnitxlQ0LhtazBw6fDpiPWXcaF5iySsq1d/Z7i+ZD
gSM2ywcarmzevDAD590C+tpq7sO9MbFTnfoYV7G8NjE6sk3/M1dBpI1YFMsJDCCeKaaxQ6l7kvHt
MGhThzlPc1tPmMFqJ2giy2ArxJK2cDT2EdsQMa48j4v2Z9eRY8DAJZoN9gW+dxbQOTyCd/of667Q
kekBJjxWAvaPFO8AqChq7u/S8invk8RZG6OIU+T+QryizsvtCaHceImvHm4k6Bg90YzPegKMdfA9
v6fEe0S7R3mmDCFystONHqM3qJA1MHkZfK0INAzN+fgGVgsFt/u3YhtcDwJMRlc6VAe/B5npoEwX
1HAH7dxk+N9bURp/RAxCLa1yTtngLP8ovjno4b8xIrWC29NGp3sx6gfQvYFXuIdd10LpD4R8NFWg
ruVO9M/A/JLbB97nk36ko9Uu2c5mbwlpTf4PoncpMWz11E2a3gvjf2xcONPe6Ouvhyt+a5Vq9awQ
oi+s4y8EGNWr0I7HtAPuimJFm2s7370Uqvlk6ImcIyhBp9M8cV+c0Jk43ArOi9mnFxO1sS6vF51p
gJAL/GJoU47oNAfbZZRI7xnGtt3EMiRrLQLnnBm/KtPnEg41GGWbRdTULFQo07Q6bpsNi0hklzv2
sDZGYJzwhgJcGJhtW0a0lwfh1OQy+2s/BjEuq757/8bOEs6Ci630mNJnjFhivBPO75UQQEGt3lTx
WKfYubPlkXZC0ml6wsb5GxHafeIV+JKgbjVx6atiTdC6tmn4BCfv4iGf2OLyVfY3S62FOScUd7P3
4q4xPIGDFhKPh+hd9iVQs+SfVVJpAVW5hQfTs3aC4HOFOSUAPZzVlVNaa74VmFa09rVxVvHpRpke
+NnEh7rYn54bGdWJlEuPE507bQoQvrWgkN+qnsyrhaDyf/Be1oP/VO5JdMZdIRSju3JQ3CHgo6SX
yaYzC/lndubx0EUUEFwCdAledP9UBuenkSiZa6bUxHPwXVYAjI9d2dkEk5raA2guwPfmVFqwTn11
mFHzsJY0a2NIwQmuFpPQreoIrTeeT0BbvLDthFeHG0V7bfWk10xHlSlCtxBnImCx4BlkKaJFvk/t
nB/+xztf6AFB3ec4Gxm5mf0DjgfCOtJz0dZhTqxbeKK4R3S6ubQfqF1pKkxxmLZRohPahtJf81B/
JKO/0mbXJRRCChwGwH39o3LcBKS633RwjWUs0BYWDkBL5LuS1rikLfnpD0VwbxUDOeczbg7aNhWw
ibOM9FhJdUVA2ksVRuvKmOckzBKiXnYt3F4VfCGkPe0jaEf8hGxi/gLeaH/E2UgKo4cZ0ocGefQ6
mcSRu92vgbfWpCxVEFBB/k1hiX2XvtiXacBPoO9V1uIZH0zYCNnMPIE5LgJ7JLhpVG4aaEChVf7X
yhZ3CKeKugAPBxlcxpCGZbOv6OQTF6488tTy8PUwzVSLjF1gaeSc/Cc2cXQnPDUjWDv8w1ZJwYeK
cICzAdcgtehOQOsK87PRUhtflQUKs3xMQ6roQFRa4rsrVnp8phV5UdoqEBaPbHHOnqbcGMcSOmOy
PwrCBAYDApI8cAFugYxY2K0+hKei7gm0KSw3MYfyAjQXrg+qzb+v3X82XfT3LAtNGsZ8wcMUu1jl
6b2LONDBC+BsWLFZ/CuZy5xp2sLZvXWWon+wSxWNFyaGe3ovoaShagXeduseQtI8jg4+KSjGVItq
1LFTz/eng7l62hIECOgnJhyGO+bDEm8/OGAjROQvtlca/6IVE+IqvsoLqQ/TnIWSgej1gaqD0hpz
3lH5QtLx3oqxDCNWG71OJ+1lLeDYpezKglePm9zHS9KE7UT/IwP1CKDjd61nF/CaNxARNvlsk7fr
C/mi58TzDsOWggyywOv9Hh2Ggkdgthm1Sa691kwz2/28njhNhWxHQsEWwXvvqUOqMqbB0IK5P64F
+Rlv9NIamnOZcnmX4GQkSyJbdw382NTz2XrH6GbwAvqrj2errvHkzPVe0QUNTdd7Ewel5d5/p2x4
+2ZQms/Z//Dki+XCnnwoCVFEl9xlNoqttWuIldXAG8/88vxlLxgNJx8/nkDDP3dv8bGlcadUQK8n
YIpN4wow9FWifaFai6ik+5bWav/dwDNLa9vqTBdmDLLHNwyp+9rh6lEWe5eC32zr+fD/FrZAsVqu
wR/S8uMJep/5lbn/JiPWTlPtY0pU2tpQfEfcdoNQ/b9KkA68sSJC58eoyzcvr+k5U71TNobQsoqb
KzMa3CJRQVb+ywZn5Vf+97aNXwxqJ8+dLGQx0UNUZNPG2h8QqyVuUHWcLkUgCmzFuUxjS2rAzM7h
7o/sal8eG8wmF+iOXYgMKqSk9iF/jlXvnqLJYu/BGzIfhycFGixUh3WZBa6iHwZBC3v9PWh/sP5Y
4GAQ1mNweh3n1JBu4H9q5Y6aV6QV//8SKgEku1Sw8q2wgVhd1YPMJni8QAI4BWRLI0ilSsIGkyI1
70DjV/VzmlKiG5FEZ3rWvf9iHS+zrD7lsXXEcd4fbJhn/BF2QQf99nJzUv5ldxDTIp+BIrPjikv1
oa5PHlq/WyRWKYW1zsFRBS/Im6/AVxv4Bl08aghFk1Scfi22DYeg9gZ7g2s8OZyfTxaBXyFOZmY5
4o1eqen417PpF5ckOhqqkmKUfb8VI/vFMNYpM38n83PSsSRx5aCgYm7lq/MMWG5AkuHIwc5FR6f6
QALMkCSs7HmSt8wgDyLvL9lsOoC9nokJeD+OAsA3GHwTJPw3x/XyHbN2hlbxgBG7vTG/gy2Zsxx/
+/b/7IAc+RW4fep+CWsxvtHDvJuOIrCkAqYCScXK7wcAO3uPSu68IU/OzxW1dPE1HFMobwLFG7xp
J3Me6M9hHwFXik4jIV8tSUUkup0sixfyWHNUouIAKdAX6l7BH8vOUCVKxFditBOcuUnx4nZrBQL0
d0+2MyTMA8YV8f4wVZHrdPW/P+8T8i+2b59ekSRvSVu+BA2Mk5pm51F2NjI/ieJwsxHEplRvldDU
jPe6RBtfndIawQb25lTo5aeth9P67BJrlv1MclpAOqizWKlDGXBxZbOMH0sFD7cv47htEvkDO8JE
uX00GCj/1LJPL6YuRzu/ITNxldKT1DROP69Rc5yATHzqihqKOjLvw076qj+orrR5iXlyFlT5kytE
62i9g4EF1HPgiGCVhDHwqwDlwnrTa+2qlm4+xK0RvoCIOfKAlTsDfuCi+dOCidpgXomh7jsaS3OI
aAw0Nl+prIzge9AwvjAU9GXP7FCddv8xGKkvUGFCzsbrPIVwoSydZ3DMFcOVrx7VsOi5wUO0R0v1
8MyZ1RY4710WtkLCh7k7+0JPvOHeXqUh4e7Ry7yVpUsHuoFuDWjyJz44XuZy4uJRII+V9JVJd4XO
6LRzHaVroZQj7PrWYDGSiSBEHwmRp1YbilfelOEDujJraZhd5AaqhfMbjo2dQQIvn8XoO0y+IaVv
SE6SyqqVK6XWdBGTRSLL+cSIKWGEV9ayzQa2qrhATipzkZQR2P0MTPnUteeaOkX0kcTETcLolBKe
MMhYunqcZF711bLflWWzJ0sTb6hJc8IZEVOuDvgvNzPjMSNg3f0kT/8i81tF/w21TVTk+ut4xWPt
TJSqkJ8W4f3xdGlXHgVIyG77/JkVFfiElA5Xw1jtTVhda0ag3FIUNVxq2IHgW37rhxn/2BjSSIKU
XFOrR4TpKD0g8S9QQTliyLmBBLrZDdBiWSm2/xkbMsiy4iDTsCJ9Xjekdh9/yo8Ew/5Liy8Ft6Aa
qVXAmZ/pxHA0UxCucFKdktxPjTesHlgYzBpefxm3CuKQRzIO5v9ngT0dXPJtH4ISI4ss/JBowEsk
WEhs1tJOtiF/dLZ8thW4YWd2sqgRn21gDwIqufeu2Th3Ty/jDTg3Oa+X2iV8nwzNo7cyTGshENR9
9acaFrvRF/KtU93AX8Q6D1nnT3epZw/oGjTm1w8aWaW6hDwxiyrZH0koLWjRoTASwmyEzS0UoGiN
FnE5HMnx6z9Xif+n4erEOVfgc5UXgR2pl4fUDeTGSd/07fIV7fCI0Pl0UijvSlcLA15D3iXVKbcl
LjNzM+/iwqtg2e/5yvMJzC3dRkOz306XjnLG6IwijdmhkdK20oQCX/JoNdE/+1iXvBnj+qC0yW42
Cuv0NJtHAPyyBVoTIUWzqBExwHkMFTaHYGgx30aD065uFscI3XyoUQMU8dXdROaVu5HrhNa5HpNc
VlAoXeqM53xGFA2dzERdD3Vo4RPqOibR7X/Od/x0jOiRi6sV5CY6XdD1rfPBk4ve+gC/gjF6lisr
SG/d2KC5Tr+h3of2nXhLo5hfCfaO+zBEA5R1UFVuUOlxlLYd03Zj+J6Wgi9I4DIUrWBpmFSQB440
kSdv5l368SXSk7myV53kMBaHoOYs8vxwGF2huElhQNzmlyVSqXMu01AcljWfpHqKGXh4ghBl1l+Z
H2oxEoWzqNJ0VNOpvyA5xAGwSDrsZcAtFGpOwaEsIN8s5Qdd6CifH7FnKT+376AJRVzz63PbJYP+
LjTstlx5+5YNSZXLyIZ5zNGEN07yGJDDLt5T4/UIfGFpyuGNmDlAa3Rl/19z4JXcVl0olRcOoJL+
RRdW91iVtLehf9jMSTHTf4srGPDJ0iIl9yikSqqulSVlxWwAh3juWo7CEJwquV2FmvMBwMBuw8P2
MG32lLM019BFJXDsfaQ5Wha6N3PfPO8I8ZBq5ti0KecuTE/AtdbkMuefNvrFrj9DVMmwOmDGVri5
ApVaw5X/C2uMMvQoQztzwIYK3YvCgUKoW08ZqBWWAQzlt/b9j1amGq3NclHUx9aIeXcG+/4pv236
DcD1wlaCY/s2XPd7tYXSrdXJrOQc29F4y/NT5TngUg9woUydPjf+1xlFTsQn1v5hWMjahvyyCCzp
/paGQzWH2PxjWolc9vN6kqloW+hTyUHs/C6V0LInEU0nuRhlP6Zg512oPiQY1Tpcy3/NkanUZOct
Mcav1+HNRo3Z1xZmXxCgt9Rf/APrGwv+M89dPLJ9OyKGLCNY1ZBbglQOgbhK+4SQOMLwr99/G/7A
LIsPnnOVKjsb69JKslYTgYfkJHo7semjQ8itDhCIt4dVEUVATk8Z6KBdOzPO3Q9arQ20DfNvF2hD
00qadEBSxR3IVaYD/OFVgronmXppnCP2veQB5eT++WQ2jvMCRQHYUXmSzgDQ2Mcd9ZTJmgoS0Erw
1wQ8jjPDYmOww3cq1kLYAocZKSPhwUesM2z0X405VZeRewqhczvkuiJbfSlD+3C/wQoLpb2Rmxly
gpsn3oJsR43wAkWpvkSx+yxxiVLq1JiTwxgfFg8f0GF/dCPYxcp+dip1e61OGVlBHDyobC+U2lNN
PSL2zBGWZfRyppT63yay+MsStFpptDJSj5KmIP0cevhOu1sLRYMk+Jm89pMMbx5FWUbb4e365y3Z
sxW51Vt39Zk72xOVg6Vcai+/7FwUCJhqi3XjD0kayrw0WiHNrsTTcl0FKRwCrSzBKvWd8PbiPATn
gZpwZT1JXe187bLL/3GF9jKITxVMfJlFzha1KkKgj3Iec4T5HN0XTY5vxa16vH2Wk2MCSBA8/onP
938Ys3EVdjUrJOb/I2pFvs9PTQkAfgp5q7Sii/eGlYC5ZzrKRvsPYKrsrWWCUF+zwsq96ioJukpr
LbNU8Xq147NxypDsdCJYS5mRIWrfzoPZnka40awv7xFlVCi5D/JyAUus6UEUXLUnRgF00kAUhFb/
y21eVUF3Cw31vCkp0i2dBnHB9WsEzT0dwou3GTg0k4VH+ftG3pJOc9glvuZvZNeNeLqQCztoa6jR
uwLjL7DjhyZgw1whyU32+GvjLAXiAv/dOuCA7oyPQsgCydWUz1iA0IOpfZUBTvA3onGu6pLgqXCo
XiNGIIs13bu1HONlbqW/t811erKuF13gELsFO4CxRV4ejji1ySf5HEYHkhnL3/q06Y4Slpn+mWTe
xTpRBxwPIRRVT/XiI2YLlgBye27L3NQyZTZB8jAnmGuAnurzZ46Gm7UjC49rlhNKbZA2O1KYFGI2
MOeJBrECrFrQ8bqyUHoGTDz+hlE9A/Pu7pANcyh1mPxFojFbC8jI0fberVYP4VxX1x7/QmmOXzdd
0JeUjydsMGkZ7yME6LG5uYVETjQZ2l6O1FOrpxdHP0Mt/5Bj55+f6rHMJtPwkZm3UW2GX8Gg4Tix
m0KZnt6gImgt11NoFCMYD/8TO6Qu24qNRl9U4xlHAvS2s6Yln7sQhegcKe5p1u6p/49+iZNWKEU8
p9PhWZ9FXCl1yfSOoBR8gwovpFUEdSCazfgFYTLkboI8MgTuidmtB0gixynqsxITE2LORCTavt0M
QIY4xvxrJQFE0hKQkOfbe11MirvSihpoPLB3x1STGcR1w7xm/QUAdLQeXSjNRdE0qvhde9IO3/w1
IeluBbr1wC3IO/rRi1b0txGQbpaU5tDqe4sKYWiJDXzkfn9iIIajOfa7wzRbzq0MjQev0LqiOwVP
b+2i95eZjo4ySMCkGSkMtl0XLIHuf1x0zyr2cAGwQ1B0biMiVbv9zvtavTrv9seklPYWCy4ALDCj
vsDGZounzdGtb3C6sw9jfvsuxp8oHV0JJpCW4mqaP0iJ31CPjm9TUlaLoit2MlfwEmoKVGH7A9k6
4M0EXbhKNvbCbuhha+K5fQFWyjxV18GFopZiAb2dfYRdPHnAD3GOqYxxdVjrkr+J3q+GaEA6bO+K
XN0SjA2LxXB1mFvKUw+ZhH8SH1LJfzMCAPxpIvvDhELzkiqZpNa6a3kZAPRzguqQK4Z+2PnNGZUO
1XMK70XDi6aKTT0DgvmNkxZDsLisA4BOAcVvfBgnRQlh04cUjPHoWbt+YwkTBzxvCIaqROw84dYP
eZg0IGCtLy5VjlSz5wVXxEd9HmzwnB0vtz9qpQofd2euqkxA17E6gZn6Qz/w3063h107qfvqJUew
yQOr9n7EWdTwi+uyrWOytZHSp1dQjG0englatx67l+25lIznfEZ4B9W0FqG48FzyCIX9x4mwiCw9
+7xPNSERfZ+tqhqlV1zO3GSqrkp41/G1lFMx6Hw2HdCWkyZu8MoWnDQzILUGr7AcNIKcG2dLiMtJ
o0LKZbFVgshyAmj03GrACdTzN7SM6hluFEJB1rZOjI0POGriB/U67Wp8d9/mWnV7RhDQU1s/nVL/
d/a6Q5ZjBQm8pfBNv6F+F4aJyDFk9P7eBXJEHadyj8dyBVjfEhvZV3lgfEuMEIqa4ZmnfrKuCAJw
ZY70utrb0/dLi9z3OKW7W8VbdEBeQzCAVV6AAS6xgN51uNAlUMfXwTAAk7WiGlpPOok5ZkaI1hba
ursG1QMQQMj2lC8qVtr9TWV684dnIqGP76OXz+It7jmjEqZPasH9WiQLeVwhC7qKYQAgs5CF0YYc
TBxrFU0I0Pw6WynjKn7JwKzTRdtcTkQfqpWy8XPQE6kHKyvS+V+JuQFyoMK1jiAox29B4YmnVlML
yMqOWqKJqTjxcGZ1QogbDPVCt9LblGvT+KMjp+vX+fromFON4UGMLuRtiXBya4X9+GYe74WV/WCU
C+nDIgctRMEBiqVf9ksVklzYvs04RGKNDKQCx82Zx7Yw2523Ze4dKudIq7z3u9fuFknVbkFs+4eg
RPEnjqhtd7WqZsn2D+VzjonLXbAALZatcWYeR69xxRTam/nmN86SW7PrkaIwNa2w1nl7jdF9187o
8A4dDbUp7Y1llcdgMqcS+7ZJhhchzEPRyDbwSzxm5Dyp+C8TEYmDO84Bpi+5D7iUDnOzpUo3V7Wa
iNwqepZpoUF1qnCAhXyidHWdnGy8s+Ubb5VKNbZw647/2a7Odyelhz2MGQ6Q5v5QEFgYheVZjckZ
2j4xHsRLN2DQvsGv9tfmgqcZ6d2fJHXmdVHRNSCsX4eKiGPI+ksKMJaPyTl9HZEKDq8dO7hBZxix
jj4VTbNNh9NskQ1vHgKcggpf57p7cDq+MeMyunBldT8rAz4e4LpA+3GAcqfDOd/ZUfNmJ+gkA+Uy
3m838rK+7O/YeTYM18pd1jxC7TEu6P4bC0L0vWcnpV9ZmHDue4MSA9rR1sJg2xo51s244l/vbCPm
YomIM4PWSSQo3OI4aZnOluVsCTMDHGTjKA/Mk+cCsNQI4yMPnREAxJpVYEA7vDFqECklzyTN10oS
rcGEVVM/WxLoEU5FCZIvP6z4jV8E/QKNeNJYi47rwRR2ee+m3pd/4kOML+Jt1vq4q0e5QxMaLRNA
RBzaO+vZgIysxzgBsngU+4x5aO9nMiTf/X4BrmBDqRD1zBaa8OVTMc7IfxWUaRSRPJIVXQh2N9rp
NBjFk56ELFRLe7pDfOn8HjT7w4Psw21qkWHcWMdFAXRTBtK/votyNa2qEd/Z77K2ZriHWYTxwhVd
y/RqOMpj4r9Nmhd8QiyUkkTKIfIUoCW8HtK8tiCwa+lQjqPKDXHww900FicmZAUxngeooFttCh0a
oiSYlhP24XOHoJIbAvAoEaxeYXVU6F3kN6SC6E5r9iMjWYSfA1dMhYQs59RgQ23l3QugWexsQky9
d6WLTYzxRuUzxrrqJaa7CroxljJUlyH3HzGqx3Zu7gMnbq7gJbqCEsT/V1t0TqfvonrbrTptpfTw
988c3skFMcuJsOhwz4QFZFZ1IxsOxUWXZk1D0YASYH0FYpyRyScSVerqeITj78SL3uW6VRsj28cj
Ee8CUmlNdQgijnKMV7MLTkpxhxMRBN2G+CPWFWgzB/AuvEz/LJEfY7MOC2hUxIcHYy9M2pP4vZAJ
h+4CxzjnxjfSgYYrejGuBgfKJjq7S1zRE4+0D4U+sC1WWtSh+QHcpvWmbdg7EM4fzuzr8lMUqqFZ
8D4tx49m0VQPrthm5Wf57HqViJ4mS4BNy1jmZPTlEd+4ShdBRq8odSE73jfgUZZ4W1NyAamTA3/D
A3bQTucL8WV9DJUYCXFfulnbGFElcsYwXr4Vd9CzomaqnAf3soQx0+1j4XtSZU5vsHLu1GogJ9C7
tFvpkWOZcV1o4Hvgtx+BHqveIquXCi/xRKfmK1WJyvrox/80MI6z6Ve/TfqGiUFido0AShejSL1R
6Eo1g0rC23J3osUJtb95tSTiZrl3Oteseei+hory6KiqX8FeVqQGyZvDGKWJd55wOeW/WyMjHAmU
jMNzJdf16yEsoBNbfxQ/IJXx6rQ/LLCgltI+dWk2dciJewRSm7IAYrSp9cYTHk2cbV/GDB6IUDBL
jl77IGVMbMzHVYD5R0GcdANGRZC9p1hmnzn9PvT2kTO42wR0U0+OnEhrzS+EHZ5ZQFi1hHMdpp8e
/OF2gEgC0unnS/3VJp39A4C4WyJd/0yaKktF57Ob0k/DNX+hPbMAbuVq8z2wYUXeHziOHteQJMyb
sIj0D0NfuexaZKHvnj3nZz4AlNNnNQA7A85ulbWIRdme8QfHJ2D668kZQLzBLFPQhS8k9b/9S9Nz
H3B/dSyOshLI8PRlaNVAwU5IrleiujUFDio0q5xc18chgfFBuw/PPe8x1aDO9qiIXo0lw3jqM3Jj
TYEWjFbQNkE7pEvvIRj1+avuB/nZvyHD3MrNWKYIvQc8HGC8eVJsSRVs2JbZ7JhXx54a4uJk0xp0
pZisKq2wc1Qb4KY53kv7ROyUTdHr0Do1dJxvzXk2i51/1ofXp/JfsPjCPNMII74QJ3T25p2Xo//5
/4zomzhTdEnnvyJLbdhJWCZpfWh1yNH34HHbfSDq7ZMrEIooxdccxKRgfKnTFNAhGKQLAKuFHS75
c3EOmFqlWu3hh9CJPex99XJOB4JjcS6wvpnm8LHT+mVC0Vt+rYYqW5GPXTrWQwW6H7Jyy8g8XP7g
poJbGkNAFPVHhmWraXUUCU513GI+YIVvlTEq97TIIgARWSYJonR6QoQbF/Eo/zp+FcJj9Jix5pGa
S+wiglUU7C8o99VtyJgXNNDxk4IFDxAV57zblll6CkML/drBmFNcKR1R4G2PCwhLjE83JoEPQMtT
ts3Zxj2bQVNgD54/0S95ystk8HFEfRddZdhZFI9J7wpATDw6UNcvOeWDZmPGruy9vzd3EZDXVLtt
bacgqfxE/1DJ53K4kmy4qCmGQQ/SxyzIdM4oEwrKiO/lFGdqFAj3ZQdlnVmsb9TFAoPL073U2LNx
X/BHsH81zcIN8Q/mXTR8+DKJ6uEh+SfpnoeY5XAi0E/fS0PrqoOV8g7sMunpwjsY3+jv8x20ygkl
dBzPCpJWaoW2V2YBZhGKmKHbR56LGNfhpty3T9fGqHApP4J8kucnT4lxiGpkj4mXTnQOZYnr5ATK
v/dI4snI9TkXkMj0s4+mt3honG2chCstLYUPqnhxC0X8jcE4shVy9C6oPq7WpwzGMgFzoCaAkJjJ
vL0AvdQiDVHfkGYxTGYFt2U3jcxhvtXZDf+5qFpsiYPp8ywW3DVxkp37ypzg/KIT9Xsg3U/2wEPO
TYISKHbu+fYlY4LyeTP5mi7T4dMXAq0tnvbwxOcmM1BZaxXuZgBBLiFdPT6n8JNdioTbyK0QNJpm
lcxZICY8rgayAuMQHXOp+v6QsshxWqnE+1K/7Yqli7qYKqIzH+z5m4xym4HR4/AMGF5FHGgLY/2z
0MZ78TAxw+QmuC9lG482Qri1cgFFNiL0Dm+4ivBi5OcJdM8QSehPFrvPVSAvZuaUJfvTj1Dhd2wS
BO7yk/jfHUIdm205udpKqXVl/TAFEM8HYKh28Ioyttvy+Nr/76WS9s++vxh2JM0m3ws3LMkyn80M
dZXEscG2Q7ScIshGsEZPkPqSWKig2R4TR3/r2lC06e1RvN2OumOlwX5EmZfS9hoi6Fy0L2raw0DT
XNvPwkIjX8rJo/7BXnn9kh907v8DEoICi45JZC15XfPxO28w2llGLLqBPiH9aeEEuNMitu/xULYO
OPHQlFH15oV94xw2+bsY+gXxyqQ6jyiOsJPnhoeNGQK5ykrHQo9Fm27e00Fbe2CHCI5AvTLF5bYK
o8J7XbqPtoVko+IxDSNDw9A8tIvtD7n4b5w3F2Ox3Gtj9c4JiKWiVezHmiah9ZqgByFa/jb0yw6u
OPVzKKvsOYDr1S31NK8A3I0lB2yxUFMRz6jtmhsA3HYQMSUodVhsUAu/oKqzpz483ZV1jgIQ4OFe
4NcYHkSDK+rdKE4zVmHwWIKx9zIVU2hQzpnnJMd01Aa9lb5liJ81bDqnmsoxRr8N3UBxEW4EGUg1
dEPiC7JHlt8yj2UfPwij66I1tUVQUVp+sDhiAheJpnvBTzjAUG4pGgXZa9YqslpmfWRy7lec4MKZ
WeOqBNQlWbaiWlAnzMiUOEjRKdiS3+EfZpN4jvA/C8JQtrR8FcMnK+wGX9aNZv/08mphV3ED9GMj
Paj2BWPHGPZ1qVyoX1n9ZggCEZRMp5uxbxciT2pJTeZz5y17AkLokkqGt+NvcXE0NSwiT9fjbUPm
aA7bSnM/vKN+o2oIJURd6IiShKwlpNhkueOj8/4/ZT1l1nOjuOrfurpqXB5m/7iYSmJ8j7xZuKNR
d9qjGTWtWRYDYBlZE4diNGI306iXIn/8ABbluU8mCxF0CJLJDPsUE9yJJbc6vMoK8bjma2Ar7Erq
rutLkeRbpGTXUIEwKlld0hhQB4nra5qAkFZXzYQmN2SpdbSasgI1Lrs4XVTxW1ht3sFrQU5Zlfc3
f1BaSowmiamllv9wRVPXczqUVptMObAHX/s/Mz6k80w7VMeEMCEmU/7wZ+ZFvTf6Pb7gB3LD4JB2
wzrajCiOeUh/U9wZa68pQKTNXmuDArrX08AQDJtnt/+MDzlyCxRYQrSOXRhjMpcoO5M0ZhJrGEM4
DdDIBoLh0dWji1hnL9XEzOkm11i4lu19G4yXppMlhqn/5sonTjdkfNgpdXQa5hKcVbkLugMCkmIX
rxne7SjzRPBS5KmMF264GYdwGbG5qc6h9HyigGMblztRlMLIKVgjdiMU9hqWLsDtrNXsUO+f9ea1
0GwC6fFH5a7nFOTxxaZ+xv80zF4GkNzoUZgEJNQgQ0k8Q7skB7qL1N/FEstP7cohpCHQg4fNmiTn
rENTS8U7uVZeImaWhWcIoSNhprG5OQOq71H06C8aeElG6if/Afa/4iRMeT4wtsp83Mqiu6cNFtka
51JmUp2VRqdc7ApHU91qJ9VA3Lfv4Eh31QD0mtgRkglvVTvhuWY4HCvK6FZluybTieEVJdvTsr6b
8ubsrD1qjicG1fR2bNBp0cA0kYsy4408cdoqrF7CK6qGSzZqyejAUMxxWHKfz89tOUxBDe5HJp4o
YYu8RsoJmWw35dxRxD3xHajxQh4ozZcelD10BvTccuTtjtyWNCSK8U6NFdBH7fqaC+ORRmLE+gKb
chPTYzPuqCwCaXQxeBvsi7SP/xRRdK1CATVwRrKXzzVJArFbRaTtmNAJDX0l0GplU4Gg/5bSo8dT
0857U3tGdb7h+T3lHFJBkURiKslLQNHS+3iuppBRzII/amr+FhRykTJXHxGEpm7opz6d/nLv9Mj7
DfZ7hxlPgII0GATfS69jnRKfNj/SQZzlKuX6HVcCxmlCzZ5JSFsDMNA0punja/MrqUP7YF+hD7e1
nwbKxp99uTZWHVFNt4b7dkE96UKcNPoEOqQ/Esh7Dh29DH8g/02fiqXBQmkm0f5PbYJ8qH6fiKlV
alLn74h/T0dwXcKogySwK7syPDgmdNB75ZSXX6noUXGfAj3wSVOEdzL5SnqfQ2mwYJe6Mtwyhxqi
MC1Oh2I4hVbGH2l2PugGXIOMmklRY87kb1b8HaO+IRakMMN3mfhk7ReSWXIabWGmPtmGtwJYMbax
Ul3CQJ2JNPPCUBTWIK4xCLce3GCIYFpD7aYXpoYJeUV4BtC7tJu4fVjNyTZeGdQWntCpJCo/tK6t
cvercOkDaiA5ksVzMv54EfGM0ziVoMmUVUgW2vgdIL+xmQ9mXH789948GLwqENlKvz9T6zDt43Sj
KE2MO30/UMODfdUrdHWnduUV/wO6Uix7UwwriUaoxXdptWzQHORU5psjqEb3vYmpQOQisRDo5QuE
YgUmWf+tMdVqT17hLDm2uNc5JCQHvZHYf1CFzd/n9RqmZd2zETvQfOyxhLsSDo7q0NHsoSjbpd17
nTJerTthXq4glBu+6c3FZU4uVumBjc+ZCm0EvXQg4yEqfFCjNoW+DVTcMYvLcWB0Cvj6L2rML6VS
i5Ts/EDfAOF4N2SEJxT/NWXvySYjE6Wpt+0mwj0AwGtoIqOsJIXyLuNDl2+A0gKWERRziGrHUuFM
wKBoGRl2o6SPKiC2//cvpZO459cwhl/oTPbo0/d9/SJ5soru1/hL37pppEwmn3goYaS59cf1w01l
0SaB6dYd06pL+K7BRCAf0Yhg6WPS07ghtsk3ULEqqd5IDlMxdzHaatZ2BqF3U0fRZLNXsALF0r8X
/WS44GT9npkgUw6OgtvO3XTRKR4JLdFHNDxJZv68n2IgK7SgcLbIfwlBOgU346XaPBFasc9MKEjp
7ufUPRvo98dFmJ/zMELuA9kTZsfrxXKZPy8afxi7UMMxT6UjAybo/ykUyxvE1OcogJ2CgpFKy64P
9CMBJplhHnbl3gA7EWo4uBzS8ADotU22+rfK3SR9x8P65N8HHIfqQDCPDxhsEV0UgUinyh6CIQRO
S0re0kGGHgeFgZdIJmgnKxegjp5kcjmuVOn+EWirBH+I+v6iEDZCzto4JP+rzibumQiGs+RERqUU
8cuu9J7QQjTlUQoMtrsQmPgoIgVeivYPVwvYJWwXWpPsofJZ9qWYK56vKZZj/pZCa6vvvRBJPjIm
EZRh6wtpa3CHQARRyYpDUDa5CU3XNiwBYBeP/GJZIEyCWrXaggO3PLN8B5OWlXWBDPkYOOxsenOz
jPCOQDcr9wsIiQsscUsYpx/IuhekktprZQpPASGXTj6kmQCcM7os6d+aQoaSJJRWVcR0b2LZj2Sj
Yj4kg3ij9i+fsIN/dfdGdupDkGQOVPNFevVr9DYrMdLEINnGxDuxTzRlycBKghkdkr/cTiM2brmX
bVpDxo84IId6xZ6TsgsnAQkUASeL+6iWznHrqbu5TMaNXzUKy3JFrC784rEAszlfoQlkaLxulqJD
+a2fa/ZYS+0LQFQVQjaHDshRu5Hx0CbUKN2gHFrwyYJES+/UGb3b9yJQxCh3g8+niwF2W0HJPjDJ
sclSLlXc0nVFDsqdwJ2F8zjyxRzRqgIBx00FjG6mUZYbue1u7/M5nD0SoYj7PTdFG/pX5Fjaj1ox
qVn5oxfKBOo0gjOM3TwJ6gvlNvl/hOlQtLa7gemC6wH/ovei6dJSr12ZMSKlZ9aeU1Kem6fTY8gY
Ex5x5ozzDhINrFJywnYZnAIP5LYEl+Wr0T/H0ApjgL5dP7HCbJmcQBi+weI3pJdsF2iRCZr6aDRs
JVwtZUWDGBXHn6NuAUWZvm6wZcI66iM0ld1nUh+ULvHD5DNDqWtGuFTHjEOHZiY8Oy8Jck+cMfPV
zxuAeVEcjFQuQa7sMzclOxk8bY6TXQ7U8QpDAAg6HF7z/fLbNYcMZrFYMm1kfNeWQ+9U0b1UkI9S
mJcvkVsownDiC2qwYmEp9wgtwYGjvkenEloTg/23FdSEpBkJlRjjdYiDLOs9SuZDzQhtIRAuMeOz
obVDm1j0mT8UxNMA+aHmUb6aO+7Xrh3+X5mTk04rRv9oiwlXO89djn34NJsYjdFwRceKiA83vWyU
qjR/XW40jl3iqWUwv3ERwuY+FSygYBmf+a9C8o/htsiS14UPFUzqDmnez0YMdDXvij0Z7/dtcu/d
ZFdHiALmJLsbaopfpijbnvfq24aDPtTfrkIu8/FffwaEjbLV4rLqEDMI1LmFy+03preidFtdLdmZ
sLNIatxNb16wbeRZqkk7McQh22g4Q185Y8KLzoUPE6Dlh3R8ofjPUE22+ubmCDEmZQaD0o+oyFMC
Fq59NGI77a5vtFVvbB7E0coydF1YiKdD2lnBFPK5+RotFTvnhTyhzuG16ks/Tt2i/52u9w9kQdsb
XwE/KIbdooPkFcIBw6jRQUAwIMmYSvQDXGeIAxWOXrRnhpfp3asAKa2V+JJbCOSdKrvUoycaRUj2
KGlx72ewFyo7XnR5gUY/aPjk72eTvf9k9dgvCB/Ihre7oCxgbjEN2bZf5Jy3EmoPd0/bUJv7jwWp
Ogr8rP+Jh8U6QeJmnRRtYqBEoJ2QepgsNAfwxhv+IsGMYf64g0zwGdlniDdll5GUqZ/YFiekev78
1L2fnV3o9Dr3WdR8y1Yd2meTkxS4aRVlaVmOgLF4+nYAYHaC6RGfRDE/D/oEO0pXsO0gIMWylH2c
MMPg/oxN8Sln4dVvnilbtno40bFfN6TrfXT3vm1OJEGNGnwPScdHhVqBQBsA+cZsAfXrfmr6M/HM
JnAnyJxQjooQOkv6fikiEnM9thYbSzn0x7FcptsTpZn+xkTCTSH/1II/hqLZHX76Lec+qeALFHiL
ng+bwDtV/lD7hRDxVXAUkYZVCEhn4v6/tQfA8LlHTl9ejIyB2/OPYy/pGjYsHDF8woOYdGalAR9i
eU8U1/Vgyx5uHRci51SX3jF4CKkjSOLID2907lj5px3zwHQsxuKZPbdFVRhptu2V5LHcKRIuBrby
hHiqVF7yzVfu9EZjoRGAhEx4O/95T+Hoqhv5T7p9S9KdHEJaqRED3kCowTbrYp91ThCd2ouLrA0H
UxIM/x20o8hZSEeO0KjJnSPstj7AO96IpotMsI8Ttrmsu10u4giKCgji04QByaU5G3r5nFJhp1U9
Xu2XPz62XBT5an8D/UEG892679PhtWuum+j7/ZOVqomVjj0ujSg3+pSfEvQRwvpkLNMDbuENPPbN
6oM4X2DCIwaavat3A1x/6IeZ/LLqdNNZlyTaMLgae891Q2dOGNr+pOaenUI8/FFfUWeZWZ6tjF03
v6t6BkCOVjbBADSTYeCl+VDziPpAc7FKuD081iXIao3lLJI+H+BhK8ue3Uln/Tuo07agsNA3VYRh
LfKLf4+nxBqHjCCiXRpYbFFBIOctjX+B0TpJd0azh6PnNqNMhNvE+qxjTncVJKcmcOfOaUisjE7v
JSb7mgmRH90KarqxnoFg83NDyC5QJ7EDPpenK5t0TB0vm/++whOo2ng9zFOBFGvfN2qI7IBuhKJC
IAWlYEmzE0tEOjlHinT29xaQlxaUv45+KILOfDKnsPl0rD5EQWgZsY1EvVeGRt1ggPir9/7WMY/B
XfzJfstoLFMIwWb6mYjBtuVCkMRvgbjoJe3qv8bRYzFiktuEFYrRlWUFBcBS98XxKVSQt8YvPLWe
TVmhajpiUlhXrOlUhiWQqESXQb/J/OjaeExiQ/CbsOHvh+EY7MeOsjoldIyWEO1eKKQKyCPID9/j
6QdBHxXCqT4PjuyV77fvk4qz+q43CYmz33DxGhNgucjxytR8sl9cr4H8fdDMmALhDyV/XYfjzhbJ
buywwKW+dGMEzK9p7KXENCYweTaxrCMuPhSEL10KItkD10efFGsaSjyefnedDFqVl6t74J5RrR+H
zNsY/lAAHG81HIBt04wQ+MwmYZJjzyOYjE6+GVBGj4yzc6O8DlzUPliI0nA2HxvD2/Wvikyom/iu
Qy4D70aCvjnVC1Pj2Eoqc6UKvhMCr0OvfTByY9EU1whUDx4QOSQAGjfGT4VZApjzkHFar85P2Pfs
oxvRGUBNZF1qSy1F6ZGVdwLySzk+LL0RFsIA4s+eVUzgxiNaDNOZ09lIUTGPnzwDlhUkkIYelkjR
zYXhsnuQgW27QCoM4EohB/07mW1tFJ2ODeVT0yYDV52BpZ7vhfILBvswPmpQNRI7EdTMaa3NkIdj
GOqHiZt958DRGPWlAehUW0sBeJz9YxPwRbuUUKMfq0RTJlJjj8v+/VJR5xtUNBzHwrIo2oMNs1Po
yrkFO9p3TKlopMIrEd/RWSKqTkLxD40lyVpykeKv0KIuaaep5p63D//qlCWFu5TduwllO/Cchz6p
56aOG2Ub38aF7ZkMtvB3FBh2UIYrD1jamkWILTU4VZug3aPW8GKKuw45HP72QHFVl0rnSkQ35L6r
1cv5RT3ZoaxBTEDXGRT54X8XzZYotVXFHrRy3Q/IbQXeB/MBGJMNxGnuJHMoIMrbbFFyLBLXx4iF
ykdt/IQpJ7DXaVd9YjR8eYkXJv256kV0c90HhdtO22VHUzesT4YUz/sMhCKzPAvnuqqBlfYgtg9M
5nc7N4qPwxUOzP+tZ/9PD+5SE5k0zXRrFa6HleVRdCD/YvwceBG4Efti0w4x/Zqzis2CUusnB4tt
Z8I1ATnAf+CnTIZYL9hbgjtA9bUVkVlHF5hr3Q5Zf/aML8+a0dm6HdSvvXwpXUMEdKMlzXaZUC2H
jDzQpuWzriniq0brd0ScUCCdlpCaKlgbtrcSTD4n3dpsQnavMZf1kVRQS+0Bk56PYh5K6XY/ecbY
ssTmDVOoLzak6pIibShJLDFl8nTHB4ALyYvSazRaYTWnXMEH2HDGdOzMM3QwvMc2bb31FooN3Tv/
UMFTQ3qSPPfLRIlKk50Kkjj4HHnHYGvQOYQEc+e+pjMDdLdPpQIhHy7AYdLN7cIn0d4p2Vz9myZY
321W31PJrQrcZQpM6axN7TYLf+C8sCOAS1i2t/yRqOvqplJPKsYtRV9cd8xm/CrXconXCtG+MtDj
AGqQLi1FK2N+HyLAwdDaGMCXfarD60JoUQTVzWEqpJs8bkF/FG6BWIQQYgT8UWkVGzN2YYI9MeN8
HuLcsUJjKJajpRlRfhZ+jsFY7XHQ+/DVgunsliixIgVroOBUnryCMEcPF2B5vPBaathmlXwbMHXU
5Ii4+akRmd0fKFyqgIoYXfeAt6dTeztIykOK0xErc17pLOdu2x0LXKxImTXFNS0eto1ab5hjoM05
tA5Ig7LdsG7jNm8HREQcYrlQYAdceTmRaEnK2omC7m6nspgTxXJzEqjZoVHgfIgvQLx4+HXzCEz+
WTnBpQe1+16xihQJ7BPxU6B2qZjKp/KuBXmOWWOhY9yKQmSDeNC8DgUmky413+js4LJ7xGWnKnsR
sO3UX+RhJhWV9h5tdnRlTXQAMZ8wdBRHQ5c9bjR4CCxqAkRsZafIgEh1/85EPdHrcyjUs2pRz6RK
itCMhB16FjM7HoDTlWD6yD9j2Q7o/3VbanmxmbMD9jD8DjLMK9vPdFnpZu7tCjLUprn7MFuD8LEs
/rmSZEta71ipxFRQIIxXL5UfI6P4g2VH9efBSzVkSUz6PRiJZYBM3e+fOKZkt/7OiJkb0whAumrq
bttfk+u7NMwRCOK3eQ3zEN2rOt+UUMt92EPzk+4oeNxBKXmffetFN74i8/9LqRKMD8lpKB5ePnNU
tUF6m9UwVjgaJdFjK0wniywTy0VffRqvU4yr6HWK6+xSxVNJyboA9CUQWZu9Sqr1KQjF+Dx39/eF
MkS7WrpbPhIiqiV36rzDbG2YKZpU1VxU8zrD+H7TJ3S6MhMj9hl2fn8CgrnetB0apk3SRAasSRbj
bQ6bHMbMTqDr2omyomEKfmZ9vbuXFm9riyQ+6140JTBNuO3MxtxfKBOpBsZrFMglkkT5V8EqiF7S
NxkoB1QN97IJHVKrlUrdvTZ6tSoQQ/jAXn2W8ow2GGe+by2c+b10o6DeahMOcxak2kD0bopjLtUZ
9nm3AZrvL7IZJotaBXBAcYdK2xNeOOqFc/QcjrzlEATJnKVANLSzFnyOGThbZrdABb1q4yLuSZp7
Ibm7rg62HJQmBmizZTUaZweFM0itKJilkKk2hiiNLjXU4HUmJR7xzQEBWE1aLETaFJwDDn90bfX8
Eutt0fc7Ywpm88lBlLx2znVXXAO5xl5vx0FQXAqtqF9j7wJAOGpJUDrLi+xXAddlGaLs0/aOV2mu
bzf+YhCLdQTkY4xYhSaZOlrIXF8TXjGjQmPFuVLndkWlM0G+JD8woqNYnPeWDU/Wi5+hcyi/iE2r
lqJM1JtKPbQWA9XJ/vxixC5YGujCLyMeDZvFDcpCZIb1s2HXjjpeOgcwRjs3ju9RU9JlDDOrely8
jAhsR+DlturdXvdq4ki1/E68t5QK71eT447qGmH7cdiloWe4yaRXk0IVuK7OORVbKuxCbhWhiyAO
xTam57WSWNKHV2kVK6+GiVrvHQAj0jzhwz1CthRleJTJ9VR8l3sDtJmfwns1gSj30mmZbCXhqZ26
aSLuEkv17pvOXqP3SqAkFma9smnqrLYCjdxGUvm4bnZrwJNWxtIHPyw2PvQS02VA4Em0ZPFREBVk
AKJ6PaDzE9sD4SAA/LDIIpDWV0HLtViimgnMDr3jSN1PoQ596MJ9zHq0cGFSOJixXSH0OgnUwrnh
PtK7yrp4wzXigkCx+o3X1LlXEgFW54EXxOVZeuic72ILy/ZVCTtrthR4yGlqEGnqxYw5+mL+n9S4
IQrb+d61/I8GFWv79YWkBazlFbBYL74t+pZl7Gb8Tx5ptmuyrVHeqD4iCwRnrTiBgUtMvxiC7oVh
jgNDuFgPhMpi0RdO+58sXHlLaMbOCO9hWP8GMkbRYfaPZEut81e8+qH0vWnL4thx1QLnv1agDipm
GzGHKxUbP0OOIFxPZ5aPlG5kvTs6eYi5O8+i8QDVs/sFKk2xFtIO+Wl7OyYWrVjqyhfj4EJAC5a1
tPLehB5zPOYlvDin2IAyPQ5VNR4Wilswy3FWB3jC61Q40eBNCDfTPOF7yLQ88IpWZjCD2snvq8Uw
37pZ4OZH/Oqp4iQn/Mykp5cbWcXp7RxtwNTYiA6r4NyuP6m/16svmzmCtu4jmuzdvZs0A4ZSS0Zr
XKWH/r3X4uvivFio4NzUmB6ttSXeHBEnndkrQiQELXhbMC6DMR7A6keTYbdOjvGA8XSFz3efsmiS
uFjj/bgL6B9AB26VMMhENtxjAF2R0OvSgWCo51aSbdk+OlqiUXD6IXyHzSManrzFemL3dz39VNl5
O5FBwmtkCTm97cXBRfRhn6Ld4IBftN5bKOMkeiYMKfvjKWutzkPxoFw+ko75nUsE6c7hC/8mO00B
AUmQ9FpUuuXDnpc9IdOZn6E5yd6lIVdto5Nj1jzcr3I8fNosueUqcciSPs4v4PP7uYLilfAa6niE
SySbzm+0UjgGXBnlZneBw+j0RQnzEwP5ram52wSZPOhKLKbqgFR8MnXFsePDcN6LSfCwfM5WKfX7
GL1eHOJMPcL3U0YmRcKY9w/0RgxtjVNY7X6IqtXyxovpoKwAMKgt/JfR0zDsvOJCeLh88IbSbWTf
L+7zfn3zixTMewVZdEkp3tsQwGXXoiKbuNsFo6IC/oOXqPRnxUjMFjDkjITchV7m46KIoxcK581O
7FyNs8sml5+pp52FSaGffDadodnqg1ixPxGP7vRLzZhhiS8TxJUmYGU4aNC/1X/6W+CnulDA3NF3
PJfU7topNbVUaHBJbS0btSHyZ/ffwSI9iSe0MUtN1CjJySGMoj1w+Xzc3eN/q4kr0+InfLelT1Pt
TWN2hemTAvJaaVJemH8NJgb9law3OZqAMdmkinNjNnFXeR+HyqKVZlPzZDgoZoRrsXW5aOd8dgf5
wHrBxsWyMgipeyTtv/f9W5j8C42y18AFlRSxysuignNlQ0SQsFqSILYEAyGyR9FY7KCOB0mXvA4K
y7SIKrjVqm1kN5SNWkCMVFsZMlgSAz1Ha8K/lcGtAfcabp6uJfLvXUsyl/WH2I6Bt5g7N8YLZ4YH
23/jNIylrA0LRca75i5DbkUUuYpRgqFReTBV0uxJitYYVJO0YyvFg+28kUBHvO9uISIge9y3MmsT
WdvH3eUx+WkNehXmf2ZLTPt74ETbce8HAsTvnBKguD7Ot83iaCFNk+1XBJuQo1ScRqlDvu8P0PCC
CJaPWi3kTgwdR1f8+O3hWWBwE/5B8HbBOIPrmNQUpABZ0VEvJ8oYFC9lEa1T14e1ZHgVZivTmsSV
g0I01upL56+Fck5Ts0oSyr+7yoquwUFOxfYceefIgv6KAdeCrnLkbkb9hXFAthSppo5Fgud2awBO
PngvipRfuLq9dIOzMszKA09gZD00cKR1febzffnrBveoVRF9FikhCF7n7N3zf5ag2gF64SRa2kMO
wI/Ya9fSnEczGnG4X4ut38bj8f8oBE8R1m3JYqJdiD5cUrV63awZbwTZMU0xBVhZ8y93uwXdy3tk
M9cBhNKNMZJXkhiQdMh7vism9h1yh+v8K/cIP/ODR55+zxfvi+bR7CQsUKsSQhWuBxXx8Xbw8uX7
yIPY7vq7XnhltHgYquy9PZavu+pjL2NR2OE1/rzhBzEpPQM385BSMj1fR+RN5MVPPi3aiIvQkgdb
CJVxVq8bkIScvFXT1J/6pI+RRRhFib3t859E8Z6TAvqldftTB9Y3QFA0d0Ejg97fMsUtgeToOfK1
XLGaJ9djTR86JhcO+TZetvZWBgrT8bvwdyFsSyKRs6Ke27+3qX3LvIiouyJ0k5MHfAvXxU0hb/hE
bnrlIQSjFwppTH8Rh6nQ+DPfBinMB1pSsthart/B5nsjjBHNUXog12r54UxrUFDpAp9syxTl7itw
4mgi0jTdMSvnLLOy9Gg8Twrh0osDLLri2X+kSEKcFdwmzdo/lnWrzlUr6DEwpSqyq9HleU/NUDGV
PhSufxH57hWphHOodlJXo4QGu270e3XBtHw2guiJACHTPHEjSUaB79yFfr4V1yqWssFsrdPEBsTr
i3XPRF9hoCvOXhLWR5wDCbGONaKkEzuPyUjkE4B8A+6IpBlXzxY0sE0tgJvYDyEGj4tjHh/CIbBA
egbj2jjf+fkJRL5g6zidliVZofav3wn8288QJ1pxY4yeSdD/WIlYAPBbAGsDfbZPCo9dYz8VaV6f
AzBJwYVV3cspQpfG7ulgc6vnOV9w3jkKfFAMAxCDxn9DnDJRnkeI9DU5664Kex3qpU89dLeFHxNV
mPQwgJHlMa6ePRxYobE4rkf0VEJHvmXL5olUBtopNTaXVB2084MWYVOcYznjO0e1QhkMRhSjSXwy
HGLFP2iXlBIuYaQ4/an5YoVgEyzoLLvMp0cYiIgS2JmLt9Mlai8qzAiFYXPnTEr8al0+C/SEQHNx
Mp1Cs8fNkLPB3D6tMe4A7tH+dSlrSC1vsrnrnzo7IRtjiUmHfGK7A+kjFEzs96CkNomAzQ9kzH3u
00rTafdxR9nL61Lbi6AweWxXhuKvtOdIDgPax8TsMMnmtRHcG4COO+z5Nx8vRNLMBXbB1XWIhBbV
TQv6/0/EvquUQmw8oT7AtruNh/OstJIGFyioPntSFZEc4WC0A9x9Q/P0DO0GPT5hO7RC9V7x6M9y
T3GFNWuWiiyLuqkOmh2d9KqaDoALRGncUXgjo0zII0GWLi7kaCaYOq4IuDBKzC4CNbEg/GHRT+Aj
S+xCNCnB6tL6jRh04gFJEi6HGdkJ60KkMWqqe7B+UftK78Op1lQF0ouQGF7gpqrlO65Ybs019TAz
Y1RAnUPd/7nFTvq5jd6P3pyRvaFvZ18VfgqXrzlGK/EbL3vq799DVH52IbyTUZEuIbcIJyG93f2a
d2teDepxP4KaLMOazGlaQHv5qyJtV0AKJcFfRAFkldxn39C9WP1120b+dYLMsy3Ov35w6zYs0TxU
OarxUtBpqxfXXWuYtejxMC04l/XEHPJU/NlNGRwtvCLtxJ9XDdDG+RUSfM63esdZxpup/AFdSUtD
b/mGOpb+pfpi7OBkekVeG2lIFh281hgU5SIbzwuGDnraxI5CjgSMEa/w6paS32R2eTZT01CIbgGy
2RmkKQ6cYz+RYKMGvDxKi3oWU7I6QfRnqM47XB5Cq5dBGMd1GXPgx6cejGSMPzMkZ3Orad/pyDqj
lH98Auo7aoGZp/peEvIQY7rwd5b72rmSVKvjseZM+Et/cfmpPk7Bs0LnaiyxVnCmqf3pn5EsAYT6
RFXGmkDZflZBMHpzf8WMsOrgnvUtpypNuSG0yJ31gALT5CHGyUvq7zVNg1qIPZPZFbWXqsx8k2gV
0IB4AFclIgNdbhMydFJvLgwYSThniB3IOVD++aBy48Xsx/rVwAsDtCdoqcCkHljsUGGOe0IfNt18
ZAt5awswbm2r2MXXVM/zgFsUFzhoGbn1uRv+MtalDrLa5CMmunstbRWOvARKxX9N0bHM1HY43fOE
MHC7kB8dLRJVzZ3djwg+hgxKc10NfZTL/bRygHW4Iq0s7Gvyzia6XqaQ+6wCkSjkWZLaJVFIs68B
Q6PTWKKfS57hZeVSpVKmWV/p5qC4uFbE7bnT+G0OL+Fhl6cT7F64P3Of1wQY3oPlKVgCotDqC0w6
o4dK642CoJyEWSmdvEmv3hfORqwaTvnHvUTy4cpCon//T4iF/9u9MLlU4o/o37I7CMjBb1YWuntj
Zr8DdriOXBQeVTo/ScQnD2FVunBiU2v89mkEtmZnwOSh08N13faC9AILPP22TdNQuAscFp+3FSYp
h/gLnv04st8rPLYuSGncDa59vrK6eiPW+j1U3JeUvoqj73yDJwEJs+8YgD0IH6gdu/ZZjN+5Y3bB
0n4yfXBy9xcUQ+2KTsrGn+yd9yLPqbAyvUa6Dd/E+EuihOJoRYOJHuigUFimhjQm3rX5ROZ3Mtjo
hjBXVqqdn6PL6Wim1JRQjw+OjW7nIzfj+GOh73/X6teVb8XiGe9taDnhnCD/wI8WmUkfDjd063Fi
6+75M8F2H3mTiZYkFMoogImsNy90epabXLr2e/guDkFiuTF7h34cRHyAr+q7mLgiicrJWOcQDejc
qkECu6I5JynW4wGt/Spf2xbnCN0X3k2+8wewTxcFRxdnwN6qOPIP46ykaKgyVwBhBBHW4kQZTERp
/5bZC4f+gPQd6AJ4MH/jf1HbcnSvM1KKoSmaFmrlTc7I+eaJffIwMK1EZseZdkTIaf9QZSf/55vq
+Ayc7YNwJiG2knIFsyGXrd3VEGGoPl67eMpHGrZaHu3ZKMCEuP0jkutwlmJ87GojPgyNxKKbLu+B
Qi8HU7VCCamPi+CKWRf9LCtqhPTlZG3tIu9AEEcfrzMEI4OqXjOG/ne6gg5OiYJUqUsrpN4yEWCl
GoioxXjs7Yhsro2IGk+zK9I55vE7d1naktJQevL4Pa5qklLV4KoAjYfMYIgnYh4QjbPkqArDZHZO
ax5XYqZgD89USVaG/htvFGUcUHUXI7bHcf1cIE0o1pSnKWiiBldZe5qYevdgVRnsyYYE+oScqGHH
PATapXfAkMiEGVEHC6NwH2xgfHFvP8K6wuzynH/1aQBpt7TeuYjQUeiHUCZJaqIwKTdrakcPeDBL
fBchv5yAh6Ko0VydocylLZTD+8E2mtSmhNpKmV6jT6/1DXeGDZj7HclrooiT+5zHf4/ZgSnGjIFk
iECTDZpEYolbwh3LWzCni8luaee1Nmu2+inTPARoIOIGaYrrXrmAqTwy5z+Q9CLFMuWrpklhKYu/
vps4cxbOBFenNtZ3PNGXEqQtxOkN3z2yaNpmfipoDekLKZ3Y7uY0AYSGf1RHbjrzEVMuxx7YuIB4
7T6PV84vlAOOhskxdHBrGdtlofT2x7xvSATeSLaXStfoyB5Ar3tfxY1YAVxJm9apc5SekH0UaiSs
aTyN6gaPWoSGwbNHLMIo3rrzVJjouK971tQbZhfZ2fFGBfs5zvJkYpZW9hrKHZqvnr0TbHdUASz9
vg3QQWGEL0fvGmH9osc/MiJ+1jbatRC/+guhhY5Xk2v5868xOq52tctkGxWYSM5KpmZ9X3FQhWoR
ifwoqNe5O32X6BUawtaXYIz/1ChwrjZix78ceLYkXPNbMUVNTbhN964hI1J+ME6R8dlALWaBTUvx
mQEL52l3+Py1rUXYQ7Ers1+s2IQB8CTA+iTVRmAax+cepZ25nFtRRbB4XcbIhJhHTyfpzkqazofZ
49ZHebTctKhNxals1OlMakQzrfio0zjG1VCNaM+Q0w871Pec5+o4cxhmOKwNcnFfeLgoo/z08EGf
SAGdB6WSxt867F/R3MQJZIHUqmNa9tyXq4j1Xr+qdGl4zrIZ1fO9+hAHDqiJKDRUAKhY3HO3lswt
095yqwwpgCknJjl9Gs8jOd77ne8yY9tPPc9i26CHsXqvy6x53TGSHVt8ak8rwPujr5NxQurylOpN
pH1eGT2b3UE0xtkbH68ONERGqLCa7VN/FZ6RX0Au273b8QV+1Jv0aGdVGGnXXCfJirs9SgyrA9Fu
Vf+/9xnA9fmRsz6+7hv8SfAt22zZceQHMbOd5/uTKcRU9ySmMJFbmrdqxj0+C49KeIHWUhyasXD5
pNpQkd00kpfxEn0ad6EzHmPH5MA6JBD38q5vFbLVCfV0/RAbgRH+qpRlRTGY1r3WlMgt3itq0sl0
ft6NiCuj6S1Cf0pdhJpohEtgtdgRMlEi3/tY7sBPm0kLu837yAwFYIYbgQ9savEGgmyGSF1KQp03
mkJVd2hGn59YYi3FTE5OzzV0tTH2wYb5vTnqI9wbbplQVR8JhLsBFNYog2bBeGLIEDBZUuGTK1K4
so6ux45nlWXbhSUtSwlh02zjevbGaHfvk762rh0NQwWL9D0IKxzwf9MaZMo7fjlAne2iIh2y3I62
+NpNx3Ek0T9rU7+ogVHSu1M738yWB68Nv6CjVzHqLvpjHcyUU/eUSvV1VpoyIa43Qr+6Wgv5VwQN
ZEUHQjAPnwyHGep0wwJ71jduuA5yhk0ExsVX2j2K35aY87CyXl8PLdfWGPIYBFdZoK+rakX09t4D
DE0md6K3eXi4Ml+4FMhab49xJKJZTdjEjo+21aNV8Lrzgc5B0KpOiDzabweOqasbaso75Aw5JsYh
v+ACaRGI85JuFWjJItTXRDrUI67Q9kGmSBk+ooifrtpzKTFfBagR1ieCg/FDQQPfRieyUz91OmdT
aZU3ExnD4n622RmPNe6AUjR50gCLim96a2jZFKwqmREzUun2THXrNiY8niLmIyy+8dEtxk168oAt
3/w4GYqNnxMQKmKSTjmH5B7V1tTXGuCRpoeDpj3p/Qaoewvw48NcoD1S2QR+enN+7nESWRWQ/I1P
h8/MWajtRhygzR0sG5qwFW+6KasBSidV26U4czMAOXtmqgRTjzx7cncDWik4VuIExwVdxUxRtvKn
KjP0v9jTKLARVmDCYqTytDIEjvaqGJ8Xp3vMaWTiuWV+LCTsK/lave5mptk2DsMKvNrc1PsaEJ48
wCCoFt0VdYLtRgsFB35/DX5thyI/T/Lo+SAwwWj173bMGTVDgQkO6HplmsW8chdDEzuFnMa1OKf5
6Li5HY+1JMcXeO+5yhILKUjGOMjaEP9/joJzRH+N8DgmXXdKO0+GQkel+oalYsWdHXtMpzQnvDqy
RwZRH/QYgLS9Wf/Z1KFVRooRRhaOKCoqJK5EOlOJYVgn0QumJFBiFriGoZtBTGQp57njPS4rOgZx
jZtfpEBSYiYfI+cjcXTO75km5NE7/tOrMsIz3YuvbS0Jmcdk7ewX0OLleJriLSZdh6HkAsCML54v
rdhbHe1FwSe+/M3OnL0D6eAr1xnBXi9cPlTfJhga5OmMNYWT+jgsCdmHH7nk423vsNBnVc7bRfbx
mCT+DysLAji4pLwHEVOXiptJV/wJhfRk/Wvbnc9aKyK9y/1taOy00UEajEtBmwSVO4XhGblweO7V
jyU4FNY7Sq9xLTmmRC1aDrH+zeTgPkfd3X2tfL5L4EwNBbK0N0xqaMdOs9bjrhuS6PQqQvLpqqlM
yWG2z0wYsrriPKAcNfiv4pmRFhqv0QBFL8/iyL5sbIq9CEJ3nK7X5JpX7pMJZG42dKMnphZfqf1R
NxQwvIB4AAI7MzVNwUPAkQOSYWgieu9OrgIP7dVsQE4qNWDqJJjHEaGtKex1qBAq+2HQkRi5fb6F
zqAQRZIZ28GQIE9T5k1o1bkG2kCmJmA1ZBK8hQ9cYuhxgcwxEHT0yD5+WFYTTdJedAwFuWqM+tx/
5uMR7GS78VtLY7Prk/CXEQWMVImHKjaFPa0WvswJRS0Ynfs9fLPhZj52Q8F8zciwRLG/mP75w+y4
Y5OxtDCt7vnywqDuI0miRw4CSC4Ayy5NyuLU3o/XYrM8mJFcP5SP+HDTYM6xGPYNgj732XNA6QEa
4JHtoydd+4i2ytRx+tNLsM1ZuPgPVIom6sahIzdU0qkteAdfsqWsyJg4LOcMSeU6sGzCRGwwcpLK
H1UNUtkX5P11V8FM6URTBnQrOgPC8F6zBFc742MTjkJLvPsgs1LofuVSO96TB4HmQgebW0MnUH7N
XPC6rx2rUn2ICjpCmBYB2uz6jY72ow/k8BvbcyEsv40Z+MhKP+S3NDbvHKHUjakLmnuURLylrnFe
bqwSdekOPu1Ao2hTAxOZcmSfwEW4TgF3wNKpwh3Yrf3oCcXgKgy7VNYHt6ObEEqBxx3/iNSQ9s2B
u4bynF+AwOcM0W5+wUcp1aK6emItR8ZxMYHEkz5AQS3+xZBOlmyJIGFVhJYCMCxi7M10jJSpnjWS
wix4/CfhUT1tovV8yXJstfBVvoGjjYK+/M9pYIiz2A0JTCJSuJrn6UuUgmyF9J0U1oaocw7Td7VZ
NLbeiXtZUGFob1MbUy9w4v/KKvycN/u7oTIev6WYXvdLjcH/+yxjtCddtkl/+QOQUNk6crMYZ44l
LE3rNkveuuBSI18TjWC9vvcrPYpFrF+nw9Gbc0pdOVkqRHS5SWj7QGVT3VO2ayk3bgtexy1GOgqs
WkH/HyPBNXA/7dtNo2/4xTw7GNdlqmfLtIz9HdSiG/qxCRRs565lsLAcy6+qXYCmxK8RQWusfKCK
M9/LQyZjHUNvycsx/8qXAgc5fGiUZ//WJbE7WP0LWT1ywQdgJDoA9WRovozsojXiKz2M2lcit2JT
UxKlFcYA9S6ObzNHS2glT82EraKJFwxeF7QY/RJxnZ+H2IlKmnXf5NkUvZ5jVJJfqRxJK0MsPxtw
/usmuVCgiUMFjnwlt9ZTVE46eGK0k0BK9fzv1KG5Vq08U4oZQZQ/FZTrUDdH2lqmXEYGtxZ4CuWA
OWGoEqsqxvxJR6Yy/FsMMg9rz2fW52Fh59Nk7joN2Q5t6qUxQC5UldVtFX/Ba/zHQZvOGfx9kbd4
lCvOL0+cEEzRItOI6GlgxsVilG8k1Fsg1+GxLBpw2RoY5Ap571yQ5v9ggkFYgZtSakwOQZoCb/R0
n+9EgETHu6EinV9lR+/YE5AWHnwNDpPeNjn97o182W+qxLtkfnqucG4IhL5yY5dpU2c4ZbuWXXNC
30Ust3vBiOdeVom4wCQ9gEvmjxCxaeaoIQcBcAE1/AHZvSPXsyGNsf05Ivv9cJ5ww/GZRxIi1cod
KRSqDDRBpibUZS4VlQ50mhnPzGtGmr/U9G4Sz5TKE1XHCU/HyCByvTzyzDvph/b71rkMN96KHAwD
8jy2SrCxz6oSxqQyKCcRvw+37MewHMxCzE2p35uCq5T1VgBpTlN8UFpjYDaio8SycvNOTECzdiBP
B2LD2bIifriido5Pf8A87J9XYHq1y5aYH4WkkSfi3XRpkBjaPX/TMj329S30BwvekeWMOR2wyclc
pQQHTVKjm80LVF+W8CKzRnjk4IPGeyzEtMwxkL1Vg1cWJKLdxt11qS26+Szc3P/gbyL1PB01UOis
o+ttkpRk97aNbByXsedQEkLUpeslc4ktwS5qnBs0kQKKVwghQkerpCYj67UCorMcFsnCdiujWT16
OshrY7woiPQDSWD5UDKtZBUrsKx8TwrD3nmQ4wjKsi/kRbGuCrVsR56PiI84OpsYbNuLibV65aAR
mXmBdqvqlepNdD5tUd9HiQsza1GkoJJUgsZYn2RLWZonlAbqkeiuLcBte0Zjip78FUCykuaEr2/Y
sSkJdSOgnDi1CcB6MOFCe8c93SLnY8LYGsHZyXkijehv2lX3yMCt86weVadiHYEpyn/aECT4kX3y
cwWZncIgO2TENJPRo8EOfDkgs0ZnbKyrSM3aRecMxj1pM8Q4sN9njg6Tfc7HmLr62dK55YizCgJ+
bimWB5Lrfj7jNrBvMIIdwISydjIiOlopG52bDaFKd6s104T2UiytEnGc4KvoZ4CL8a2dnUSCASvE
KX5k34CWExTZKQhYBcYTCA0qsBb5k5501M11eOQZGo2mCKLXmWgo2GogTAhi03XoUMkStm8yOw7l
21QLdnsrzpMX5jc88YNGsjAqo9U2IHip+Yrr555ypOFUnSxBIkpI/tSxRIKF0azcIyvYkqUTrxY8
f37P2xFqJtYPKwBj19MUY2Yp9fFMGVND4vP2GNuZGX1T+MLiI4hJC+c82z+kR8PunD990qbKxXiz
S1SFS7D6MlPG6HpMtkZuqsZEo7kzBvUdaMehSVEgnhTh/oSWXAy24MhctLS8cBHw93HETcwBrxid
BoOqiHViV2CSQfJWtNz5oWqm5Mpk36HPRwoHBL0Qr1oJEF7xkIPtDzmjCRjWL6cUTIw10Wh3rdSx
CQASX4l5JGVX87w3GHLNGx+Y3z5RWVseh/DxXDdVJ0duiouKuVMALNqjSf8hE/E43zLK+909IC64
3+BMmLbQD3C5wtUHru1v+Gd3BdUq3iDR21/B/Z6+qsCqs1Myn/xH0lPTXS7wIXOt4zWJ1x2QxBGS
5RR4bfU3GY7vVBpBl3lb0rop5jShAB0YIDOOFV2Kxo7IIcMUVX/pAGHAopDlxn0f1DeGcyRjxCrY
PMHLfLWz7/ECZsJt84QKffmJoq3MREDbrkuj5c+GC6fu5AgQPzGuQD8WqwbfZcDrTZ119L+SjRjQ
oovW7U+YRfGOOErG4X9ROQ41R76OmTHoUEOeBdXQLjDjrbCFJcweYIcGQw6Pg/tmQwM5W3JgVt/h
2mHefMsJnaVYATcSzw82TrkMw17Iz1jkHuR+MWFdwBDAEWZC1zqqFtKK3tEoHkpDRGEp1iu6R6pR
Mh9T4zHXy74HiooehbEbCByXnHduiP0kEBqLrn2cKG5QViEQEYjXDmAApJgcD3OGb7wvWHi2WzaK
XMgqqISIXG3gB2XoO7D2QHYWpU1jhi5fnGDvPEXTLRrg81AFnrsfyjjUDKDAvQ1mdvcTFq3YHwSh
gRniEqkNMQ1M9tp//okpNjPIq8GMPtA9+fKg+s/wA6iy7d4NWY0NbfMNR6Ew8Oh0R6vn8wykcoY6
tAX4rHvgPFiTzper1GR5nfNWpd45wGu9sFN4axNGqvKmRziY2rGT1UFJSE7zHNmVaXTR+UtruaOm
kWXcEqgWCdbMR4GCUIBMZ0dy+SkLsZx+WlrJOgu/g4m+C28ySkiPBClOD3L6kmNMKzZMER4BN+kw
UFeBJI82IbXyyatfk1PIn+GRjHQfTa1BthhMePVDc084lUvz8bcprGmTQoHz08iPjoN0IgOrBHeU
70e4i9v5YSl2k+aV08gnqaZl2csvCCcFZRZgaFVGKEeWgJoQhUW8Vj8J29zpeR4i3TzritDCyRwJ
I3IlKfJJSP/WruzS4Ld/kTq58KIBUhot6/VX04gG7vldLPenlVdr9dfBzeJmzrz+aaOC+IlAN4mA
q8aCGEqwSggYIMx3LprlMxmXxVwcxjRHPtg9sSUNWqvvyEWnniPNkNBv59vhyPCAoV3bCc83eN7I
sCJwjfbUGSHzu6yU7jTpC96cq5I768faPmq2F/2xLSsYxAoJAQQrnDweUi+Iie0t8Hqz7yxl41oA
r9dMVQJEr/FTl/DjLVen8e9/U/sQQEzVxE3+5zjSSxs0uEZg273DPSAQzszg1ndA2ID+DT/yvI1T
VJBlIKqrEku3yIiick58Kmm4+/J4a7HnV1wvkHX4F693LPCBQRm17MDM8gQk+/xqp79RaIrF3kOZ
xgA50Y0skWDISriPDBFoWvJNY3jhn+IztoKabWfjpG6AZdt9dDk6Z5lmlcc8n9X+YTt7nOLPWMFc
KBrUl0pAihN808fsVC7QEbdH+ZW9z0q8HH/74AvqCrm2DQxS4KSm9g1z+HhX82kRIpVLGxPVtcbP
sNy5WIdf04lwV0wDlbbYXESJ2cn+jcFqQ6wJZp3mKx2zz/NGUcLsKCZ0pk0MP9OElLNtnspunU/H
P7vZRZDSVYi8rFb2JF7SH/Xcqna+kL9f9uEHe83t5yjROczhfR79xy6sj7bpPPYbDW+zYYHJFYKG
3iWRzZldpJ4SRxXaI1fH88hOgFN0t4PawAgn3Pa2cN4k1vnNW//RDOEzEICAH9unMx3ACV0xxaQb
aGmv5mTLlxvUKG7c9+nmnoz2omvGy9+sFOP5+DRRP6v4cRd7jw7JEma8gPpHiqJJnbnqjVvIIQvl
ex2YBR1ILlATDKME89F3vNbhTM3glnS4pM1asRM6QV1tnYD/b+/roUsCnzBQGvysLiZsH0O9iqYm
IcOKP1TDTjWCVtsxvXzzlCnCKSiDBEZfM6ptmMSeEhJSaLxJBNRNX8d1sLxTagE7g1RuQ+VtiiOI
62pFu5z543NFp8g1O9LgCAIuHDy8klwiIf0cHiwIDVCOTQ+7OROmLxaMn/rLfJgKB0q2l4xxEtjr
GpNLhNdNDRHQln4TdELnzjIaoZ2crK7PwZMhOfp6lUVhHtSQODefTWzaydKPLZz3HZbbV0OePxJJ
wtAckXMJ97PyBEK75mU9CQv9V1+9lsHjvgLKcK91BvoDJpG2krHubDH+5Iq95b+jZliolKmxy+1y
vPgxXAUuWZKlxOj+texW+8WXX74DPYTgaG4tPpW0kyFgWmat7BQxphsJvAuDrVnVL7Dh/fJ4I9a4
1TjHw0J9MiiMgwrS+8BOR+Ibkv7vCQubJCEi5LON9pVhlUZ5DNcSCz4dD7PKSI1OVYMnmQWMX9MC
kWNWDswhzAlmS6YMAzYTP+tVG5tlLbx1DLRcVPIWW0DEPHhuYf/IyqO5MAzeyLxmDUtIm4QcCJ3M
eiAX5gOdPk6AXJ4/MHwlfW5HyHB1PvB5b3j6UN6Tk4Rs8Ww7F6RJsOwoZY6sGLiVjUxCTB0xhVBz
8M0eUTKGAApqHZzS0TzHVlvuC1PUG5/3eirCrYpmdUWAyNpQVp714o2x3hz80TYUzyooP/zDjt0U
YmpcYX0FdNACv75s2x4xhoWLjST5IPOWMC3w5stIiH0E5V4v57pjsOsaN6KA12qsW27gqRqqmnSj
DmL0WB3XR9fc12XW010nNPUHtiNHQqbayFtgjlOKqilT3erQLxCaRyR+ObvO17an3OaL89rLeZzL
a+SF6kM4MfiRCBdsez+ciy8lAEIKpXwLk8UzdMVnVICSOaZlb9hWaMskjxj/giA/PfQy0VyFhXeJ
u6653P6tGsaMZJAyzbVDVej6AWVATpvg1u+SF2Cfg6Ia4wdooSutk1WJVYsIXf8Jenc/BTyDotNw
oWAOxlwA60Pb4y6pwhF9LUe2+/ckHUHL4FqYs7z45ywoHrG6kdx1c1j/i26vLAeAWvc7YXAkKJ4T
MalxZjXSwHMcVsxfq89tp1YJ52OZre3T1bQB7CmOm67S45277sEONck5TzRCPdXthw7sw5Rym26k
P5iSbgRi0chpQfD1EohZMyiqGeXDG01zZ0BDfGlzAGaiVPvP5+2RdLli6DxuKi0YBxnCvfVl6snQ
jVACouGzPYTyyZ6WoTDcj3ut8X0WqaRxvY7FRWjMHt0lKnAAuUY6sJ39HbQtzDojkKfsRixj7AK8
zPaWc/omzcTXwNQ7iQddKRFF9FPqhYsYAtqKM/K7jfZsmWJWWoSHfyhO7inhyERzF4AmG4k9Br9c
MXtvI6yoXemtNJrzn+0yVtiuastYpk2CxWXKj8R5dTnj40MczwfJinS48hh3M8OQxzWdxGRTjFmD
CAPg1yhwVJUeb/77Kl4ooOZuEeCzjQzYVH2nQTWgOTEsP3MDdTvW2ulGpCEPSs7+GR6Tiw5sniGG
NuDwv6sx3TklS1TuQHd1grmUDcAIBjOcZcTfjD/wXTCkIBRrDLgWME0auvd5l/q2xqq2dGS3yeTH
exEPJAe0CjtzK/VYwK7OpeH2iNVwmoy8ZJI9rrJb9MPWu0mUSG3d4T4e+bhxiDV/+ZWAN6Zse7Wp
Cz9/o71EV23D8GEweOfPblOghRIufZXz+rECmGaK5A6zlzI1iedk6BMJ5Dg87dYvjl98ds0WqgiR
gkp5BpB8JcOPt1XmJ2ndV6ABqJtzCHlgbDkTts8qdBluWhjFm2sIsNnoNJLXvRRNnB9flD3QBgdU
BTLQ1tJxJ3OzMhLKPdOn7udTBcGTkvCVAyPvm2KRZf3ufTVuauBTvANbRYhQurEuxp9cRykeD9g5
+i/1gWK001LbTYoHiDkTkb36+anobZrgX/hCxtG2qfR6H6XmD1u28C3IZOb/aJ/o8gXZPdo2GnNF
Wtf13ZQpYg7bGCBM6agaD0rEvtVJ2B6WSXS5ECa1FJlkEiD2ZHQSF35p6DJP8EuioR+hNj6xr/FH
pwitk+3gLwfUBzEDg38di393MpmQvMW4H9lGFQ1YodNi5hJXM855wurkm7DvXXjacI5E+RwTQAxd
I92OQv7oC/3qhlTrqWf6WFCvNaVQLo1Aw4OqragFUyhkmAR2WnBhBbV05k9Jfwyj2Dllq5tkU0pm
qYpBvHAll/T4W9Yg8fSqcnZTUyZTeR7iDKtpY1fs1f91/PPGwEFxx71p7Bxdi6uJQtm7o94Pwa8n
FSSRDpKdhcx3gVOD2rmIzDYnc6LohFNhN5sEmcKqcJqMApJu12a69azyXM7JqEX9pJ4EF1hGiPRU
TJEY1nYZWolUkZHk1lqzR5TGagTr0rhPgjp1u1TOLC9tgypj+UrJPvAYjycFSFrF4aCXlHLk5Npf
QxtN22GHQVFARVQmGvTaRy7YRMC8haVg2IKRprKZ7PC+FannPDR8i9BatH0n338JoqndHhxNjJim
rN1zyqjsDiGPfhfnMWu999A2mFzuYYpwgxoEOzMOxSk3jIFe6LyyyrwdSgvN05iPUXKx8JZEi7/I
v2UC3Ehq4ddSFaEF1+xWbQ/nW/hDXUxZdQdXpzby2ReJPnUGJvO29M78goHlj+kxWpNMkzmVyUaa
yZTB4Wb1rja593w/CTVC9oKxSkKMY9zxd/CyDskwfPY0ki06YYLZX3xIM5qlSWYrlexJAjVLG7P6
tksOj9LbvJprAZjkdVDy691XfQFcydHRcLPdVHj+BlM/Y/84U8QU30AjJR+GZxMAklAA7ips6YId
vy54DyH9hy3bgml+dIhgVNEm7e3BXzMztBpAY9rSKicziSS8Xg6dHRRFW7ZvKLPofk4ot3gmd4ZF
ht+9O/YYHOmgWTseG+pEkolh+g1z63biyVakj0yVtEFvJewfEoz5o3Bo86WLHeAGb1Y7rnoiH2B9
aOupbqrIarBuf7Q8qVH2hZOzYdJjCLHqeSNZ28R6/MAMrtSBrpRVMKhvTtUoLDFqpqRb2vgioBEo
W12K0g6Q4Gbbx8URfFR1ngEQ8wtu/GBSYRQJvRt8kwwABJZbpo0Ut7DGwE9LuRcp2slCfXogfVqO
ok5xxdiZaYDCw3kRW1dRKwcKbm2964orKAeG2dpCYLi3dh4frhUYFAR/cfKJZBIIR0C977/DWPdC
m06WddxwLC1Nfm1kLXGYk+/iWynVQDrJjV4wvYyTYE1fEpCFzv5EivtloM0Om+h4m7a2e+yClHgN
DH7V6dWDI2DUg6ZCe+hBqZjcHrMnufuCTwuDG6o6LixUpnmeAhZrcm3/CInxCb6pxrB2JD4/l2Nv
JAEnuY4qVAg4NF+5hZUGLlrQn42lIVMceyAaXxjwK/sJm5Uk5KaNiL62DNfGA5kZPbqmYJzyRy0G
ZxiGmFBnIBRdM0pLZmoXve5cJVd7bwPp96icSPRv7PEl33LmOcilxiIcDxkji/MSUoryHCzR7jWy
hrULp/DhtNkSewv0dYfGR+olkYWRm7t5b0Oo8jwQs4dOD9taICYMPcMuWoO45OUP01gQ4K2uJIEN
1q7n4uysNtCc4loMsHwMLb/KLQlG82aTdKv35dQz6BCxLb0wId/WRMN59DWXIMewgW+OOuMczn/0
rxz/+Tw5obUwkJVL/H2ayU4ry83Rv9DFCcRxoEvIsRvvP7NVBKMAepBFe0LfYPqVHDvLS+XvC5Pu
UP3Guhe80jV22Ko8WO9AWoeRTw+50OripviTWoQu6wAXf0415KQdCAyj4Hv+h/AJyd4qGVeEqj0s
PQibH7ftDWc+JiJrvnbf+QUZt+wzBriYKc3Kx/mljB/ICAKNl/3/p5W22klLlhUb54VA3ooqENC7
veIv2aKw8NR5f9G65d4PZCVwfKofZxROoeDLVwJaUwzvSfGkB4Ll/mOo47aLwDnAXhxeYPUj8uqz
0hFbL+7WwFBFqTzZKKcSLNdtFuz0abTFFOYWeybcBYzOGVg02K2TJc8+qHoO0mzF8fk3L5YesP+g
ocYcysihn+l+N0UIVIGlrkrFJ9tPQr6Qaef59l81usJV/uFpyYXhiAcp6VBYF71NZD9co3crLbah
A1Zx0WhbcwPatCLV+sF/6rbNTVTS2HtyZujISHvEgZy8s/QL1wWjUoFytLMpeww7+o9s4JTMp2rk
tFjgf60wXWaf1y4jBI3dT/jgGfGwAnBU/3X4Uk4pmf8ljePafa+s1ZgcKbxdyZ1sud5hDys2leNU
nI1/7r2PGX53GRAPC3uUCuBM7MUAGESJ4ctXm2dcX0Qy9PiVfbWmAoZJSdy4xt7gNrsSX3PYJIJu
hvRjPk7vSxOzjm8Uly4Sg3JEqLhDFMT74OfxYXGntcyZUaK08WJScJ6StR5uS9v1TLVbUnn/JjqR
7gF8LdeJhqrMafsNqQxC7ay3u8uFDdyhHUfwahc91LHuYqS8JCYPJaDBWK+n+s1Wowzwj05P/52i
CjQPPiuSngmtNWR5JdpqjaQ/kw/DS+er9w4fCwcuurf01FZpVtSEePpuX4dIdfIdxXDKk2PmL+mO
w/t3B1tJ8u9mqxVpDQSVth+hpAbpOW82lIvk/H4nVBHHbmJd31qWbYISUCcRwMDeSMcMGZG7NlHT
rlNCsP9VMqb9Xx2LMoQq7R0Nb4fVe/4BPMcOA09Y3GOzWjGmCyhmfI7KVB1SPrAvSTnqWboQqmwS
gZcqCpbPYrnzpS0ImU8EAsqL1mz7Zra4lPJfRtF1+yJTJ/5ygSq2BitZxIq1QLtSgCIj2EZBAnyP
5P8xqE2QYFZ02cjvZVYNy0fHKOBM/MXFwnFoMnA8SWE0u/42UdzmENJsbyibpkAqscmYV5wTh0XU
EoKGQBhyNl93cw78YF0SG9IHe6muOLZTfZ6nKfPfRjWn3gKqMstQaIvG847BObo/Zw7xn8Pp+wBR
ufnEHIEq1ce1UPCyc3WiLQeIZq087gZ2l5yXxOgM7e+iz25PLOVrYz2pyEUNgvMidWs08tThu/e5
8MGdAmOkdR6Nac6cwjQcQ/h1STJM+vTHqO+6nOfrdVScxiZ+9/mwpi8ltl83SEBjDRTtoGvGl/eM
rdqG+5KxCo3c8cJ0mQpUQ/dhAQqnvtwq6lfxklguMw+RMsHD/MAnQaRoZjPt6FJLXRYM0jXPx8PL
KyVkkjPaXKSUu613eENm1F3E7cFlKpcEQ6u07voX9LBMnfKqZKxrOb4Pc2EkDQ9BtBNC2X3z1qvu
CJSrNDjDMD0pzNaK1a4f6rj6PNL/62yrQiOaMHglmaeQl/KdTRpzaoJJa38CQN34RKJDuo+n7Khr
S0KQmZsJxGeBoig8qLdlUySSopn/+MoCp4dcz/wZQBlBrHJ9mkRH0sYQ5vSxBsd9S2+HFYCES9k7
ZZYHomGHrQgcDq2Tw13fY5SxldXsbPQv/vo6D55sfAuH7pDrYk50Yqv8FpPk8X+k2v78uW2Y70Fw
hgcK5AUzv+DkvHXAtaRTO5IEj3nrn2GZfxChkzVEMfTROOTbpqu8tUR2uL2ygWy9kBW1tyrustDw
6AFTjoZ8Xj1YhxXcBHw5GF5j2/Q4u5MizU9ERFUbYfgIswzdK5sxTmPuuFnLeM5KhyOm0Ttmp8pf
WcOvZjTLaHj1BZFyC0K/Ls19oiCRfzZepH9yWVRzbw7LkoZYhlSJd06uBBYn2kN0zndUVoWOne91
U2UIz6HVDj9iP1deUryreT3srrb+hqL25q7M02ZAl7YfhXH7P4yCJgwaQoZTGfkewwxrR8plFwYy
EiAqHQLgF5vmYV+3dMUbQyTbQYygg9a2wkqq8f9XZA2tqYXtziS4y5Meot1lCVRDjQCWtnrjDg88
ErIiKox09LyASiwVl3eAcNSfC/UbgNT+qBexzkKmmmmeeMjprQNsfuCvlHCWyFXm1krm3sNMmBqP
TE7bDm3rTxgkp8eukL0xRZb7aMfi21x9SbU/RCvvYs2mDZMzQhNRtAZ1D0ZMPEEDVfl0Cm/h9ISt
TvrSO9Vt8/BpOss53WXqcREx3TjmCRTj+jnnxSNm9IPba7efZLT/xY53kFFmOxoFg7jVce48NVmx
VkzCsHXNbqr0BO7Lc1AZ4wYE4esvXM/T/SO0MKzOTW979GDSh874M+n0y+QzcALAajp0C+PbPO7t
iLYc7+Luj/mCcLlR4T94N/gKwMQ3xI5wdvA12N/a6JWp7DaZfUJE//KaJn88/46/cgg0dIbcrq5+
MVc/O/0k/p3ubVB+3QMjKM3zGJd3qxlP3XCKN4mHMIZucySmyRmkcoPvV6WBDk/awWnRnGgZeEV2
WdwlO82u7JIo5RqZCwZ4T8caAvPuM+bmiz0HGH1rELvrgtgpouJZvKIB0ypNV7ilhFq3/+uyCKdV
PuHG3jhPa5+CR7HiiCdrypKK+wmczPtlX+htTmalvoTQ78U3sk5mYmW1OD4w4yDPQVlgti5/nthz
Ng+7oeOKfjs2lcqYVDuCoMLp07zqpcBHoLvETp2kJyiGyNbgrhh4sxUtYE2Rac9atNeWA6xMDlWg
Wm/jjlLjkBKIds82QM2oq9VVhOeO4PjoY0i4MHK6ZXQL08Ia7G+iwymUCiLKucYstyAGOr50vYFz
SKh7Ub+yTKAidsR+ve1frxPmIJgDRXxDibpaaeU1WBLuTrZwQCL14888oTtH1EXz0/efAM3wlngT
X9GGcYx/pqxHxJ9f4oLqLbr6AEjsSAzhBMRm8FsEys7q9Y8PE7bhhRr3lTPbl7LtWA/Z57Tx+NIi
U2N8FUFJlDv+LFK518QwcLrJ7WN6BYqjzp/2Y9B/16B5DG2UEgH55Nu8RwG+j5XXYLSnbxXGQRv/
k4xN0anmlosPhgNN9ySn46Z+T19X4Tru/k7hzKf+QmESSh+yzgpIXRR+zoVKUEVR3amQjBteou0B
6gqulOoOq445/eO8IU4U3RsBzwMkoJzKfEFBJAY3QYpQPnCh5T3ff52m8/Eh647LK+E2E7KpROwj
yJWVnzX5q+Bz1AILMt1EGAlqltylJp2zzfE5Ho5DndT7aUmLtlhflk9KkLohd61QpwI9WwvUjUnq
9UhuGB7Sz1T0LvKdYU9GtQpQSd9AUpJoCGLC9fCl1/jyqfR3Utq7rWN8PcSo8cQfyzaAMKujgDU7
ODwfxHq6Kf3KrVQgt/1JK5agy0SDD0OaE1wTaRNiWi0yH7RsLjSzX88T68jbwas5IZM5L88p+jU1
rZlTwqx0byNR7I3eIIQbTeZBLDDYpSP9OHho3ruda+8drjpqpyt2ay/UYZW+m4E17nYqXYUxDx0O
pWRWOa3ETjlt75FL7/6KWlY+ARSpu1UBTvnNNJve8MRU7inw4H3sNhJNjypW3j6n/L9tdOqAx7Pg
phEAazNKDoqAR2ES1PY3TP/MXGgmrMipwnFtRODYIf/0TYeUfGpKUpcmLE7/uwUcaZq96vk/iOfo
abITnCLFdljKwyIHVpHmDUs369y/1fafkWiA++bVBilRbF72h+SPwb334EfTOCP6By4qO/rnyfuE
vwiMdsru2zQFarvS0Sen+QK/5potvW4DBooR3JvnolukABYyC0zFCuJckOALCe1s1ODab58bb1hW
YFh+UoKP6XMyIh0UGySAarKos6StKISbh9DuVGyXLKCqeNfat7WJZeyaZZxKjTVhlRoFLydSZ0QP
0JPKwnURSG/tZ+vKJCXoGdRWHMbDDtsxmksdnfZyTM35KQvAXiGB6/Zf7HMjyC/yyfgyO9aPpjPA
G+k+t/T0Z45R1vXiR6G557lmCvKttH4Sk1kX8C/EPW8MAX311EfSIVYuZuzTEb+KcOj9ra7kHpVk
kf3eustqSvrXc4F1ICSpmxczTBLRz4MJimi8VNFraU4cHsH3ixXakUD17NBXX0xAPeDScLZl0iAe
Uo8Dw7vsfQhRUcNEUpXMBJGNXl/BfJ0qz525DAHdvo6kwGqdrCnrjDF154FG5KfsBxOiAg1r9swx
redFj39oFHZtYnb418IK09g94cCC2AYu3tYIyg9uWLzWR7Z7p6R935aTufwyQOiAuGSy8Mo3diqo
YPAp7frYwY/efznKsOgaJppWHE8WARgH2mSXy+k+FdZWl9S8/Rqco8+K0PV83LvGHtX+/byAD5bV
wPRnE6A5qV72xX8BRRRQBFoKhpzb/rtJ6RdFiO8/ZXNPRrPPOp8tbMuJPYibUM8kWJPjwqVnY0GI
mtV5MHDzBXWnJwULGGjSQl+bTL9PP8fxewoEQxAQm9HPIyZUrQHufhB2nESYJ1DV1i1a9Svda5d7
Ux/RXN0UIT+wj+vq22Joinxk1f6S60SMg1YWR6RPnjrJX66K4JfLWLvCCKMrRyOX3dies8VMzADt
UlnTMLY49/b5ZqZJ6YU3K1sEKIOury9BJ+ua4GWM8LsHRc2R2coS6ulhLmbgtLJDYLJpZiumD7vt
Pi/ixgGz6i7CxJAVLRLuyyPpjPEGWL5H725/TN9iNkgx8XjKDAMj/udS4CrIedfKAf2fzp6FF0y8
TseIA1f+rdwIv4gAAMUrZ6WoWGJ+30oTUAtF0teW5sJA3wwn4GCRd+BPMlxDW8VcrHZvM028PClb
UxU2PvpafpaJzjkpLdTjrvS1Kh9UVgzx/Hyh5JYO/daHmdDYa7RK01JobGBkx2NiGledHSjCkQyV
HjGYNCTh/0KChBW31c8kVP6E0XjGkDDtgp93ljVaa69BVvMOgRnB+fmfKXHpvWtpD/6Mhr20Wfvu
VxUwiVlYHFlEsdnDbhM1ox1VYRNmdg39NG6t7t74q+7sOhNxiEjTWdvAkwClAnlOT+ei+ZbOun46
jEnTLEDcZOvtzqgX7/IOwKSV5ZmoD2sybXHmgMcXEV6rZELIoLV67BgZlmytt/wDFN0LK865hZaz
2TGyb9rsjC2QmFlJqzq+lpcXQXSulylaV+zRzGh09ad6phiERjg/9usqz/1temn1QgdUD9OUicm1
py02RnB28QKTdsRLF7U9wNaAvavzz5Gf5ofAmArrFkmEhRF+bevn98OOcsxhcLRn5q8kV2F2AYPH
xfLKUeqL60yumv7B1vgFkyLZHXUwsyCZRsK2Ln4Pdc4ou3BQnEIQXAGh5VgTHm5RJhprzmnjEqh4
PFVg+CblQVo3HrcNumhA2cyR4/R1zrkgeLYaqmC8Z8nU3WFtm/dQ7GuLfiomn51HansHkHBYAA5j
PX3R5fLsoQtxCoGKmrFpOCubjI6+396jQtqWJkkpr7IeX0eJJH522Trk0a0qYH1z2v2FjWL1n/he
pUewHl8kt4u/3Z7/1brJkT38QRqAXDsREHSHgEFQWfgCX02P+QGCiSzFmhHdxOA70xj0fXMbQuOP
7lxCh0smobTle3J/Cp7obARMRSsiTKQnupxFEu8ai2iqVzwyV/djs9fD+zmOXq1G0tEkwrmsV9s6
sFkSRgaFE7JcusEx0eFTODAlpgEh/gF2xNv/fX8OqgYRTq9xJfMSyQVtH6jiTJo6t60XIphY2HSr
dw4RVEVMT6GtIWBFrbN14C3kGYIZFEqjH3u/8Vr0wwCuJgM99w7VLfTO3YdNP/k9gzNJ2sHaC78+
3C1sRM20VBktJQyt9S24kPreyOEywz4wV9dhH2r+bwio3MZUmTi+JazvRxXc/EsfqWO2tXJ6Nbt3
pRG3RnYI0kPXYnmMB1quxh9tFIw2uNTpjRE2Cs6Nj73rNlh0W5MznIEvwC81iGHVcEkb3HJ6PM7B
f7guCcWKkBZLhmklkMLsQ7Igv+tKLcXD+L4o4hGCN6S5B39y9kuwiDvSX5QbWueSlPyqML4eA0zp
epL+CH57GGTPX2gZcK5/Hy4vcUhlqhq5U7imFBYRW/Ef1SAOfNQ58KCNrfI/ce/gpScy6qH5b23Y
wJNgI1IbM2Y0Lb+GL5KMeo9y24NxbunOKFfrTYEBb50WPm+p19rxy0YExaZqcrqA+DXOY95tp3mq
Dob79SOP/JBDUAL81oh9WbzUkUDLRdLpU0s/aUd78K2VHZLdwI0UMKGrBCWjYBej6mSkWONR0uLF
ls56wZjI5c5VExuYU/WP4l7fPFVaooxkJb+4+/dZaVUFDQtXsTmplQ5zSk9jBTOG8NogthsNfIgL
LFDf0+b2Tpa40pbAd6hxI94fNBBn1mJy7kb3OaVYPVLAruaajp2y2pwJi6uu+/RNYq2uWpzSwvTO
KuGEU5Dzjlh3DxyHikeDB9xpsAGE7CJzOXZWfbreIRWMS6xCyYEBMMyXWIG3bODc0ftmOLa+8W/a
SucleuAVjKwii3+RZV4I2cJnM6JyEpaIcXR9SkxgHXLssq+70M/e0v17+/s+TzelsgS+xEV2bJ5j
HzKHOPxvibQ6MWR4Q+PO63Dn3f0/6FV6jBZYHUOGZMJN9gakCmPrbWIOwI/k8kqsq1girCiXkb7o
8A39/4L/jGSlzV+m4Dag3D5ajy12LllYTPAO2LMgDA91FJYXLV/kKYi8kKLPTy3IyiDqA0f2ErNw
Ve/trPCd86hyoj7hmjsQTnrEnZEup/7jSdj7SpukkYVUzmctycSfHyg+acWpe/U8/bJ1Ndh0lxrM
Z/f484aRirm5hEzFGAfj6QDGO+48xmd9Q4fAeb5cLULwSzpLPcif97lt9qX7tWmSJ36ySs5PIYmR
w7Twpyg7+hke6KTmjvOA1KKxMt6ybG4V+9AJdu38VlS6QEQs0usO7fkx+fxzh5QQioJIMu2O+QsK
dyJ8nCJF7xcMA64GhLO/PqNB9kEu2g2qcMFm94Qp+RaAf5bwiZVha+FRY7FztpHxWXIehp6ax3iE
3C7Yb9zk3QqNm+bmPmsifG32/jTbC/StMHYL1bWa3y56ol2mDq8Uyffd2mFeWxfXZtmUB2fpu5Sk
s6S508qd7+YxdnIS3GaGdUQFTkRhmrSSPKDQaR6oBWIHozmj+IUtEG0tncaOiX3W0bAi0DKjtXzK
rb6nXf6LGBtxjOPq7lqK+MOk5a4M7/BDM0ra5faBAAf6UpDJ8mFQ4qVW5pFdFGIEMeNKcsbPTNKe
LDf8msFZgUKcaDnB/2lVbyoK0H9kGg/CV8s8F2RJN7jrCYr4m2gWKHFeo/FNwCdAqozKcxNecquZ
niDqC+WfEhFjOugKP5nVxkzzuRT/+6IwDqqPOJ34A1FMRhRFs1CwcCXdNH/RacIqbuoQnzlbyttR
pRmCXxq8++X1+7IKnuRd2sugNSgqs2W1mnP+jV4dH8LgXoqVEUi4bzZg5kNoWJrEsVFL6gCHR7AR
coNezPSUJ1g8nNaEG7F+RUkpNBk7icZ4SEA6zvNF67UMH8PdgRNEq1f7zM27rQCAfpCMxelJvhv0
4ezzUCpBN6r/ff7Fg1UPLo6i0c0/9KsHrbfExfikmSeENY+TMf/8yJehoFLxIeiDdqJqOSf982F8
I5lZjfRa482AQOTs70OHEfc4XnWPmlLf6ZGPVqoM5A73pt24+e3t1pHhpsRyxiRT8AbWuLsYmtVg
SIcsDMzWmdzsV2zLsLoI1F18h2mrPWP2DRfJkOomPwnljlkzcmdpyBMvtS+kHPYT7x9DJtVy+79d
mn8+bhldTlHlclP3qXMCm/KBgLqUjHbJdQnEVorBPSY3D760ugBXrEGRv3dc1dF1gGbItMxiTOG2
/YGdzaUkSairVDwyv7MajPWm/rbA9qILZxUQtvPP33eN1F+Huo+170D4Sv0Cb7D9avfk18031UOw
rZPSGIQfb7dZBijeMA5MBzbb1cVrlStkmRsDi7P+RTC80NKB6vgaG0oU2kJap8ikTZESsOyChARG
TxbU5fhII7a955KoxZ1qtUFu0WfFdAov4s03TFHxA8xu1rvg5ROno3zNRodM/NOP6HY0IXiYd1LP
0ekhJP3v+voKLjPqF/3BIXjsdHD1VmdRfGXnDTS+gobgiAARY7e8sHqDHa2NqBxwTr3Dz1diDS4h
yeWIjnDaWpxFTbGK65XUAyHGpaGjVKnw6LKUsL07w4dZqOu64J19Cd24Kb5tI6MlDBAgGzD/wEby
UETl9L+ndwbyBFASWq4TQLJN3plntGWb2LHXk2+QS99XonIUlpH6FL+2cUeaZxI8nQ0az49AT31w
6H4I3GxptYipSoj//cLxUtEKllI1dm3pLJJUjJTJtKKoQunJkLHOCfFM2p0/yXgWZaeQ71kKpXOc
dz43o5gR6ulsKk5BWkqyPQlWHeY8oNdz5p2q/z7GD74Zl3LCbAvzwUJVuBfhbbaM6crmuq/DL101
w0oEGTHbIFIG2ktwaneJ2IRi3J39S1iHMoF4hxlKdcyPDox7Jr7BIq9wEdy+LHlbRseyL9cN6qRm
ftch5I/dKUkftMWN0fxoCNcg4ZCoxkTh/cwMQWD8Yxb9SCQ8+PuyVkOvPL2C3GwzxSY6u+GQDudK
s57cfEEuuPnu/NT8pFI7EI3f2atI8nojp2I5dGHfmZV4ZKjhvoyLWLo91UO54IkylS6udu0URRdG
j8OZy8Kl/0DityKQo8rTvCNsQTlSpm2+VUhgd4hOqP9rLFQFVhFyhjXWQWb734qETMqaxEJPMNN5
N00xN1d038qfFz0k9UJfRGNIH/mBoYe1mVEt/4/AOxWwePLgIYND/rMDL/mLxKt4/bQnNmtr8HGI
zNiUaelLC/zqr8CqgI2x8TLACIbGqxjYO1a8519CjE7nkmohVTKrZv12yIy94H1tia/xdV4WPPsx
NFa1zRFQqixh1y49XPOeXsIJl7S4PZ600P4w417D7k4NlaoRDhq/+8/snGXFm3hDSYjI7ozwmJcW
ujkGlbVyCHLKzyPhLreOta8HXHV5BBEjz2UvH5TLPyMVNYWbuDWY0awApQPWJtnQ3FaA3U9jmjiW
JlYJ87Svfs6ZmreMy0dpeVeB33OTrjwcP+azhg6oxs1J3zY7xycmJXR/2iUcRH1UDpbhHaFyYaoD
sdrZ5de28WhGDMxp1oyTbMfdMGmXDc5j3lFkO1aba5qOm1Z4sdDMJ+Hdw1LIxDO6mnk0wqTmMnRf
VaEbQR6ZB1eWg59ODC7pi3V3WOlIarf+zvfSZguS1IYHemqhkRFLXscGb6mR34CO41oBjunnrXcS
HQNAupIJZhBZA/49CjQEGDoz4PD9tRDk+68J8blhIbfJhvvfLbTeR+z+QjouLDQd45dVyHAiKHcG
48wClFZNhVmN10DYIXRR/+PvQ7WSH1OIL0lRyns7zfI7Rn+Ff8LqvxaT4cU6w4X+OvFhdcUwKOaU
4B2LCU5+q028p7AalsuhGtmhA/hAUnjwgR/64E/IKqwVcq70RLDMCGrXDIrvoWjMOinQN2+YMgaK
fIBASjWJ7ilyWbrjcsMOk2ihZ1bnPS5SJusEOGh2/3vvKI98AdsCfcrXivbsM7JgUVMHEFx2Rh5K
kIaPjbs+pkQUIAHvOv29B+qGfjtFaYRQ5jsXmqxu5tlB/F4C+Yn88FeYygExSOnYqn651YCz8pVm
oCadxwk9g0/LdViF9scihRA9i+9o25o6wz0EWsALj8GgZ7amUulUAzbDUwCbm7YfDR2TftiCMoPr
jCuCHvJ8y0uHGlw5+XGKEJSG9cjon26UMo5dymHhhqGhoDLhCHGFwFEQxNrQAO1NxGmQFZwfAWDR
9Etc3mfbs7yGn1ffWPKqRD82mcCRYzG19XXmcShWFDcE4UKb/N2RftjBnyNwHE5TbJJjSokpH9Eq
uARdp39ZLM0c3tSmYMvCALII1fX25Dnx1bGj282lQLMNpdLUXB6n8tevrJun5yVeJlpZWfvGuS+F
bKZwbYhw2uEHYuin4ix892R1rMQcAkur7fldUyScb2Ul/wHN39N6CnmmQmGPRtJCtPTLCdMfCXKR
gB3q15/L5Otzski1X62JJu/wZa9n9vQYOwXZrHcGG05uy31o2OOuBDmOsZ7m7hyVvNo9OfF0dgDQ
tBTrS+rnbEwY6qVn1hhk778v3GrntZbS31O4fz1oZfKrk8eaqNc9MxE931v6KuzWBAGnao6onaxs
QEOJzi5j5eAd5tGf3ymblV+9rGzsMbrV9csFJG1m6i6DZNrX8Rq4XEiL2QGaDhP0t/JD83j027F2
5iIdMekZldUlZ/w8PZ43bvh3xszb8/FUhl1lCDOCecdeB8+B8s679aUo1MBN5CCOmp+vn+2odtcE
fosoty+cNS0v1fYOhKvOZ5uugtVHAmJupuAhQd0WkBkrCjeqPqOiqnqIcVqd7RVw5nXvj4CM5Trb
QWvJzRYtcZSfrPsdrTtJoeqIK0imBmtvlSpw7Tal3RBBhvW/0xjrwsA7SWz+xk6umsVdjKtJvZuB
fRcFAF8CdpTnzY9f3Worxv7CCvJkN4gENCtHPQ0vX6w15ElpVQw+ok90z/LOte3EzM8o4ZQShBVB
ogvwlEQd6aR48N5yV8INLETx1fOqYRgi7srMm9TZgbuICAA7/9ApAuDtgAJLFdyQFxHmqVmG2GOI
NJ0KtRqLZxMbsNyTUpOUHzJDt1aAA1O2Dr+/rFpkuqcd5CkZ8PfXpDPvdMWybIWqW8EJU7BhZcJ2
u4rWnLNC5Ix4ibscqou/jhTliHUrhKR5oomjr5IxK/1Jziu+ZQiZNQne2xxyQPJMvrQsRt1u6l8n
6SpGabfo1hdAE5bQUOylQ0liOEAZZzH6KxxuqtFG6qAfmzZ8cmwxT2CO+HYoc7cTX0PoFFKLTejY
zX3HjJ/sCwUHLkaDgN9xo6FEt32G5fHDP24h+bwAvIT11lSwoLu/eiK8ZSB8OXMPyHgCn2uYrTDb
8hlpQtdOnTYTDgebxUK8WBugZiX9syRJyb9pdGIHuGLLtNZ0tSdMFoL7FfqoS9zb7pCWJw5WQ5Vb
UjL7EvlQqipVVd+KLrhAjG+Pl63z5mKJqiHWf/kDJzqNC6+7MCQgHnL+ZzvALIyWHc3o42a+r7YC
Lpk49UmGoLx+zmuhRIrsekSJrBzHGd7zS1u4pS961LnHbA/CykvGPHzSfs0z+KsCr5kvPPvVvuCs
VWXYHpGPuu81FVosreyxDjcxO3cUN6kRuGYapMQs6PjGSg9abH3ZVI++M4s8dix7XuOj2kck9JXt
oJxhmm4fRbdVj9rqgCN5edyRdEQaXb4+eLKlaZxiLSLT5lvFsGnSZFjDsgmlU4dodVgW2sH8Jh70
gVJGt7k9vxBUp4Ylbkuf+nzjWLLRGs7jNmjikeQbq+efUc+ZX67bh6+LkQns0k28YMDUDUe6tEIl
ZtPWL/pJPZ31MbQRxXpiBtiZ2rj0UqFaMb4eLS6AbthztjDF0j4b+lrsHhMdehw35HN19SJLn6EQ
ZHZy3DFqO/S18gmodBTx6UHzQTZTlRxrkYVYRb01cSATbkNEBHueQg+4BDx7Vk+9yqV4BQsADOGQ
OXMeP55iQ+fmXwDv+sGjapZe59VbDAXti2Z6ovtqjL0zDXFcE+mtzCLwDyUgX6HdwUNXd8FIansZ
pa32MKH9JOdpwNfCv5EX5fvmxXVMIZLVjzZl6WUAR6XGhudDFWzuXw1BMKd4g6MByl/AKV/L92Q/
mdQwJdLIWLcYQBDHq+K6bkIboXIRwtKRYDt4C73ItVR6rwD87gTzIaCcQTdHZD+UE8V/mo2RMiG1
g1NtcH/7jImkGV1vO0w19nhwHpl2Te/Mc5yXF4hU7TlX4qmHPJj5u3SvD7tTmUag6e4BY0f9iz2A
HCkYy8Uni+8J4rQKoJwyb0mUd44clg3934RE7AnDqU7B39UOTqQhA5Von+cMS4kVBgfZWLe0jxCn
qFBPbS2m+1t+mJt/2j+MtePH8i/EVEfxz4SNZfFT/wYGIENrw419nbRcaAmFClo0DbBIvoceguJx
jaFN7oX38Lnyva/boSkZM749LZZyrrz38T3zsygAUKbcowqsG51NhCVy5rxsn9xaXDKxDT7qqiyp
q7WiwWwAnqSyMTJt06/y0kLFzc4tsYz5f8oUCg1sg3SIp1MFdMsxh8J7BL03BgduGUrqSZHsaN7F
UaM5AcL722cnIY3EaU08nUTYOfK/V52nm3XX239nM7fcS4UGNeFo50sX7u7u77o+e/waIAQgOL+d
tvytVaCGnhu72fMNztWNv3errUIsuTIIg5tlb41keZDP+7cpKsP81nbN/6QkZZRc4CXn5TEdwTQd
eRjcsAUNMHuw76rewgOwsbXIgHgABHBVnwzv3HJrFQiiCJLgp2imv1GGtakkgY6y/oCMtwMWUvzX
/Vk51wQpBSy7kf++9EiX+Ur9q5VXd7sQxxwG+IRh1DaFep9RXUjlZ15E2hlSM8R/BhiQKhQHjO59
miiuB3eUzOxHh74iqaG7K2Av8J298LAeWb4KDY2x1N/QgWxrn9h34Xp5a8jCHBlHpmr/nM1YeaBh
UeifGpf+uGPtPr9J8d78ElO8fAgGQ2D7R8/B3qVIQFc3vY5wO4J9+r/J3mwx4rfM14sxc3G3TTm0
mxbSxX4n+ZuhOSs+Jjo8UVTbs4HN2VQDkVlLv6LJOo4IqWsW2TYRdXSoWRYlLkx4nFHHn17zM7ex
38wxJSEzz529yjDRe8NWuIhmpSSEPtsZiD5O/9u31y4dBI3RRuyrZDLVCJdLmGUGk4BT0qcluVxg
1MrHT70hOJH9pRFxUyy+rnlC5+I8/VbFjn+r20IDPMvypXzQZb/1DW86DWcscsmRc4f9HiQ3L4vm
2NxBrP8f7BciF38j3+G82bwY1j42UeohTVmaH58G9pAy/hNgAivPPuxtaPEKQrD1SqsB5tkgLSOe
kRFRVBTY4N3ELrgxjUlW5rj/ap8Q2/TD51aYoMpHZ64GPEdU+m3I3zUUs0Ezh6cNeXMWkFbDYeuW
IFXvBJq+3J+W4fkGpfMIos2wh3/iI8Uc/1yASCLZNHjEZL7U9PmZmwy4i+NnXWfwvdf5u6ObZd60
YlpCALW8YKAXlfH/H1OS5BmbVOmsFRiM3tOQklIXSF2k/1DMhfN96v0fcFdoXCJvOjWbJgMVjS9/
5II+dsT7zZ5a6UQsK8l7ODyQ8CPGSYMRkKfrM3CIo4kcFHESYUS3WPKahzOGhZ+YNNOna19LFx5n
iGoz6R+34Y+hyvbJa7fiGYiFrrj+X55eZXlZWMNE3JbFyiBhjZWtfvETduPlb5z2Y2EUAgKIgGay
tI6hEeJATHBkeYvMi91KVgpdXoU0QXLN/qj0Y7+1ZHMDKkQsSGjN9eQ8RhOmQ7YFji1ZoxKqDyU1
x030iGVg2mWpMANRZBtEOkuRbafLTbjp4TXoupSi7E8xMyaJnO6ynbKzSwkcIivKaNVoGG/q/JI4
tYRzCHekb9G19X7yPRNMX2dUpE5geWfvu9wBH6r1Kd+KlhmtwqS0Q18gknzu6wqagU1vBCmjoJtt
4/e9vwqB6PhuZCtE9l/PXuQU0koQ9cTFr4pSO0otHbLgmkkGlrl2GSqEWz3RcJwB4pylMAKU0vtz
xqIeTR0trceRGYF4uTAOLN20CicPdBZoJFw77hw7UH9edpiyZQZKLjTkZ80kQ/+E0c6a49hwyOOf
+t5ytEqiV1uMVGS+T6byFJUlv93As6gbUmmwSOOYSfx3fnrWEYEc+m4Oi7CHF+id884u/LUxuQpT
Bm4xDR3X88cR+2XPd3sol+iV6udhovt5i0rAiyxDydWlnLrCtdJHyrqpEaTLV+/oNJoo0pRL3lXK
jhwIy9kQRE+hCZdBwpOnZd80LLFmASCYHa3sFGjM0eRnfYyAgnsPgVsbHABN/hIphzWyI1kGtqGf
1j6jDrMS4xGwvsjFJWg/2Q1d4rgK+EWFKhQJwB5cj/J0AZ97QzNW0yOixJmU/S/HSAX6gyXH0Op8
0JJou9FM/ExCMnrcib1kbQajHng+uy4IMGH+l8dCTa8LB2yaSxxIwLnvOX5692h+CUBpbOv8VP6T
2eFvhTA1nJBHLt+FNlrN+Hb2ShjCxcT5tCQisvIXsGWQ5ZH2JasttRTq7C10z4dmHUXypBKeSIo+
HNccjXLMwR/UPHVZygXvON6HHWWhsNkEMxKe5kyxFNs8v7YY/jqcUZvfsRrVl0Wly30G6DwUem/Q
JU9qBXy8QTiQ7PZurfpOOeeyJyitpR8OD8RRpKvMdGBQX4M/6Q3nbCoGkQfk0ZoDJ5SW9cGbdBLN
rnpJciZD0V75uVCPXSRCRQ9PccG8lQmSSN7bYrUCQXmKpfnGhWXr9OHLd2VWoFmZT8tGAJmRTxP/
K8OjL2aLNFWdZNHEZFLcnIYNQ32m4ZlisWdmlsUt3EwoHqPv8Xne8KILRS0MpdDfEL86/vDotKSj
IT2XNtXscpKoIpPQ9QbD90JArA3GfjE4pq9ILiVwQEnfFJhFj2A2sZKl/c+TcjJnpxiMJ91uORZu
zCQgOKSAuA9CqFEQNW6NJn6rSonxa0vMW7Q7tk8y2ziatrtOQmut1oB75jDwMTzqytPEB/t/cs8n
l5Q/PdHxymIBwAIbrzdUaILKGSHjEztdYlE6kmKM3gtEuDSXOQ/+SkRsvZ4mz5w/w5cZzx+17RE6
mqBiqQjI1cth/SMss//v6WWerVywd+8ik6EvBiDuJJIMLDVlXIPRXFzmz/VgT/ROWyogx7WAZt0z
soGG9In5FWNEHLc8IX1YqPan9JJ4cHae2yWsgZVZs2EJm7M4dupaHMa3Uk7f5TRXdyaZbgdnFC9e
ou8pq33442Kzat4UJ61QyCKoxKyf97/8ELVEAnlSKQXAOfqwbWzGnH+F5wH4qguO+nlKJSN50UxL
eHyhlusLu7xjp70dqXosTaTaGrfVHGT4+MiJ3Zh7eCUEHZBkjh448cwdIwXmNdhOl74Cs1pYzEl2
PB16pL2LjFx0LC0kCSQLLeAI3bIOAyMfUEzaLf40vtBXGd7bzZE1kEQTJCsKgJo1fuaDIXUUso4u
jOVUpiRNisjIOj3UkESloB6BwEUYIxMTEjB9qjPVeLgzqxE8pm/KaoLHl9HGz7cuQ4z7GCP+fBlN
6lvnZboBWJQ4+s45glesJU26O0DvD5YG6MZOSr0WQUGPvpMLUeQmSQK+lw1pc7rBAl+U4ceU/vk+
OqwUWJt0QcsaeC3A9OFazWtlfDQCo/QVzv6kXbGCS9pgOtIU78KtjXmLrtPWT46h9bKGB0+icKnE
+0ljoBijZNknaEuI6nQRD3F3IVVQ6JxjjabYpzgkjXO/vijGmTJPYTsfvazR62DFne4vaCbuwGS/
ufPyJvIJNomh1iRrj8MZvUCpxLew1PmWQojhvD6zmWKCMKMmD5qPW1+ElvptGaE71u09V0NQ9Sfm
ZLnYIw9lrODbTTllkOeJG2rOPm33Y8casc+qQqDlPcpIZDK5JqoJ5AbGgLElRmHasApKIAheVLn4
tzGIQim2a6SgExkMcAFR1dIKvwdFlWLdLQL866wSB8/FX8lXLfWMEDvmkvv/C0kEie1CsZMnjU9G
Z2omUDVU8g2M2nm1v8dc9LNiVI6aCO0sw496o3K1bloKGWbc9YuJ4k3KT3LP7cV8IdmgnOEctKxL
96QU4NlyCahA+okM9RrpLcMP7DQ2HEtfAlySbWxichDniekgUr/4dnMcnZbJtovY9eZML7jHCjTj
OLUbC+GGddnJIEDTdeFwUOrsRJx30AifFyUK64ZNMbbGmjZF+g2n+epKjuERgyo351T9vUhNxgh6
f/KWGPzbTfiJmcVhGfN3+Fvs/nhAmXVUT4aNk2RR1XoZ4EGfD6+hzxuxcCUo+RMXt3SgPI0U8L3L
xJ3HsOlkZlz7lzEWjwKB1T8fVwFY3NetIdBDJ3lERCIOjf/E66XP6axFmJ1CsI45Ymz8QXzydOgQ
SqMVAW8iEKBbY/K3JfnOatvsGPVGd8z32hIH2q7TXr3AOc3d+e1gCf0sfCTol+t7f3j2Zh1GwwOs
Qw5zCrElQ+mu9H6ddKbRoE1Ppxz//bbKyKhw3i1Uq1N3ciw6RVxV7yEp5nHxoFGmWS9NVgOkvExD
zSLAcPgqfq/1NEAbBU5dkTWEJIdYCNgiIbtDMPP/E7FFX9TCuXPdmHSB1uMJEISLrM5yZzDaEait
z3oFIcPlOolA2Vm2uNeMbFvYNrRrfo82hXoziwKCH+O6LOW5uWES4YKw5JoytXfkMW9ojHbC+GjB
F4Ia3rQWUMAlLc0NOOrypW+Cgx//WWGzTkiVCKGaELUicmTdAsAYZMp1DYd/LuA00ErzmlHSEgCT
6uVun1Cpw5p6aTD4OU5aB9arJpX1uaCU8dS0VY2XuwnZmthMv4QP/sJXA/rwnPBGIDj74+JpoIbV
OVYS5/tzpfeex4dTbd7Cm3rZ4vTb5XXnC07tEdAfpcXohiFDXl9lX0WP4PksVQ81vVuNjNkTyPgl
yWQjoyG4tu49I1uUvyds+t41qytb/HAHzg7eQUIrt99+ppHwxmdSnbfBv2yo6BOpuRABSKN0w8nv
j/OnyTV7dm9YZL2U0j6MLu1em9Gk/efK9/WsiScCHDFNZlUMK6fJqiSQaf/oP5SI34mlwr5BQt50
OzHI0SGpfUkSyHZnTRMI42V6Qx34WGjONeMKrgluT1FVq+R5ZMnvQ4yUofTuFQhNqzzRHJNCAGMD
g43+IqTUS5GdLH6rkBHFX6SE0zT6TyP5fs0WnZhsFEcMIcCQwo6rA7/xfw9f2iqry/9/DoH1fbvG
1NFXUGIo5QXUGcpCh3qIiZOE1s/BpK/WMaFVPhStYkbIbjKcAU7TKRfjxZp8WhUK8z7oaVynI6zV
13ugrOguObRzjWKxzAlfWYo6ZdTaaIM+QZrNsu05cuZcfCXF4kkq7Mslbiul1ttmRCUzxr+BpVNm
uGXQxMa7AJsYO82M6wFv2WJmoQcv7p2lTFXgvkTmGkiv/DNPOnfuwgZhXQeB4p0Dh1C7hVTbvy86
kID5fK6rotGnd5yJ3Iu6iccGTjgGMNvGAvpYKLi29Rj/vOpwicqy4sE94IADd1jMSI/Bj0OreTMr
cHupfModA7t6ajzcS29ZQn7cBFdmc+Plzirrif6rBUG1iffj04dv7BlEfCN4GLRukck/gKE66uyO
PIK06L8AZWpOM9z84nNP/R4lpRiEf7t/AuxEN7S9rF97uUiyTTgTWvKPmdXt/VaTR217/BK/0dHA
u1r5Dd0KlGhHt8DwSlfzkMhwxjMaDUN8bDLBsfPkOVfxQKr0LOViuIEjjqSb0jovyl1gnQPz7zaz
BoLIFTsJWRN6XRk9PVeVdng8CdShFD4BzOhY97Kiur0dotNMT8Ekgmqu7IhrVFqRcyWhb3MCdE7t
XR15odkFZfKXXHO3p5OHyPnmvs/QKPafe0wN00lyDjx5syz94MxIjMlkWDboPLL1oykVWlOMonIE
CTltEvwY/U/Ds7+2GQvw7swiqvIDoz+u5W9VPutGpidlPjhff+EHT9euCbwQLgwac06Va6SGhpEE
w5+oy4An+kSJwuZGNphGArQnQX67OhdWxi13Q5BEIdk/8XKTyRoGimRIepmx6W06PvaWDsKM9ex/
l+exA6r9JMPaNdXjcO+2y6EvYxwFXLGzLsF8F4yREX0iL4FL+Jg9ytL8Z5HyehrZOOaJO7MdG+7q
huXKjss27H6xPHOtUdMkfsYPjPJzPJRZn9ifoGStQ963iLiQuZw6ntGIiyJ+2/tE/M0dDyFU1SYs
4iPI1bS9QFs/cVUWQNgY14recsDR2NwC75cCb2uAJLPlp5bmNMqcgYBHGoJW3ZSPSq0P+CvgsfZR
y31+X9M6bdPCz3qJSPUBZ5Nf9WeQyRUEU3OL+FB3p1DLvChvftDFbjqVXABfWWCSZyiT4Qpe+ZAx
K15s1acdhGvs/bRy89xA7vxgqScnSHi4DslHA9TEOl3vQf4FXMyeUus696Iu/j5rn9vl1kxNCk8w
ldNj3J/oXpj5NLodcUQywQmeoR5cYcnvNsSpkgxaW+9mSclYZwLIh2Dlop190kbixlsWUiOqUOEE
MDq4hPo1nTzEiQxwbXgZEPya0DUUykErn3G0oUKaUPAqISnlKRW5ZW7fKb7AsRHzIfbgisFpDhW4
yKyIIxUNCejE2BRULs4cOH7C4ye2bn1L62DmcPYjPPXbNKtb6EV973LfmlhZ8bWUDLCvktXSQCHy
znPq5I1iovTfoHwO5E5lBNz7msbywXkU9fbRmPK/FmdVz54kHUkuDbPgeAF1w/xIEzxu6h3jQEU2
F7ZYDMJAKsdvpEkkJXyqID317SJKih1p3w9wJCizP9gpcXwsu+++/4Y+7wNjxyznPDmQrGqecFi0
iFKSDpJT31mQDBXRpVQOWJ6Kcm+j8Jv2VtTi4MrgKpIiID2kRXol4Nj/VK4ZAexfhnWifm4wfr+1
GNHAfcZFPOh1aqsi5MpIAycGxRNtNjl0rZEbcAVCACOsJmDy6O0EbDlkTzQfwz2SV5XmRtXh5eQy
M7j/odFx7lRjobMcTUCYi9S6L5lPupfEGNDh25GnSSl+5F3NpAQ6Re5Id2Opwri1uIm3QgXaJQyR
veRbR0fd2Hr8Q6Xhh8uCq2dhmU/k+xs04k9g9zXBGpZp4cd5mRToXmzqK5kf8YBXrwND+ZLs3RWv
3eHX9O4y63WHH9wB1lT8KSdoMleJzhZeL9b2b015GMCFy1okIUtBH4pUOVDa+Ex7PBoJFdptJOoB
uBkkRBKpOrYezta8pVd9Ic8FSTAGbvuuGETQWlnnD/2xnn0BSxrSiBhnUR/pS50sNcwl7nat6G52
mCL23GQGhsb+qkuOYGgL394utMweC5beiJtNWAMRE+hveLlNY3BmgsXHz6hw46e/RxCVzkKMZrCG
0h7rMr5M0qj8dXJ6BZoX3YMJl9sj49vs98Ra30qeSWIt00tNy0hT3o1gM014emsn+aqQAKKYJXsQ
SAgQczHo9Daq+4/4YSeHLmx+9LQzS7bMuniYQjNOeaQeXzu0zUE3S2HyytdTbStt3b3qnKAhWShE
4fw5OiSf4ZJ+H5dv/gdwCh3tWISFXWs1PC4lB99FjAs2f8TSr8UAI5ocafCTKsjRQQ4QJgnxc4J5
LR8Esalk5aYlPFRvII6CjSEZTCVHSiW57hFkpmRlMdtW2i1PAEETTwguZzxZlolIJSQpNZzyN+Zc
umF5tu5hg5lSCn8HsDIz4xaZa9kugV0CsBE5S8d86jdLxOg+BN5A51OefhlsRDAyJf+k+1md9PaV
9xkkiS/X9TFhr955Y64iX1eM/cOJWiIGj5UF/GznNiKUj0ApTRW/7KZxdFNZ6DgxJoV0sxn/pvkh
ZALaxc66izEXrtvs9BfBOR5WkAhexKErPaNDLsk/Cspl6zgs7aIhUsOCFHerZ7nbH+kzAdnWwrOp
uNPG3T43YluJ2T0vrWAR51l2jxTkPdpralmE/j/eW2UYZrSQi1LPKPNpJPFKwtA5n3su2MAv0Quf
nJeiJ91deVdfQwHNWy1yw30fCgh694YqvCWO2kELdJLbv8Fnniau1+d0lJxHPsftpIjpvx01kNbp
SEiM8I/vHVTAUWAZ8U1GW9MRa7L3tchx8unNV9t7AgrQKKh/xGtAGhkqOqQiiHJ7CqN5ZiIOi8Vm
KVAkZYzSXQSrv0i80+vEqEZvXQuvDGcWTb9p/4SdKBBgKSBmkesgOrr0xXINbt2H8wLq+0yO409y
FgsgAdlEMs26dBB/VlmPKP5WrvmMp0lXKmpqaXNfnAefA4KCzMi//mvSqCA+GFbyiu6HDPS99PTp
Ta9RJchoIviny6GRV6fzcr7jkxRY8S2HNeoUNlTrgWdOEFQi1EnJYu1ie4bbmvnY/MrMTEtYQml7
hChfEB9916TA8CKrO6Q0QbPMBOKJqkirFVBinThCR6smhFGlj/I/w5iHPZNtW0yc+cbgCQIvKRl0
gKgix47QT4w+hBEPIXiijKNh8eU7BjrvaPB2tBnui4xf8cME+q89PnGEVMLAPOoJFm/iGJ3Enm6W
bJ/zG3vWpoXFrUBbTa3dV1vI7Tq0xBoytcCvDZhUhvbbvNJdWQqMRaUfljenkBuDQEN3Ob1bSRVC
lvawKtEt7lq61paEE9/da7DIL4Ux/iU3H6nf46+Caqa+ZK05a9O6gVFSZjjySiOYW4avqthUd9tN
RnlARXnSdsIsO8qa+jNiq8v6okDn5JOWJ2Q+LcL9K8Jq/9vvlFzRnelTKEJfXbDFvpbFxdWcwqcP
2QNKHAIssTMedd5IshYaFWk3VldXpj61Hhs7xzyQIDD8LkD5I3QWq1i5KnjfeYzggVjv6UGWqkmr
GVUGcXYwlyZoRgqbvB1U2/REQOEfAW5hUObIa8laUomigpNrfJkzB8izbqDIxazsMAcyPezCJ8uK
C3DdboU7R55+LzEEJMD7mWX1kTdHhc8jltyR22nCOXW35DdgCLIPiVhcwS6RcJw3/K7ZbvF7uCFC
idpiwLYqJLrnck76uV9oJjkE2au+fcO67B9FKahDrnXdUrxcHILaIyNB7KGuAsEMvPYU338csVdq
8Qc1A4ES6A/OkDwUO1/epfHyk2cOtqiQiC8E51LAA3f7+Bi3/xSGijdYLI/aEiys45/xUFDsLwgb
5WZccnhBBsIw7kFpT7jk0qbtQJ7JlOWrOsrslA2F7UfRfD/XTSGc7PvusuY2qo10dHgYkKokXlKE
Y1NH38pUtIYsS4KiPZ0c2S3yl4F+le8Zirsf1Nn+CTxWKrSTCT5Rf52Hdz4MWbChlfiuudBtV0dp
IgYUny+UWQDZMz+iApiDHbYWCMU/cVRcdna2E6c9D6H1+ZsgzjCbBqsp4KAeGPQej2td0dBQX0Zv
AFfColBWtSObogJf1c3LlTXtWmCpVt6/zA+rgXl3BYsN3rSdcM6b84JGFrxTcEUn3fnEegiQFLlA
tr1ajZavhwhDtXgf8FG0iYR303hw/G71f3fSKhrinjSl2PdHuBWeVuka2XbV39N0FgUMniNTeJCg
4/fOlG0jDW5cqgjwa59RBxKDLMOJ4SqHlAYtj0F6kdojCFD0jbqJHB76MEwUw5scmU9Oy73StvPd
LBCQbsYuqNGrJbt3fYGEqqRG+uWP8XlCwcwJAtzaqjyIMvti5JsrvqNWIw9D3SJxwucQgLes6mQM
jaNMBgMCHRfvF/0b59MTfhzpgCoNdIMAE5jYyt6LGWpjZGxPXgI211RHgbZ5gDD5ttC5spuau50K
KZWBJ7CPrPkWUydj7AnLsn/D6kfwn1ht08cytMwCRnIpTd+ei6ILJ5KQamnGeVzFZt5iOS/RCl9n
m3bCQCCIx6JnvTL6YmnHNWVGdrbMjgkdoBxFpaejTCrktXfIiMIGSBfHGqwySa0wlcEXXrZPTERW
IhZCcpi+zd5KnME5OEnnGJ02Xl+Mb8gzQACoB6Z4INU4I5T8frYUlIt/xDlEcL8fqyGgz2Wic0mB
Bt7Fg5kdVctixoBeu/MLyJUEnalLselawaNv5nGpovWvhdSgbD8YqAwV+oI8GHkA52rdVyRmwJ8J
AE7OUiDDBQTfiwgqaG9fcCGEKXumNnocGm/UVn6+WulhY8j5VIZEGGJobEGpj2Dxd8/mh9tl8qip
0ej93ooSzO2Yx08bsicE9u8cu2ns67ZiP4HJ+OBIt9hqM0Wo79nFAZLwyJpNJc/Eg3CQqnXrDxNS
swpMHeM7Y5iyAdHlRd8bfEm00bn2j7/0JB1iMSDvQmnchWUjyFoQ++0XBtHK0u2qzMd+wxXXDJgE
xPfL08KhvHmC9DG19/dh7ygnCPxOHbqADpJWk2ePnkXhLJdeCxQG+h8W1KqkXQIMcxKcxje2qBaF
SdI2JPLXTgalXmPQqsZTp7TOaAwSC5k0Pg6q0l69LcqJ9D6/cx2MmwoS5nleFCQF4gOT8aXjflPZ
rL1A34vOnlWytRYnjkvdwBG8RkPiHckltGSEo7HAT5zKN/E436ZLFcoTNIv1t1NPBvMyuv6BwCZ+
fRQ3+bd95P7OKAl6wqn8Ci8VRJWCwkVQR53j4LLRLck385VKmBozzWKJLgwekLCEVvifz2M/KvpO
EuLX8uBjsLt4SUpwD58LK5x93FNaICz1R5l9wm+uhudMm5xYgQrLXVhvXvb+D2Ga07YCzjzCo7J0
/6PrNFS0Q/u2MFrBvKdGPx7Rul2rZEdRCiRP1jR/X1pSgmJ7uMvmfDiA3RkDAPMaIKE/f2FPDNcK
nxZyqQAgsYeqV9+dSv+ZL8lYGBqhpsHOTDR5T/F1nTqzLKXzuOyZqGSl6uduCs9ezZK1lmnxzZst
IFb/Wai4fUvYrHMzuQeaQMdbL2qBk1YOZAmVa1bGWEVBOTeQiDD3Bc+6gsIMDGlw8qN+jtd+skTp
Hjn/jIU+mjfbSMovn8Qee6krS2d6IF8ZryD7kh+k0eC6OmvRsWBDX9Q2AtfzKEcK40WjHNBID8DB
U4fagFht4FJwoY06SjsCKSp60rUbFtdGftuwrWuLqub3mmppKHZg+JRosP8IavKGC2NnUVzfGwoS
g/HiMegUgnqzUUW3CG64HZddgNpNp67pDlcDc6GjU311dRiPqAEcOLETeHKvf4uJLiGp5iUpe5lR
c6o8wrvXTn5P5tulXnW44ZW36wxbkawIGv+9woYR1QrgEHJYfEX56BBx91EoCmsEoa6KU5xun/b7
7PMsaWRUpF6ZO5z6S52SITVqr5T46QMtiIyL01axY3KywnOoTUcwyEPAel5YTANveNiukDYzeEPN
niTlbZP6wQ5KSVxZ6BV9IKERjYllFUxxg7509rXqMs2WrGRnerkWmW9+ZFT7N8kRaMaMkMSddRR4
VztGWvL6xBVNoRTkZjIEMGARnFGuIpks18+hqTx5Tf1aTL4p7FGm3/xwOzlR75w4fKx5sYuPEqYr
HPhm11rrZygIGyE83UiGW1ohjWim/tMWVDnIgpgHhvI2TmtnzTTz4J8G+YlZkSsA7fM15VcTo3OK
wlw8X8v2UvnIw7DLp/sdNfFESDPLDfOscZ/LPyWKfjYD7OeACMtaZ3fZowyDZUQF/t4s0YtjEcOI
kDHxWTF2LA/sAbyBWR48Sf5EeA0GbZXKtoOFPhh7NGAb1VtXk+4gW8h3hroNJH0Y1P1Ysps9ODzc
50hTpwqXM6GbyISxwMP+lxM57+8f6VhqF2pu1d5VFJJX6A8Qi1xcNHCruFzEQgNLVakNWyWtMuV8
dwkLcjPrRP4B+Nst8Y7HMGtchHQ9QKVH7D4oIURijIkIYcJK4wLOWB7aVK+zv6DU64buo7GS3OAG
jgT/Px8hdKC0RUtjn4Gat/0cwr0MRmefBQaoYxImVPn7sHQG2bJosK329iRpxhMT/pG59XNjm4Xy
9NsECCfZ32ZtRd487mJpa9exkqN+lqfB9iERRoF58fYBfWzEaOq5zD5vbauVXlgKtC6EmAA3Yb38
C9U1hmMhNzfb26H+psgsxhTzd+0y/0r3Zss6AWpRX47QJz3R8/vGgXXXI3/Igk++YArWkLFvSzvf
LdjAuKG9DoU7Vt48APw1TNfWgddxwudJDet4gjpuBJPlct9/6WBr47IzCHnmuWvzN5PTVwlEPJ5S
ejscV0KCBpnIjTjddcRiW+u4DybBYWHAjHcW/rug9CVj55rRGr7UJFdB+TM1e/bIE+ddb9EZD/gc
u6uK1lR8J4tLzg3ErKBZhwnBW613rUvbH7VnRN6GOMC2fuLGzp1co4p2Gexq4ct8M3BGMHHjqf+N
MDjTFGNvVZ2gmFMTWp7esC4d7bgWnOb4C6Tn01PTmPFcNqilJ1veAYug3HR17HuxZD3M0dRCVZuq
xgpswsZVgMVW6eRWDUf2+yxgjv3xUer6ojYThe6mSFTPWfYZdi9/6ZzEgr2rbmo7xiUu9yHYKR8Z
bJvtMXGejX8wk5Pu9fd2aMvVe3/iGyf+u9L6Us/5U/a6AIkXctxg/8k3KpCr5km90fm/9JwiZISQ
7vtnTCzRlzxTxnFWrioelvNz1mEp8riaL2ujptSMB5ZyYH5PmxrQveMwn5ktViSNYgr4C8hWCADa
oALdfG9SZGzE8ax6TOfph5Xpfwk0CHWJ5oWr9i559EKkO4Y/HtANZDEGAJITiPHe7Dfmz9+WYzNC
Nhr3J5kmNap7LQvdNyBkiRSufge0obcNbDIxuf4kyktpDtRyGhZ0DKkAdZgDpqZC2yIisSVMusCo
w6hJznZT+/nCj/5jYzm8jVHyIjiK6NFe8X5X2DYstvPSmW/x/RKJFelFIsPomtTGJ1AjNa3Ur7m9
N3s2P5q84H0xfCiulqTNaOZTw4eQeom0kjlFmIQXPJUJYhUglQL3wtT4iITth9al9YMHEt7wUpb2
c5qjLi+AosIADJ43pwWl77pB6Fbovacol6JLeMOGPkYRjDkosqJHq4kg3qWNi+zwWZePcdRK/p3k
sh8jc/Wyj+m6wSUryX9y8VEQWa8+xR1T7iOA7MUBiXpymuiwiP234g0I6gU2417WQThlvMmicdm2
K1WIgTqCe1KT3QnU56qmA9/o7LBKNOGp99WiixgI9yKYu6o1mLv7kLHWCzpQTImxy9npwqc+gyx+
USGEiimlXlhdty2kkIo85lfwFDY4J18c5GTpBOXHHim70uWL724bSxymmwO2+O0/X5H0qTOYx/oc
VR0iOdkMb1v2/7aS40sAmiX5d2DbD28APc5cRxYD4/4kpUIXU+7+99ag53Pnr1PRzKfzDhMEcFxm
lbxziQYgGyHMAG9+dIA1IzFHY4UeN95vx0noJIO2DEmNdpR/onh6Eu714gC3l+0AovHe1xJDPKwQ
AuNWhofxzn2J8dziwI76ERWsCzKGg4wBtYPpYGxmys2bJwL2kPSx+47CZEzS10mpLkhL9nnTTzLs
zm5HjYHY48L9l+MIHiGXoxP+A18+Lz05zLTRUMSOLRmDnft6bXKvhXC1Xp1wmCtCqRp9CYEGLLHY
Cj6QPVylDz0S8uT9RX0vjJu/HHhLI/qhDGVvDpzfG6iezrnkEabqrO3ylbOB5m9VB5ecMN3jfrT1
Em6WjRed7EVm5iDTmHynV5H9Gtgq7W1ALHSLHAA+o8i4rExWvcs8MXWqfky8cGrjJFQQ6O9c9G0Q
xf1nR9ztC8+8E0hH0rdCBE5E+awcdoyuITzcVKsn/bp2D7kMritD96IRj4gJC2vnzmj7zf0kdtQm
MsxhYiZ2ykzyc0qPVXm2V6UE/8+tHsDoOVZBf6oj8Smiejli3od/t2uwvpeJDw/AeNzHGT1r8GXv
wcN0X3I9uteZeFf/dmJ2uGfbdngPUbNkYOZtYoMDBl4yAtwF+HkoD/Ta7yfgUcFup8TlaQERO0+0
CnSOJjadz9re6BF00xaYFV9UoURaXo26e3+tL2gEo1IDmSlldpNMDtGW4SOBEGCpDQNJqvGiA/sH
V9pb4BrCsy83pH8vw7fnLz2cE++IqgLt0guGm+W6PEdbPpCT42JLnWXpDJU6txtzXXGFuNq/lqrr
t5reg2Nbt8Y3mQKkrVkzTLfUKP4pa7A42Wq71NWb1JK7QtZ/+i1g8fglYgPR1sfbrWDvk0wDSpwn
OHpxnNzTur2pGY6S2AqytE8pG5dSQG/J38zTESTdUiyjlSs8yg0MZBreurhCOiI4CQDRljt1dCyi
ANupiGEE7RA4kYWAlCssmJaVyipsKNnpw5lVA6WNgn5PQ0W716HJ8sCPTNhGHuSL0hMhEq3bMZqn
LGdcCDw3A69ms3/Kt96wRp91tHL3dNCMaRpFjZKvZxBbzDhCGVb12PTGZi846OPgtS2p/GExnX7Z
52sHKyoXFkhZzKrTddu1MS5S+RXPyInLFzdc0h4SoUPREz55+sO+916YGJYCbTKn0fc0e4QN0NFA
CzfJjBWjG2jgzVPG/p5PsP52cwCoFGG5kLcF9UFV+6Iqy0G9PXl8VU9wfrC7kswYnh7S9juq+rxS
mJuupvgIiW4AqxYibJIbfhxVBNqcHAtAnQIsJZVOccJR2L93b+A11TUrGFnx1TqIhdk19N4Ia5oS
Uxi61t35LDkUVi0YnGbQFVe4jNfWe5FeBla9XPIxygX19CgsdRhJuGRUtkAuPitnddA6jAeQ2E2Y
rSFtbJsJn5eyoK2OxafkqcmI5GsT+OcXzjb4UYlegEHwSx4m+rxwHaVgfN8+eHfI4JUzWHTn5WIV
JdbN5Hn6ae+hyHQc52cUMqKCBPPN8F2NxLhmXYLqLiT51EZmzebskAFyPaRVoo4JLSjPnRnj1sSG
t6G1Iq3mPaNnFZpl4R6O2vto0BDP+6/vosjwMT077YqfsnUaYGzR7+BHSMKVs9dn0jGppGK6qEpP
ham1xxMF4SZXJUQ39ANmRz+HbicXlXXl9fhQmLOeyruW52f1BqwAUbzmQ01Ty0Dr9fvWhjkM3ZFp
B8S/e3Ic1vFiKXywtrLsIS5s3DRyGiCjNNRKhRTu+GUKErJWisQZ2PLXiBnoHC1OsryiM2n7Uxss
Cf017im5rTPNlOzfGJ34TIqSlTrm+Q+2qCw/aEywblwQD1DubydbNjgNz9H1jJSo2EVpAQunK9yz
0lMIIFWgnTaVQ4mZICuj4Qt6DkWh6uFhrm+9PnU+sKduLSbuw+RxDn/n6oN2G39BM3DvFJv6buyS
HSco+W3aKjj3NL7yD2gzRK3wfQAY2d65Ti2/gYQzw1dfXFTsZVfCOTkGfotRBkLznvZ62faX2mTG
RMNUz6AKfUUX5ri1vUZF9MknsZgvowrD4KZqQrmPG22fuR5KKaYs1YBs6ppXV760HNdFLSD+bwln
P0B/gPuTxVcehZv/P9eUDoTWp7/TD4f6fr9OtvFx8fo63HCkD4zfQiIBMebt9Cmm0+xLizXH3I0U
Tc1kbzZEFcYZt1wt4wdPKr/V9Lco2XsEyTbE3g/n9ztLza/a/7Y84SqgBge/K9hiFwqI7lXmW0ct
KoLpm4jM20T/gf6qtF32MqcjhGv6ojH5cq5Yqb3JDIb6ismTr4dkisMb+TLu7cqqv1D26KYLUTUB
pVsGMnYc/2+XUTQlnc32HKHv1UZ5oPirkC9KksZMv8JzqRln+f4U1frXNXAKpEOF19pcX4MFRcKt
fj8xcE0lib0Bhuj7Ri3g9iKgaitV9K63lU1JzfPCOxzpU0xHYe3j9tWCVezjU+YiaALLX70Pb6ap
jzOmchdaNEubPA4L7THY5H33+oXiFk4aiS0EjXidv1KcTNE6QptibLR+89iWuaqt4fysWPASI1Mt
5bXKcx37TaiPjbANfC2SKOfjq6+Ksl2uv9f2FCdqUUOoQOVHBA9IjSoHXYBF29UhnGWLY+BKauTD
ZNotD9b3IWd7G1mGHSW8LTCMdjqYQ1N549aNq011InQueHyhaR4UMSWsTvB+b8SDRo+JLAyrFMWr
ghOjz8PBm8U0+na5PrbuZDVXbSw5+FOuCECOhE5BzqhKTcmRLBoyhbl2DRranCy4MCxb7Qi1hj0/
9SjAaC1A6wMjdRsqnrxfMwK9lnLL7wkR8KHNtts0WlqzFKW17baSHErX1xkcFNl1h9ropZutEldd
Muh1S2KNHA0lu4gcqYvFiVeV6PH+44QNQR4qy0cz1rgz8WS6lykKhumC7sAQHAxVjuPrbV4ClTdp
UbKRJAgFHY6IQ4unuIug0Hq1DO2Bg5ZR4prQOawGAuPJGSSjGB0rL0cgk6osAHADSb8K5FgIR4DQ
c9O5ns8PkgJPMJemJcWP+d03skL2d2wNYdy4DzA0HTDNQJV83umhE1FdL9Ops3odk8Geei6+qQvP
YIHBEIl+0tIY1MUrqEJdoVi/scM++AcRj0llqi1UB9Bej7P4V21+xASXBE9Qo14pYkNh9+Op/SUD
UNCyqlrdEUrKRGTGl2/rYg8bgyoZKmD9VF3xJyPhOW7GMCCcrVgEVh4ChVH1ObKPJxxYA1PC36OG
f2CbAdCDLPTlnzHBqkHr1n4aD8Gz9rO3g9imCPep1DlFZiCHdAmlDLVkL1FiTs+p+pFL0kyapasG
WpYA1CfWh5UeSR3v5lwctenq5VhR+JID6b/9K+rhUow8BeMJ/RUM86PPeMq2aXrS4KPTZnY/LxDL
0C+g8To6jQTrz3nYOBpDKcaV2JeZwviWHpYGL0+5wD4Ic559w4gOAI3cUg8Qhfd14wDEcCOEs2AQ
O/RGpl2D1ICOCs2eHxjE704VmYHxOAGNBDx8ieyRpWs5KRQSy5drfngxNoDU/NlQXtrI0DZvIHHj
5phzPjOyNFCD8PL8cQolwWKhxokldZuSZjo8wA/BUAsOIozaWad8ZQI7NMV9NbHjON4fX4V89Wh7
zIxTeC7SxK0NCRwwitzu0BLQ49VLbdjuVxHzUPnfmj7ohczHZdlGrvL4+rLMinPfpWAgJWsKbTZM
RhDL8dROFkeqhdHg0QlA/ijTgdh/jgJjtADxw9uKUnlOsnnz+cArCDKMKblSnXxjI/QdRgcgYThR
mOv4Pr0Hv6VnESL9PyAfx11JnvsDpRnO8Nj44PtrU4fM+VKHLMM8lTAg13JNMrnpPE3GxhdZILra
2q8c0R8r3ESLfpYo59a/QwTEfBqWUoTxO188vRCiNV7E/l4FIwDKCx0kBgJ7DL9eePQZG5QfJeiI
5EbSckpLc2caO4T0kuAFe0CZ9y6CgTYKyIgGlCP3KmzxqHAE7rtiR3LlYylws8m+VwdJ/KM244HL
g4LJT+4tYggZmg4I7BO+wReFLY3U5d9TA1WEm/F/F9g/ODgW+Wd558JS6qRi2uwrWoqxBQrmLK5N
w8yEAdoRU/KA7iZN0oD/3fch328aRUeXBbpvDTJNunDlaJY0BWwYCPTFv9cxt6kBcGnUU/iVrCpF
KYJcb+vNStp5pTq2HBtVNXFofrGRbp+kNjXjlfdP/bw2K3fXqtFLAVas78XLwMIea6HyGcISQ1Wd
GqO8YY9KSl56GBt7SyvY8/As5Z1RnJnliExRaBG1rp3KOBIRVfOI26/6GZfzrYMMoNfRr6A2lG+w
sraaWBWl4ywPnbdsE+XwGQyO3Wy9HMUpReipN6LQZOED/vmzNqZSrPRTINLWdgyqf/7pJ5FcnKqZ
fbEvC4RK6JaEKGlGMsaeImdErEYeed4LbY0gmHGdiq3H4V6S7OS032/hs458xoSv6OKSdWkwDsR2
i93rzG4d7ezhBz0+fPMpYI20OXrzgvDhBdRRtfOvRCJXh/s+Z5kWNX9YvkT1gaAFAh3coLCngqY9
awa2/zxPXW2ql4A3taOiSmrVq3i9Q35gdR20tMIjz7/eNUJVmJx7qK0h+DVEfUNWcISpC1RHm5rU
QNfBpKdaNrv2rNEtiKbgbydmuio07TMgynlF7fU9AGhUnefYdFQ0/QTq/hWzILDSdd7cQXuw8nU2
aL+VsrbFq16Xk78rYQeDxO8Rsdlg4Cm46m1c7XfcxyBF+97qlI+amtwyaNiFfTrtN36px6qe2BYZ
OfWfWrZikoAzuP2gMdU0VlYh52E1YgI6jgdAPEnCTD1J+Hpe19TEzOzbWnLp0juTzmIuk3pAMIiu
I6VAjHDby13BvfgnrkKGpLMRPdPoOZGB5QetdAIGcIG/parVfam8B6CkLnQdveugae/fXsO8CaLA
Z0hcEatjZ3NMwnCdavHJGfyZ2DLCBTjQtPTP+SXwvi/YrPVhno7Yct+neD9ZVvExUtoN5iOUTRyX
XKXxE2RXPOw/jTerhtqH8z0DvX+g1ReaqolBSCRZ8fzyaXa8/FMcsLBsdkFaacm+TBbNHrJ4az2L
b6LBwcCnUa8sbpYF1rq8Adfu0ur2OpzeJthhd3AlMmTfNGsKbHS5O/np3vYxBcTF4wWvXuVW0I8J
24Wo1E2pYYI9Ma6zCottW4+4yuGplvkGmhFddhpoyFg9qL6KjDR0zycrpaJaJTi4dTTh4wLk+JbL
bJXCZhP2OuzDCP2zIQxTv6i5HDxO6NKnfNmH0ZJ99/IrR5Bez4DX9cFs/DBUckuCYmEwZYarahYO
pzUK55QlgnZCLMkSVw2+jeOduRD29QxVhxHxbMUJCtg7yOHFBSESfmC3uK/7Csy/pYG99Rq1By3a
h7MdAkX17OVOjtJoubgIKlfp6pqD3bLZpNyeT3b5lvn92ltRPq2/hoi0XwOtN7MnxkvRVhVM1pSQ
K41EOyCcIJz6CtM7rV+Aj5YU8MPa0bEeMSPWig5ZNnsSOX4BESvGK6HoLYpXwdX3nS49KXyhW+4W
1IreGnS1D6QyGldZTgPMcUf4EaKUMFGyQI96ne8b4CVTiicOZEkfqoXCCf8Eyp7hNNFavE97lmhv
v098r9Fi8mrzXVdP8SjRKSZMzqEg2dLWebYHOeqYF5wAjTh8zcU47uIKQFFtXjs0e4jlZ2z4xWgx
7HifuXkq/VCMPlJ0QKn6oes1spHiQ1Y5td3firzX0MMvSbNCYGSLUsZlYYn5sLfXaCKMr2Ai7smO
fgD4O6/yqp8PTo9/pP0mthUNJS16OjFXxc9XX18Fq4S+iGJFAtYMnCZL0pxTvZEdot2Q4d1DucIc
0NSm2xRY5l6XRt8VjL2RhHnD1kzNGbpNaEb1duJQ864YFABcryidEdWlLzI9DFbWCO2Nb2xaqaOg
fUkuwuJXM5qlWQXI126G+lGMT144rl2WZPoVoIYXuwAiegRoEM6RzZ8w0w0uVBwriQa9wepGL7eb
Q8ymjFNAv/u/MhS4BQWGu35NEwonmO8CkJMlOdaxP5LXD53TLzLtEuj7i5CfZMZBNs2UF+iawP73
Wi0c7M9zWzgYxQXjjmZcdbNPIWXpfz4kojeVbSEFBzw2Trf2eKDqt98Mru9gkAzvyvlACs+B6mGb
sCI8ignC+Tnd/woVfm7hOEKuqectXL2pVCyqjYTk0mqdo0h3xA2hkzJIzLM68LtdpFls+UcvepK2
GrbTy+LVjjHhbMUpdz7pCR1XahY/jjgBF859PiWNUS2/7aHoX3Fp4ElFXdE5s2RaySqas7z276tW
WOMlbZgQG2f/Dkc/QSGwRTwWM+VkQ90IWf6TTZCvj2idT/sYdwcQRBPvfmuVdUJxOn6SrW1I9kUe
hIDNpyYAR+vlQfYgOsJEq7VsuFTZ021ltFTDZKiJtRjNA5FnG1er5/w/j2g63wuEfSMOjl6yjRpc
j65pSo98OjnwPmheCTazHIKTW+eNxSEB2A6yg25aH+cOdz/ZQC8q+Ohc9k0qiUrTCobn/cC3wFXr
iPDqHYdoef8eEPPCpl9aaAs39Nq8ywD+Y4kPjuUosbxoMFSEKTaVQVJFm6VBaKfMGGOGTj57FXUP
+hZGqbt1AGZ1+Wa6NoFixtjBaUM9TPiDDk/O1NRX9Q/XKPbBDy2P3Iq4opT60O+Rw8o9KCITXfl3
ib5YAzQArjJwEAnch0VA0KEYTlhLhVrbzFmGzIQSewCUxz39UZeAtwO2aRkPkK2+wuFstB0DXGXz
zkGUruPnug1SjNYQ6NIQhTej7GTj25IXTeN8lOdj/7kE7ZHU8xEarSnBxu9YxRLpuRiHuga52Xcv
5dqbW4OurhfpLksiW3V0tenddWrkN2g1nGFIlbMDrJV16joUchzUgE5X7HJC3I1YMR+EysgtWQ/1
I6qnVldXsM2XWQiK8yXIXGMtFknIgL2RwnZwHINWATq5wQMHS7JwWcqTvdpuwpdaDZga8JyAtWFU
VdyxpJkAWuIOySLhZrwtA5PRJRxYOZ1R5+PI2CpaPQfR6qeByLPXXqL0Jsbe5yDpBA2yJyjD4Wh5
NUrdKo7AeJ6/Ma7/vvUl4p76aU+7spnXlNlQ19XwtjHLT99f1U6KPgxiK/HDqDxIjmsMSdQczS7I
FsDo9hPk0Ki59QI0Us9ZuxZ0LDTEgOl3XqwSpdl32GhEvxXmyDGJgXr67dCSKafuCZng02+tIJYN
JHM4QtHom7dwI6F2A1khGmdjIAlTdjKj5vJ4t/Qq8Tzwm63U/nnqPhS1Fy83TEy0L1UiRW/ROrCS
b2u1bxjJdN7bU5fHsqDZ99DN/nUcdUelUhZR5ABMTatLWpAwAWU8TORnmGHrIgLlIzoQa+maUfnP
kCYxKE0gJo1qrsdLdIUkwUjo550YYmGDwHPlOcMh7xNMSbzjZbFKOAN8jCads2njWvYkGKW7VhVD
lrLXSHja3UJodlRgDvW9BwtmQisoW0hjEyYdmALmgLCjd2lI0E7wl36ElQecbvAi1Y8mAiBt6n+6
icLfLFWVZgh71labAlx6S8z8hWVC1UTeRBgSxpgH91uSZgqkcdA7wYd1SdtjK8szgBG65W2Ltuvw
i+x4tdHvVqQ8Cgdxw5t/xyaYVGuOBXXarB/QfHcuExJws+xgnPYJJhpwMgwK3bHE0Ff8puffdetm
Wtbkdr6A6jsIE/Enon7clRtyXfUyO3aVmDOLDEn43QCD0OwWfWfTRCFnMfEtQ6aayEuq3eEMu2x4
1o41xGEzojiTQG3fAr7kKHKa4uXEngfJvJCD0tV4iIKwdw/YXdw6CMLrE8I2kWfmE1ulLHUi4t7I
xzog9SVTQ6pHCSejBH+FIjI192CbF8xuGmh/m4GypXTTumbQwsnu66sdISv3h5rN5VRuFqgbL9CJ
P5vOroiCA7sQkfZorChueQugGAsT+tz8Csr+i+3MATnQ9UxYRQlTs5rEAjXevXdZxZ3IfEcgx+Vn
syfiauUF8dHTsRgni0CBwPGqrP/gO00WUVnjtfNnlmWX0rCyLmr91Y8P5CG6qeE4/UhAgllTGnmD
SmRnyQFcYcAkW4Ir++r2Xpn2bQcFfVeDJQDO0WEwqrOBvQYanTl5yqQgxR/NQPRjnAzV7cFqk2CY
05u9vgmXrZbsO9NoD/Y5bumtw8VH/vAXq/4GgRFNqapwz5svef+HO59v3edueZsJTR+ORelE1GlU
ZqA7OiWKlSBHmPvraB6ZDwoEnfUzFHeQFrr0vdhNaOQgIjr82Dv0pL2I/ORjTbG9MfMTQuWu9+g9
+Lesx6EUvAhe7LOriludx7IWwBvYMVesk2m1HA2cI8pyHxNdGZyX4UzJAS5R9KWkd7q3T61fuPtw
hbh6MmRhRarXiazuopOsY2QN0WZrmxRMc7AvDvcujAKKZnFJ+/PGhA3IVvoLXIbFm6pWX9OrKSqG
pCv20T0W1ppwGa5oEe5/SkESrkNVZiTpty0rrCedsMCrllHmw/K2s66KpUYJVTgmalnOZv/6yHW3
tZnOO6SMZO23EIKysNpGC0AdM1OwkkBypEsf4im6Y6k3SJAQ9SKaiENy0T92ECZkfzuCajoVKiGw
/kkfDUSlRL4HVSdCyBB0XDZt+AXE8sg8+E0uZE0mgulKKJ3bmIVCA4vHRtVeD/QD6DnpXRGjZw+X
1S8re6VypCl7Ssz5QGgJBQ/ozb0UU3MsgGr68nSbribesm/Q+gIjjFC6KWwSjzAzpjcK//nnRKOZ
bi69jkNjnI0/T1WKTexgK4bC+4Ds4Ae4W4/bwk6jiF/wjqGqIp4z0PRHfYq+RAVtS14HhAcGV/j1
IssoUaQT75T2CvVGLGt3S8x5KDIJGRywwCgN92EL+gbgj/qDp3hHCyMy8uQsC2jbxMZcOciTwvLz
3jR1BT4yd7VQabUp5TzAaf7bhgT+tLrDBFzyqzlOEYYkswcfB95YtPIgT/80oQkSrX7E372Eu8EZ
RoIkOb5S6HNPmKBL6BAYcvc5wzYyOl8pqoVXD/rCPNrc78ZaNPGGnZF9/jvZ7MACJwSuwvFz/4Ql
JZxF02UVcfFy3nCFL5C4LQX1LquL5YtEaQFQ37bA12CFkuHtMe+xNmfTP72AVK6nWm27NAs64pXq
wBns5RsYwjAyhNMXqHCpxhbXbkpXxfWQl/8cSUhW9HhGtTk2O/fxPkcvHyWrUYSECVZ3/DJXITsY
Fd2aItJJCqeiXags8uZybg+Og27n1MiKvXfJGbs24rZ1L8rnASlicljrxY6PR5v3CjFZmGLktTkV
ZE66/7jGggnTfTZfQBZmyce2Id3ouPY1YpcbF1vDnDzAHRAifsTpdM69RLYqdZu/RZi4POY4/VTz
f8OheSrZJ+ZlKcK+K6Fq0JGi1IdSQsfGUiifZe9HzzlJvMjiOXvfw5LmTdCIpiR0eov+emcdlDtd
5RlEja8ITcOaDw0RLc6yVIDUiJ8h9O82DF85ZJUV7mD/lW1HMpkNH8sALTUvuLew0qm3rWg+hUWO
jWUKef+M/yiLH+imHKV3jqwgOjKyvShKOSWjNCB14lU/9R21+zfMA5oyi3f/HzQqySUvG5f9QfLa
nANmn9KDzBHeCGG0ci6LHVrmcj1PCbvDloOmQOHgs0PKwZG1WvoG4jdMnqulM21hhD4OA02XkYSY
lXVFSqD/JWLsbZZcsKKPYtufmaxJ1hfdZ+dpfQzeKyKLzZpHTGZeNB2F7CjkBGxKPkuiLAAv0Fmi
C+/rrcmCevR58W4TvHFT6NId7VOxdbeSKfliCW6cjKUBTBTJo5i2iefz/kZ/Xr2sTbBkw2zPaSzC
Trescbe2bznjUC+ry5iNBDaUtNnJPuL8UacAaBspqsIY6+61remKdBow1pLD9bMseqi9NJ//x9Bz
AK7FuRG/2VwPEQFBX3C8S3vk0KdYWyyXlOA9/dsHQcUAE8Wi9tO6w55de2zkxTdIv7K+rH0vhe2R
eNjiwmuWcSgBdg+MzMlaAdWX4W97NlQT2YoWwtij3izwVM0ayDQX4fLsINjShjj/IqiH2+PwaPEd
u/VUD8uTB4vSoK8icm5vD2uW2sHGEjKWX0k/GG6cpengyajzpfey2DMscTjHmRzAJ9J93uNzg03H
GXuSBOtYR1/HkicUIalGRfQqDXqTh3RldkLU+zpTgK/svdI9/HMwrr2m8NCfANYG0VLomcK0VPgj
oUITcFYyXkhkFKONQhFjCXZLylHSYG8Pczax0VAC/LNPg8MJcsraKKUvgFnkn76ZhsAzFe3BjpYG
ZrrYRL14L8YTmP+F+s8FniQp5VsNnaNNKpA+nBpPHqdR/ezLgUc4UyduKDWZZ3jUrDadxt8ng0Dz
negBnMncy5ZU1S3U8OsaUetQ9QRTgbE2UDpsgrtN9/DUrgUHZbq328fSTIM5V002+l6E01nqlKQT
h5aSa6Q3Y9JKYmhXBQamhF5wKov8ZyDVChpTmSovYVh7/nCF2R7RSL+vZDajsXm45lCAsBuJBxZC
8yBPxNtDod5HTSAQK5GOt7VdApJnUWL+3/8ojKwfrP9cmVBPUQzl/iHWfoFRuS99+537BIiCENSR
3RNGx9p2kIwPcWTTdazYYJGOA2f46pcMkR8mHJkU4cguMtxa63wgl+sXTT9kNrXbpuOPUX8QFBbN
81VKT445B+CWH7+85126P3a2hGBMCkiY5Wmqysyy3C1BA13b5wp3vlZ8oUgOkLRNNue85avBMkdj
1f3InOZFDorE/XG94/LOV+QR9lXrjOuIvxFVK7oQD6AhZ0mk4pRZTcLPFr43eB/qgIefJ617vl8g
Xv778lM3j1PDEMPNX2WXn4em9qVpmbPJChWccE8QEQliumlsc2eA5z2jaSCE3siI22S415wtYAty
Wye27zH3tQB0fwg/diVjmk6ILmXgo7K5UfiX2y+kUirWdW5J+S4cS6bOaDO/S86AGUkgeVttFvdJ
rIfotBwPa9o+k8flqedd6SbD9zDhKtSZfeh9tX9O9r53OaVjv42WM1EER3IX1XF/uBg1eB3UEUeS
2GzaQCADHL3PlP29qrflnflFg7VjWUC3qXCuKL5vKzpC1O2znTWEMVif6aQk0cIdPG9dk5ADCeZ/
PD8qQSI9nzkYfPHA/ZEQvlqcDx6JrsU2fIn7/fBeVnk4PkjwN2asDMI7emE33ubNMToc1HM5F2uS
ePuC6AlUqnxQAN++/vvxK2p18g/A2Dna8GF1zg4giYJb0K4JPpH+4hIrztUy9ocHJC0vbm2jiGaN
2JSRhe4g0/hKp4Bu7PU6lkpzWc87KlFatEaQdz4F1MOIteJbiKoSVYf9/CeYWS6VIBiDUWwbrpDX
5hdQt/l/1cw7+JY7Z4wOP1YeOjVEe4C1dO3JEJimxxS+PgnzshZKLOXKTwBPu9MSBIjR6nLA8q1g
ESMogeoKALlio9O4jdMMOOFuaW3Zb4xflXOn4J+serXq398xbP03J3cyRmd30EyuxlL+Ad4ws7t3
Ar8ggNprAcovCkvH3v8e0qPMx6I3+CI10hhNlTpt9DPlWgudtL4mg/8ac2vsdB8vUhvJAsFswCyt
8kQdIob+hlxcbfAr3lngA4wvXtoNvfZXUrT7DxqxJ4kZMzvE2qhpU9KqqYfh79DPbLyyT8tfKXwC
EWHA7Mo0kHgNTIE3TpwnCFZ1bA+2mQ+CfSJTA5/DUQbedVropCmXyEMmY/A7m8Cyl9Nis5UxV7Ny
3B0JimwfYlKvXmnczTLZhWoa+4e02yyMePDh3jcFAj1twyWi+xpZGoQW+4jRoYU+W7z76sNxyA1/
5znVJyWdEg5yfXPpZbwYWQul7Nj6HU3e2H8H5NQc+WxvMLtkMR9lYXWsUlUCdh/Rb+O+CljXP9xL
kkULZQYCwS0i8js17z6t3V6U7CHbT/XW098rYLbIZJRXqRme7W0cb3QA6k2chDNCE18AzY/g3llU
mSYwHIHi+UBshQrwGHnJFAN+QFIOL8vRCt/jxb+UL+Wz8Jx22HPV6m9TJVKOqJUWh3vR/3wbRSgA
JY7yog/O1ufwUBbDgeIzsv4J1NlqnDGrg254mREm/RK1Ixe75d0TJZYawSA/0PeKSQ/xCjyHLk9N
VniuQs9fF7VLIbVgDvTA6vGy/olTOl6lD2k2Hk+tbPc5ZpWvRuEKH0EkrdfONtnHyF4WOUcqr1SQ
mKQk5hRrx97LLSVvk1PM64zUYJhg2BxKimLwFVdlWn6oHoKBgfIihb+N9xNX6FZutRtyay/ALdyc
wpnJF39NwrZxTVKdXzUPK/bmJBQk+0DRKSx0MZOd6+1AZ2EeeOOhLM7G70XcjzKH5IITcAOmEZjD
jEijPCot13u3+ySVz1Q21D8e/XUq5OlSXVHno7Xb9fQ3fBdxGJEmjdJeiwbmlHaKbSBrtJczeuzk
vCpUjI8NW8w9Qq15Cj2IakS5XQbQPbF41SfhFkdWgWcnECr2JYwFzlW0YShkh14r6qNOcUk+/qfC
5TJ5EeZeAisrKKEC70/O7geWRSZqfDA4jGUrpvrp2c+qntRCy8rEMm+SHHL4b3NGcNPcTuPQ2no7
mSMuaUyuOqTnz2jlsWimR3HrVygsz/+FdbqczPumnQoxWHga9sBHnUfyi5i9nlXd9r+HnvIimih3
To4Z6u31+1DppqEvLGOOKlW5UyXldw+7DXT/ZJ+8jG5Rgm4eQyHEXv03zScJ+DXWo7WDmPe02S9A
CjOPha6BVQi70qctS/tFpw02QpT0uhGcYjLYZupQAH81n90ZcSmYAepmU9D+enErAiAIdb1Y6WIQ
OMWFHwAV2wJU3jUtlug2cMU5ToR8Iq3RXB7j7/Z8gHC8f1LP34nCOL8Y74YSy3EShCVEBjX9aWJS
v3PE27TJ78Vl6W2Db2kZ5KqqxSEwgPZ1RHkNPpCc/FdiGerAPIRs/lyU8Tt+nKnsMFkvgyFmkf9l
vGbgfYmbyMeK1yR0W2swQgaukS2bs1mbTWUAHiD9vsqnR2fj0gtfZaoPEKXrL65t24HcaKQ6RWH0
0+/zYsRpbvGiNXw4k3nepHTi4B6qKz0zjiHU0+kOBhtTjQYRiITXJ/VqWDP4xnDEo1DC7W0ce7IJ
u7njXnmNZ3Z6euf+KFfiJ46ICMlJFDP9fCjRu4aIUvb9pBnzzMZHCvQoBuHePeogAbtueqTY0uue
cogFDBqn3U5Sek5creVod9zmGmAbpq5swP8h/VEnHP/ahfRAeK7Qf9Ix9AKni5qQ/T8hdVM9TZGc
4vq1FeUD3ZdnfJoBJoG8ch1iRLcHgp7ORImZCTPQR8VuH9vfaNYJhKpJjBx8xbVzfM/FqwP9Up4I
5slVm5qH5VfuOj4oYfj28FiOi7Qv2V2vHuqFPigo//SzrslKJRfY+hO4hcsLsOIDtY706B21tlon
yk5J2me4nsaOIGEk7GPrMBJ4V3d5MlGWYIbxsl2XR6/05rrDR5z4OIKww1JMPdBoIJ0Hln07VewK
1ORVIzoJRnsTXG9Z0vSEEYKj3leRuQk/SD6aph6LN3pWUwAFV6K+BrEA4m9IqAiUCq7z5mNbkwob
mnJNTjaKs6tobOpqEAQx8L7jdV4mHptR6a5f1zBIIqjrhZtmacil1hqR30IKxwHufh39GTQaQWds
dn8RgETk/rkEg+xLvgjAqf7VhjVTJYh9DUA/HOsj0QT1ReyP+3QdLmHSpBExzpiUEpREqaUwR6cK
qE2DDC+hjNjj9WqfB5MhQK33v+qhBpln5bCjtiYYbOFUX+fl25u9hob2YonrdPdJ8swjWNpO5pYP
K+mT5BqrBPkRHANomlLLysjjJQ4w2x3MGEynelbq3epeYF2LZ0HUn1XeUYqs/AYHfF3KKTTLaLmu
NPVP4/Mc/ZngHCSO3vMek8+Ck6/xZUnpqoMCWLoPPVF1s1nbE8aTgNbonXdVUw9poHjU+ESDHII0
D47jx+JSCyFQvIX/gLd1Pny+O0m1sck3Ibu4hbai6MF2bqnZQTQiS/7TjrrNZ1GDEpw5d4e4hBdP
3lu6aJ2jf0Pev88bQ1D77o+cIxPeRT9NvGjzSzTOwUlSP7qW517LP4+1eypnRpyRN6WOW2qEYxBG
bJ0HsxG4S+Fo33KMekgbQH+Wsuy6RB7ij8Bb/136N/KXSjc1IqXnux+0Jj7SniU8Xo2sGrt5f2Yu
CYsxlDngfHh8grIyB6EzNoFG/HPOZuy+mCTFEEcwHWmEu/4/1CLg5tGHhyC6nuvBPzLJEX62BVXA
mwIqW6rDJjusgEcoQr/86uWE4DVaVRcQUSd4Na6BuHwZVyhZpnzjF0Y/JHFqMgfHNJpFAYL3MFRr
PtgOQ4vX+FDmM/MbolOTgNtPJLGw8plfFCf0jL2OAFHrQcOk4k+36kj7r+dFEZVOwVHCNzC+U82K
Ce8+zUOATzxLDj7NK0ntNVVEWySvlDvgJen8PTVweMWBd6HqHE3hKGDFWKMgpK2ktcF4xOSkG+ZH
WDAjoFxUfSz6oIQm6U0KKIwCRjnbp3iVuJwIfyyj60vfiIgO50Abcv5DyRVGVA9G8+P2UQfP+ouP
9Ai5zke5NK9eDj0rrZ9lDakElq8UnSn3dahrvZ6xZI5AkVgLrfyaoWpjaM8Znrr8KuCiY6cz5rKH
OGNVlWJKIDNsRUgDVhHjdcAJCG3c10EmiYyzRJL/Ccv1to457A8Q7NsClL8GVA3CrorTDBKs3twX
oW1WXGj1QVbMUn1ElCQ99e/cHmc74TAflCjGvoeYsZrLLSk5268M/CXKQ72fYECWATjBvDwqO46N
C/zoTNAvgYB9WWnH2uxU19ymHKPxfIa8cUWAWw7V2IbrXxQRH+6Oqr/mKVlkjNl0dhnrJ/xFcuqg
kO9eLg8EoHoJUlK1YkcAJ+x1JSsLLUwtBydmOLyWVphT0NiXfl1QruVlxgAotpL0gE5JYjfxMDRx
MIagoke2N8YEYm01PSIN76WhQxqJPQuQg4wO6oqSWXxauZ3POq+UrVwHm1YNcXHSJKCThLIYroV8
YN7yGrnuqwyIfkI7xKo+Z8OxWJ9PI2xVXRD0IkyfTv7RwtsuIstF59+STtVnoksBDSpB+lEwViGW
VSXgoc6/MGltqOAjOTOQ5uqjEEd9x+eu4gYf3B3HgCYkIXTXualQ5DuxV3rkvW0SJbsYjjgyT67y
c0mW80GtWV8FBJJusUMhMTwnG+yQTZJOqXp01+ruvyTDE6qVcbe/CrumuiiuikWTdQVT5ROkkocK
qRoypbQSkqU+7c5Kv3cnKAM1q9fX08KTDzmOw3K7mGnOaasnb0RoMM9VWCl0Ol6DF8mmy+Blvp8p
PtqjapgEyeZIrjhXjZWF13CmkA7tHtFHrD9p7+LvAGVWmE9ypCukT68+D6IoQf2GuPjBbhumR0Gn
vmKGYM/fpYvUrBlpuXsViVWN47q10dCb1GtzcggDygcl6iWQqdLhOZ9AYuPg2BsS75MEsVFu0lAC
ameTdwFTkiBEAOu3Ojvd5FeHnOCreKjJUHFfaanXWivNTLnp6SotaKJPDF3ZcZLktveneHNTI6Uj
3H7xniiVXbjEUKNWlexsIdrBRtOgKb5VNLqZxAN2Wq4YZqN4F3Ok46cGxOah/Tof5OYS17UVc9zS
ZVCdJbOm3YT1Kh+8shDz3zLJ4jjS3cjDxvSGOy2ZnGS4Drwx0ZocqHTER/PTg1rqwsPsuXm15A+w
pRJZf+/yYiKsbB9EoqWHnl9sT5yhDOfnL6/VxIYdaZU5WOmgVHxUvJE/Fxr6VvsoeZhliEqryxEQ
SRerp9pEOwuAsMWG0evHoZoKDuWrf9NCCYLi5vfXjVUy6cJ3nSivU0GHhrJy+1APmhE2ZE469OYh
SWk2dGQFbeyFqO5AlTS59GuAP0ePZ1NKiv4Yeemgr8E3iJhRg+Hsv38LO+vKF6ioR8Dk0VFYgMx+
oOACHAt5OklNpFD+FeyD/kSDckddztyFOHiMyh5Znx3VIE/bAVghCYIMPwonx/cqIBoMRRhSS7Zd
H6XKuuSY1GH1G6+4JE06vAZ08w0Unuec3Gw/F18NozSbQ5C/jYBa3NMjBLdUhpxDEmtP0GtGx03r
piqrk60Ar5zwScNutM1sgY+OELJTXzmD6C9hhC4LUb4lZiL12K3gNQRQ+fDM4qZGh9AJYB2LFHxk
BOxx9XJIEGmN6ZAKQCV671m1CGZlLuwXM+LX/th8lkOwPtuXPqd9ueoReaRdeqNxjxAePbrMU4+G
d8S3kfIxkA03jM2iQ//M4azNkaYNv7dQrqovRVh5iuA1Q5e8BKtuVNTP2W+Hb7ieiZmtkRfDXCHT
1Jje4mrSs2zLrnYQycIPjdKAakoXgaSoEtr6PLt80kUO4U6gOe/YRKO0doPyEohH6lF8pZDMtyAw
jn18f4J3YBWiXvXPRUMOM0e3xyVlMtSwv6OC72a16GRN7TmHo8WbHySoqLY2oUsdhEjX9Ra3st0w
bfdWmFK4pQhOE8LuBk3jCpCPKD0WCd3McSo5Hs7MUMNtIwx8nkkoE2vkTowvdiDYam1jpblgiHmV
3bL1AJtdSvS+bjRV9DbS9ErB8Ogu1aBCbt+iJsOb+73FbYmWPUMnIRwmEEwwmtuVUyl0NSKeeRRg
Lm9G19yUVcDK50bZrhVEdU41t2SJZ4rrPk68gVofnEQNT2HKRq+guD4idE8cwzaivs/3meYEnBSA
FvkQUJ6/9wtozvouB62hke9i5zx0HWxutl8sCNNGy1yNIQAzaDa4We9LSN7K6gSc6py4nc3CVQMJ
nK2CFOU3ON9qBhp1Vj5a5bcoFb6mDMsWLY4MFlp5mmIuxwmUVFe9/Xdu9S5rlR/Iqu9WEvUaEzL1
uwRomxPz5cM8V/2/XLbubLiJtrtt3MAnFo1dKDTQUu8Ln9BZEJ7ImeHQZtGCOWbRnDjhifreDdRM
ZssgNH8TWoAZr/4grYxMzDDiUzImtQDwSSskn19dgCbm6u9wbbnXUgOXzHxY53hh5zXaCQd2twDc
Saf2Ipl3l7a6oKeiIDhChPdFsVJ9UxnMmY2Kp6GPM64HALuw+I3RlAHukteqxYdYZj8vPDFhS8dX
y1Iwhd6HtVQ79Ym8ru5PwzYkJqTxRElVbtLcu4ONYlgDC07UW3SUE+rIv5ycg+KvzgcoqM8Fjjte
6GEw2ZlwIasUgMnfZFv/L8xOPtBvOyMkH2Y4r3LPMTXBhWrBRoqQva0O+jrbDP69gYdp4dsiPkAw
J2STUTMqCNHYO/Je4ALq/5sdJnQ8V8VLZwvdNDapVa4Ey4xyL+KDVtcsre9NlSqUKMYq/37/UQsU
hdjFBAGVgxOnqmTk6cc0Qcy4pSLymVWNPGAWINZ8syuO2/wRsvY/BQhywbrV6RHEz1Ar8qH5M8H7
Kp9E7scKM+kSbewgV7ugzgutWwQfYaDyWkd2izMRtO5nzpZxOLK4LzkVgY7up1wxewSFb7IcMXeA
eihp0NNbVsnDQ9Ng6hN8cclqF0IHLosnCeSndQazh6lMRNvD1BZz7nV22Usn9PBy/Hcm+9VwzJ3T
wKZTmHpZ8bxtN8u3uHhi6tM7wq1eD8cI6hSfid3H4Wnf4WEoea3p4bqRrjVizf8/z18PrqeDLgdt
JbbJbfndJgov0x/Vefr7Bi0a+9BmiRsWyTs3CIWuiidCobTafxmGTrs4KlLnGd+oaf9X4trO9/gI
pUnkZ/QSPyiAG01YmqJ0bf1wDDeI5ZLctBjpB82LZxfGx0iG/MSbf34WlgCq3tC90DxX44WEKafX
QyKfR9mhkU94asy3dW6JRA13QDsySjMeSe0sP27hi+74N/Cqzok53+JLShsFXcnDgwa+0czRkVCx
shmSyGtAjnAl1hNR5h/Mvw5vlfmXOedk86qBX4rW9jGZvkIzEZUBuaPzF+mewyBb56sNctd0CVNM
WzxdB+iaMi9Cdwvr5/LpHdDfly7Tz+BocF6L9HvxeRBx5KZvaLyBOmMtmImerbfvoJ+7siy3rEiw
2DzjUJXaSNMHZtX+Gxz1CC5dk9PdE5NM3onHxhUJUApxZ98zWCSiGSA3AleM68s73MAa2Ikt7M/4
t/T4Rz1axLNCju2PQoXuAX90/A/QMb7+hWeStOH8cKpjshdhtxEA6sTmbP01KJ5/iPOz+/g4dmh9
lYN5yigfY3pbsMeJksA0pUOo3lgxaR1TyG9N53PfM2bq9kyM5U1fOyD68MhVnjyQL0SblKk65pMm
hGovXcCpEQIXVtsPOfKYgKY9MJT2wdrBlNI/nUIqouDTrmxt2aTTYcH/sOEfpT3BCggPux/0M9L8
5SdxStfk5EfJ2meRJp3x2xWSVsTbJH2qqOfNFZdmK5H6lypaz1UNcqgui6DBdwGGRU76uUz0fZ6I
LHaHEKlJ1wn2KnNChq9W0j/bYTZg13VJi5YCY5B+MxiI09N/nzSgyHLWfq9K+yE4fcV17HhkUNyE
6yRWmid1GvtCs3PD3gRT/NJSY+YXkwS/AUy5ZqJ8RdieCTeTB31oqxXfTGPLTExU5zX/Q/xMjblo
6DcEls/67hbkH7EM3nxWZoO6oU7+VIUIihXX5tUW4ls6XGoUNNkyX1M0tUwwj21fQppwaKSiIPPh
DdOx9WjIVN5dWZVS9sSgW0VtlRLjI4AszF01SoYhzQlvuo11Qef9qjFsKq0Qumh2c12u9H3wRxuL
TU+zhs3PpGVUYBFq2ghW06RrPZ+aA9ialKF0A2cyZD0jpYseQl0dCeCRdqnwYSg1+9PVTm4/yh/R
rPt6ueGXAPeO7DgMdyRPuueJ4/oWICMpM6pKeThoCtPyqGie6uXpZvMRr7t06w94mUXBJ21Ec4xh
XvUVMN9uUngXo7GOd8lP3p4X9tOnZ8mVmhY97K759p+z/tB4d8WCm9DKxHUGB3AoZgcucxvUhgR2
3UvpWktstUlBa6KFV+isyy+CmTYXrImMmyNUci9yWIdw7M3WvSHjwWY4PtPRPIPz5UDHftPB7tKM
Z+k5NXrJeJ5hhW/ory5OY6Lh5w33TsA+HUMSZU7WbzdKhioJBWFWh4XLQpj1/Hte7Lrcq1xxQh3R
ytorETXMcUP9puBtPMf486OEtGTmNmUzurfUk1UOiYXx413wCut5kPyR4oj/bfpjl2NJuTMkWxD+
JmAsoVgxz27xafBd1bAPl1ACAav7mg2P093nsmrxnKYsEnX7bzuIdCzeG0cpt2GjheViMZw1UNm3
638eig+00Ismw+8tSCMs5UVuiwVL3fTZria0A8W9Nb81DNIihdC7plA+KXmmW64xAiXrEOiqiS1Z
krAaOTltVEiFS3Rj86PscpilJLpdW5vPWH3RfO66hJOO2bROH2dHafF8eAGvMqBxQvKazzyu0OOp
lNSTlzVYfM0mF4M+SnZvYwMs0mU4Osyqiz+NsKQyTht1cVP8oDP+aTi9lLBEpKV9KvQ8t+k2YoXQ
m780W2PydytObrqJNEb7a3ZeEqaPSFoA4EH+w2ONpozaw80XuA53zHMg9ODudS8QoQ15zboRBz5O
lW3yzxbmfTSRk+VgoS6D7uP14+IRzjeGlKsYSYlkvkxgNkZ5p7HSYfwRsWzQjPGdJMMT2Jr6j7p9
VELCFLHFAIKZbU09tMtGCpHiCkqMtxvVD1fJTMXxAcsaJOJR5+1PryeDJbDqhyfFK5DNxQTF48Ff
PVHP1jtxTjQQ95mkyEO5TvppTEtQtFLPHPTGt3qjED2v44+kCquw93Bln7Hs29cExEVy/AmIxf36
Vma96VKqGLaS9Hw5TNryB1iFj5lzWudirBZkUGuMN5dB5hqTG38epeh96y2mUlFCrzsiqZOXFq6u
x8NgRy3+qTLHjnVl//RV00Ebl1FE+JCXYQSruFPQ2cpOqpgYTRBJ7iyTzk27u2jiwNAo9M8Zi53k
DUmtHyiRkOsvaVDbJ7h6N2k5xoOka+AF3fYm0FP9jU550Y1qpzbEJtGEM2g1rZB2yg3/6J3Ki/JP
+1ayg+XnvWmZPIuU6ad1432YXfXbCPyk+C23n8WqOxgIDHRVx/DB7dkaknp1aogDxk/3jsBwa4NH
OrqrNjDZWQNqmvXfBzeNGnRCpbyWYslUUtFqleP+XhNBenleU+wA5sJdYFBNW3DRHeoP9tboj2xg
6a+1pJ7E4cQdj6qpabOq9YSYrnRuGM3bPkSbRLPXH9QnRA5oHZzLo5dvowMedBjF59l2OOP0G0RD
ZuJb4eeGKRZ08w1Xfg6ctocxZX0Cd9+TUwiG444ZbrkwbX3kwkePUaNi8B/1rDDNVRuRCR26eF+z
tCIS6xAWCWa+ew4f2R53lcmvWUTOKBXFJtljPdsSO0WoYDmssy0MTwsKvbubqiTWnddbYFfUsQRZ
mX5TAjDU1SoVeKex8CuiyELChBTi9l+JV3+Aru2cWdtrOFMTRzfoGfUewDETgmJY9LdOVciHgCXM
4+mpv7cNU4XBADTiPlpPY+k5uNeWB8EXaVTF6mo4zNPxQrb8rWeqweK4SZ/AvLSJVnbgH/tCp7hY
TJGmjKsvzAd44frr1BYzVcbG8CP8jBUbxGpDuXt9LSVnnd9oXD56GRMnbjsa0gzGH66aZ9nccOYB
KJD7Jsbe09aSCX1guSjXK78Vjq9zPr/6ZoANWk5HZJGh9Z09iOn3W66dvQwEwUbR1a1pXcJ2utPA
rMr6HXqZr/fUQK8dvVHtYkQTL1wCKFedgXAFGAyy7cc+plavpeCa9dFExBAdS5ynapXG8oxgjUEO
NVy7iN4pLHcJYI9qLhB7XKWfT3J+eG+PlI+f/wORcBpo7AydT0fHm34iEBKnTUSRrY+IL2e0dajz
dpfwG8b5oafMw6XB2Jythso/R/2q6hEA640f8NraEAd7nSNP81GcrHZVI/6MAmyqQgJL7tJoDJku
4UeVa/L5TYkE49Ko+59S/4ZAm+He1ct+KF7CH4R5L5J9zFBJ1YJe3LPqzLEdg2dNp49f2P2O0C3S
77YGL9/twXWJDl4B0S0rlxuQq8Y1QbpzEONYyOSsWGU7Y/Gzb/gqR9wA0LTOeefqXgSAI/Afbaxq
596xR40uIYSE/KT5NY1a0IoaRWRxCenmeXTfXI7N0yRByPLVVgLjkBa+pyIGc4bu44721n0U3tA0
u/oQV5BdE8/SF6w2jPTPXCI+ICdjngSFwJw0R3LQvvivzNgCxg1ZQD8Hvw1LMaegydklyzCKK1cL
jXa7oFGNAHcvjBsNzuBBQgH1DKwZD0XqobDVE93IeCCHLyOJyEI14zHuOsx+zYN2XpqZhTOso/nw
iD8FA4kZmh40pd4W3UNYUhYq5SIW83KZC8teIqRdqvuo6Mzqg7PC2snVznWyjRHJeKA6bKSqJ85I
RjMAIqoFHx0sh4cnrBDSoOL0a4Gy89qaLOk1jd4v+eqMwHswWNNzHPPQKE1WsVMyhWKvByvKx2I3
G7hYQUH7CBls8Mhhr0Nsmjfgq+PaAMyR/kiWdp1FRtX08i0iHNbj0lnWQVvRUDsMonm67v0zFoRQ
HuzXs3R2+la4e3NKMmP3sl7DoHP3MWdT0am88dXqsBUJXTHFhrgySYB9L0kBrNW2hwVtYTFBw5vf
Lzq5BVi+Hnai6sbDvULXjSFJh00hq8kyOGr+ulrl6nE9YoUtGyHOWsovkV0VvRvy95WdVA/iAnp2
UqlD3Oj2egdMmnYtlvf4ZX5jYFu94w4JyM/Ff6l9waE5zcU77EY7+9kshNh/KJ/gZTl7NX1qVBvT
KDXbfPYAPxmtOOyCTrh7h3w50KySSGWW01oDZR+CzadDYndMLJhKIwUPzW5r6ws9k8crXP7Pe0L3
5ZAzOxsgmWyuUdfFm4nz+HiZb3Xt2arL7BNbmPuoaTq9S+5wv4jjiuTMA/gavyY02REN1jB6tx8/
DXjsddoHXmaM+4mftuzGLXsmphfaT3MnheEcXhXpL01WsslLvXT1RhgAaa5oqxz1D+xGUjRCaq4t
nJ3KB1pyCvOqlS2MxWjuhsxM4e7yXPqe7Q+Hn0ASs2jHUFiTtnrSao/jxmQonGFGUqh3yxsEPC9y
7FSZ+szLZx7ctJpdjg+G55eW2bVSBly2OWzLdn8O/C6MjZhV/9pM1cdcjAmzEAn9WzC25Hev1vyX
XA6PTvxBj3phNELmusmOzg+x+K8HviIziT6tBXOmcXgg+1bZmtTd6dGmyYFL8KaOxnbJydVSlVr/
GCGa3kDyT+MvbUTLlLVtRK+eCCnmvFDLKmLA/QvOgo4PmZ2S9ydjL6sKH6vxwt2bf6lq8ZgorQLp
RZiRg7MAmD1fFBegYadAsUES+3a0DwJNpDH/m/adaMecEIHbfAIhPdecP/3WF8/uFqvIMcWr5O22
69pGBUr+hBXXeUPpnauF1CRa6aA2uiQsCU2F8dNW/gcQB1PxyZX79fpqRz7UCcxXZ6GNzVwFSN0x
1tY2CXTdXtxghmrlT9GAh6QlHEFT+ZYlwYDgLxEWy7AXb6GS0UiZ/7ve+w9Ue0c2g43VHBbgrB7I
G/C9eD54QLSGKXupW/SVmzZb6mG+EZTKMA6VpYd8LtnxVF0kEWgYxXdgCqzfZnMiRwQzIxhOSRhW
lDt03E8DNB3kc3VnlzDCIL/1JfRKPhjOchsGuUTuTR67OlJSrRnLGEPup13M1YbDtcOiGjzgnltW
3eaEvdfyFh4L0XEAhNfHCCPRzh+IS2jOec5ChG5bEo8SptKt2Ul4PHGVcz6lTp61nB7l5J+0kP8q
K7oJq2+DAk3V9etURrZgrNdEiiY4/zUUU8WvO5Liqty7XEu1uAGSlhxpSpF27SCro+n4PhlotS8A
tfUfCWfknUZ7hAs8MMrzacR1TlgOfqHMoeGo4QSg3WvctYdjRbLVSzlTxFLeLIOtj0WcoIuQhSi/
ee1sw96wfStNdwFHhreULvzscsW+0t5KN86g1a3S5T7JBSp0nfAo5Ia4sBymDjm5npNBn0kPBisH
9e+sYwVFLZTp+DzlaBDyP3U6vDyzpsCN6R7EfMWOHLi3NWQHrX2EmrHum8C8sQPbaVigCVIYmuW6
C39A2zQELJHzWedY3pF+DirtmT4UzOWxIahfwi3tvqXVS+XXrhO/yAXs1YqtQnhPu/eiMgakcJDB
OIPNAjGFRtjrGqbj9OTIBmcgdL4atidrX6AmmlCqQsXIVq5PjpHvGl7SeTI7yPDH3AfToEWEkceY
go2GhUUQpXzWCN1sHj89Yomly3kokMldS03cmidKrg1pQcAzDHPeKK3rro//P66TVvA9MCzTbewZ
UvpzPwFZED6vqYFHhEWRooAvNCg+puaSNEO1i97XQtwBj3ZEL3/WhcxG2QiTJuLSQTnohRilp2NJ
sIvqndvKZIW0n9BzuKzKIGHwUWy0VRfnzOw7Y5o5b4qiwLqspSI8D14sKmdkIu+c8Yj7mIDeTfIF
TCR0+iJ+b//BOqxoJQNnhMLe1jBLbFenR2BeXI3YiPXM3CrlSs6L+8B+DbKmNCcS15F8SjkRhSr9
f6P+QFJZlSMgfecAzxBb+xFXm6hhhEVFuDlNJ4q6WIro8K79UVVfh6pgdHGQ8xXg+xostpXzBSwz
bAZth2ExJQ3KzVwiReFeldHARUiqP8OnWh/YSrAscBLiWGfEV+/Y5zeRe/ZgqCQaGXEL0+d16Kvh
B2nEudGGoM409bPzbIiJ/zYeZwxVvRVquVr2Uqrt6J1C0kGMnnQugroyBjBRjpGC1Nqe/b5BlUBt
3wViymmdqOM0U9UitrCpQqs17APt2wWg8N6NKzEWrIup7zKNeP7R+q0p+4vfBRbibw9P69Kdcxwq
YfEoI8rEQnT4xlaT+1BoAyuuqAbo6vx9J+uBqDaDnB5g0TNXqtt4Nmi3v4qh8x1VvTo4hR8GAIXt
ByrVhO8sOYne43fNamCpnBTt9pJY3HCpWCYfzaFRshqdXzOqAF1H4ZHE6N/luld40Fds6xme0ec4
7v9DwQ3fzV2qnWKAP3c3xb+ro5IMRRug6tiz+N9O3DKingwbrB7lBB6KIGGuGQ2RZ0klM7ZtNNpK
qKkVI8c5XR5zP/hVCs6BNwic0Em890WnNjD0lp9udFLz6o63SgSC/8AF1LaN92HP9w/KH8CIt0ES
mC4sR2eEx52cezJEAvNdSXICjSfVjS8WCNPQvwQz2BB0BtZuNh0LFPum+NETVsyzmC0ISt1FJI96
o2r6+Xp1fEVIwBs5IZKXDKwjoDVsPndWhvaBR7CSIndZ4MbE/s5NIc8aZl+TbW+e1GxMYMdqzaz/
VWe5+qw3QsV+9W7i9NqqBjU7aNEv42ygQK2AtsNw25voSqvjm6rGKebm33LqDT+qGwauVssAI2VX
JYtcN2HH0KQWoDDLagABGLOMpK+fl7yAgABZdISWoxru0OpSMCvTw2+u24yNam6+5PeSc+Cc+G1C
tRm1ZxEq7WSwZ4+8/lAfQwBdEoM7IfeE9wR70aFc3ghpSg/Wgx6fc2cg4lg0RHAzzSFQ82Y/eRze
K699BeWvKDAJDF0VzTmppTDrLo1cvbRW5LrCLFhvBTUnSNa/LsWXgVTcW9NSr45FLSF5uU6PrdQR
F44CF82J5B1qjMFz4Ey2hTgzipUHTdC33yFn7pJ8Vx1Lal527jtIJm/epL99N5ZwE4DN9MbtoDLd
vQ3e4iT+cKJOsZxzjBl3hDvkzUW//a0R6msGRCs1ygsK+N25sjKju7buxB5FZooIM2qRE9NF1pFW
h1/kYGbfoAT15ZrJxqA7w4/cfdyUEdww6CBW1TDvJZIQWmRCcwI/cn1EBrqK51oHbcxqZlDlYHJA
zjku+SYyvAjfWXI5s8JS6QIA9hsjWpuF4fQBMjCV9tB5jLtGJUrRRYKbde9e4NQZc21EdZIMAlNe
Zj7/8gUUvMLMTl0CmBVwALtqXV0EKuNlZ7wWezjxKr5Qd6oDxo/iyA2F7CUGk/Uun/nAf3+fXIdD
Ans28f2MYmtRRvfA8S5TA9z0T5thruVC/VN0ak7MldRj0kRKRygbkL+WBv+S0sbf+5Y/e9e0KzOA
4aDblcw3alEir3GORhiJYlrgpObsG57lILZdfYKEr2xkbedVck5/s09Xbdg7BbnLt7s+aR8NKDtL
XS/O/brfZZzFxLi46XFjuo9227to6xXJzOHxfSBkqmREMgnnDwbvOQ9dq8PCbrn1hWz6Om9V99iH
/9bi7oaKqfJfnxrfKYcD+wMn3gUJS3nMYmv86flMDRSn6b5ufpyfDop4RI1WrlCc7TvafQYtqq6P
n0QRR8hkEqFoCbxJM/QauqOyhGO/asN/wrLNNREPJddytYe1NM5+spXa+a8aV6BkwzH9ErE9Mdz+
NoakEfOXJr9LmCj7ZYHN9fDLyKCB+nKa+XIMvWF4q+lk4Y5e3D2/F3/bgwyKw1DC7JNFO7OzVZNK
f4J4f81f9HPvDVjKTl7KO8/JqHR+oNs48YtSNSL+LGspPAFUjiEjD+1LrY1eeBxqRz4sDt/mPZKU
wnaPIG9MOOVPvu37EazlPWuTngvDpDB692rqvFXNcFnsgoPZo6fZYeM5W85TNSDKy2v8YN1tF2XU
oR0eqbVg4FHGckYjuS0uvmVwgmv1ms20+zYjBudEEReV5y9/NfEc44TfCYFcXvX3SIPbeLY19vuA
cnTEq3VdPO5MyUlRbdIaAZP7tbdM+FdQcngS1cpEW/GJfdUxMOQ7HcvPHfIW4r2faPi/WJdV+zh7
BtJQz8msPb5lCJAb8iIDkcaO+H07X2RwGecQ3lJeq6RRFC0n4kw18pysYCkUHQVZkYc1AQFElXh/
8XRkSiiBFE66JfhWWDtThiEH1ZyAVz/epMpgFP2JcqeNv8pm9aWySYkUQb9rZPAkkCegTlsokIo3
lqr6BLW9iEFVZDthJpNbTFOlqPo9hxLpZwLPmERJiZRAAIRVk8NJh1VbB+lPbgR21pLjz55ehjRB
UcdVqyLpmkf251ybHqyoENRnds9FW7YVxdxlCqwWEErZmhw9KAP8ANY2u0FtNuRND2vvoFe+P94v
9IfsVomMlXmwbO77p6UUCeMf+D0/61Ug5892niHUKCwGCO1TR0dXr7EesyMM3zT9O43Ei7Z4g88u
PI16xcEInuLxg/pXUNvwDG+mkD38bZgINTvo36kwG0HBgXerSwVOGu/GOBFtoNEdns80/Xs7iMJK
hNeNTt+ZFXC3M9hDyZXSNj0p/8h0cRXm8qfUZnJkEhTy93AIDlS+AKljZQYB9NNPsMAa0Hyw/3cs
XEO0/5s2ItydJyXIEbpba+kN+l7GTb/QRiklddYNs5+TLhjiLMJ4lIlxDVAeCa9amn2VvPb+zE8M
FU8VzWvuxjbJqMHF5AGwgD6+EnDntp6nAwfx1T+Md5TTTWgu5Bd6ZIKd9iSPyXeRprH37ZxVtnDt
hB0ZQTBcIrxgCgcpkhGDlt4d3u5O3J1nK4OEJV7XIqM/IQ3QVHQR6HsNCxarv9NfClYMJFt7CIIX
2oOxgj04bLIpgUKU8uNy1wGedvHucP5VZcWmIbqJnt4aBQmLBSS5t/4N6M2YhWPr1HOQPEJqWixu
hurJtx+FWYYhSTBDePzRFXIOmvVTRhfCfIanpbKirR3Rb31WW/PbnBPdZdnWO8Kx+CbbMp8570TJ
dNeL2Yc/sXH+SVwBvAo7Vb86EhfubmcmbDEAnWI28ExQgSGQBA1DmCpSX64RC+EZVCX+et3GpS3s
VReI9swS2OCWTfY9z/TWsXHk20YK2ZdEoaj8Omw3aNwrZ6BZoLDei5EH8eC4cgBxVR8avqT2RcZ9
iIvCfSYoTpOoMKuEUy6ZP4odWNE7Xmtd5oK1azzR4SfgtSAftdLe6yH4ff1GxUjKcdh5VTW71YjM
/mMTC0YcRC0wwWLXicmJU9ZI2ex6ou2sdoprGNTYeMSVrTQKIBw1hHQjV74iMSmBSdLYXfidNYUa
Ezouap/rbPZ4LnrZkWIGFuC/4rbeNRWaxW6d69WQQuEMgSKe41x+LTtYkiz1udm32WhkNkHzRJxO
2TZTRDOcz5iAsZYM9Y2wpM2+dOe59ifIUtZJ4WY7MUYXTwZynEpRzkjDpkPtJ1AatzQTiAday3Yn
I9/+3rfSBpBADhIgMbtYGLtlCVvlv9AZEr+9UKbJe4WqGtDcY1hJ1YsWDZ019jYNDdbiptqvZL6U
DVWnrLagmHmDrJjrIIsabuUaHf2oUjv/mJXCClG8K66jTp+U70JZcdlCXI6IzQz4ABtS/x1mKvSQ
v2NrqeBRE/pRgoO5SwIFys4iWDzWeIJ+kkBojLh/zrYh9AwU/mYRZzBb9c5XCpbhhlpYQi02RYc3
nRya/BCQYIP0Ct07/DRi7ktSRI3ldmNUrMOjIQnwaR9Y9m/TlTwj5Cr17rW87jWE/BtzNRrEuFPB
5pNvk3iUX2dBLdDIrJFep/Wz63wMoFyc78tUdMLsAxs48PLt6Z+qQQiOMXLHj/Mqh9YRQXufGRaE
MPX9Hp7TafFReLyucXljBeXOncqNpz9G0XkMS+NDyh2fJQL7vxaO2DrNxEz09BOFos/is5C8bjW3
mleqslkwvcl98toTt9gkfZ5M4SZXjKrMbD6FGingXV6qqMp0ir/F91gGj01NgYXQqYo4DJUXzSTb
VYSSN+A7xk9QzPTJ6uxJtU6nbwiqSaBjvX/gvexW/q3BKXKVDeUSNKIVTkVvDgR/mBUT3TjQVWp+
2Il2VYwjfDoWo3+IlXB4TzASs15bPjOE8ZHPQr/Vhj0dViDP2/njmEIQ5KNSytZy+VShSYToksG4
AMFiJv2g8G+2sNjaVLq8+OZDTlSRrLQaTt9jUbFns/Cv6I+sdnjHQ3eNtaAR59QJIVC8wbOGletS
2newssthsB4soTyQipjKNlFO40hY86WdReJh7pCMLjf0jeK0fJb9ITSWjyeF537OYJr0aqJ4GiSO
tUzTN/xuZF43C7qWh1ZcnYPpRmLziYuKcKEDi4P1hNxzHBt+AtCAJc+we9BFFg1Q7yrrjpntbmvo
Wg+EfBn/oao/YvK7pe3zqkXHcYbU+BlDn9DifSLtQ/gqOpL3XEyj7MOXVraR93WqulLAiCIKbBFm
vLqSW707EhWy0ZPsDel7rNg4SINIiILF8iv2XV/Blrha3CvyUZChAR2mzln2ZUeZOvdsZrz1lv2K
2JyLoCRu2WJCB4AvMCrHh1MVwIfXfsA48vh8RWA/VY8II/6DXiDyk7vGRVnxl6m5U0u+xemfHsCl
w7ufI+dUyjBcfAyBTIK7SJ5M7O66s7cyvSwuZr4tFeEu/K0WZS4pqXqgp412jitdcjk3pcbZIvf9
koNs5acFm++6Or5pY6hBDPkW6unwN0mxPKiKZFD87ZIweoqp+Hq425ABIeBt+qBq1U3HZwY/lCbi
ZuIdh69yhKj2j0DT/sRc31eT+0NYH7AnS5JBOcS5qbha4/a4kjzVyLApaY6y0Y7ECQDIx1zPkLVW
8/xru2a1JXnPpbElo2yo7Z9xwoR+GY3zWVuMMAUwrUlfQ1Y6+NFOPtDlAFOMf86Yzu87X0c5P8GX
1srDRZmEXKry66c8h8lXS4dH247X+TeO6nCox4C1mMUN+bjq/aJpQ4UHQrXmhXp7kwUGli9/flXd
1mF/lpHR0JUhdYGLsB8n5OgBcogDbqzZgHEbPCtLaQOf+Kqfrl0js3H5v/oA0yR5Z6Pfd+0azfPb
37QetyDASSp3ruD1uTvy9AgWJLjjmhHQLIBwbEqrtt3MZIsw+VSNSK+GxAGhTJpDAdCQ1Xx0eAbf
OzvJiwjTGLkzwEjjBolsFvTzUCHPqrxlJGONet0IFPHAH826iFHLN44TFqceYKUQjyOOT2aLnHRK
Co1hEWTAfsdYgbKkgAR13pWlc4qD9lscuSHgDGHQ63hQHgwAjVOUaeQwv3FN9RvNV1qajo9DOLlY
v4Pwf7cdaQHDQAB97EeXhIHI3OgeJEnjJ549VQ+Adx0rEI8gSME2nn8wXtttcwhPQuFO2Y7Q4y5x
31vWyz5WtZ1uTBFGBgAIAlAzwGtK0Df5QtJHIVzRj4bDY9E9Q5qVefrhLCc4mSduqruXJMEiDlXk
eoctRmH5dte8FEOcN2UrQ3Rb293fRx0McLHlTiR+SgpCZ6eqGNOizXkrvqntaVeIZTTLkT1z6c1w
46vzBXhW8vOHLMmiAItpk33dbqCz82EtM6aUhCgdgmrCmsb5THyulzLmseNrbuCqAxX3NABmaLRH
49qXHwt9eMFowdhglmfynhAEXxFWGEEhllV8G7eWGpyYYd0gR8XCqjM9Te219DhKuBnmkt26a4QS
/2P62BS+b+u53EyVPMM0n2z8LbT2rIpggI+1ZLk64NTsz/gZeB1OiPX6DHchobSLEI/qZ7pOGTDe
vX/FQfacMfdvZlVqIVaORJ4VXf296xUqu2oUP3S9Ffz1+j+7loEs/n8EYEMvJgOGAftMAf6YKQZv
Hygl8dOM9FMG5eLN7UaZXFZBusnn+pGUKIEmRWeLGB67feciLwAzBN28Q9LwwUBNw/0qVGLF0+3D
0i5TZS3fiwlFrWU7rILXHJQOBl0pxraQt/p7y4OYhjTNL7iISSnu0cABvD5ufD52qkyO0Xn/N/sH
Y4IdnpAfAxEmphjKvMEmYINqfKry+0Mng6YeCQlmTRxR8txW6EpqP+5j56QE//fxfLiQ6YqBX647
y7amIA/DHSOha94LQQcgN0aelIWQkoWztxr6NswdVyffR5dQbNEBCgARYforktwO1SiuuA7PDm+f
LDOYxbAEh6wEdenHXSEO4dAmw6vri76EbO+/4ush1Bk+nMESN+V5XsEhkhY9oi9uX1iDwc+lB8dB
9tZyPhALcmvYQIoHWZxsdMZ+AqGFH0EuQ9n8VOa1JEKYlmUJTBcv59feAJxLR21hWxRzjkcAOpJi
cEri75P8U7cNEDKGWXlb8/lyyN34Mc9XpoLYoeUnCeDjVs1Z31f8mEZi8R8n7lac5eyIXSgas1Iz
3MhEgbwGODZ3zbFxY0ev7Y88xnIGIuN9FSfSG7JJDxMliZCsNzLc9ok+oyOYpdVHoZsxeMSjG8ZZ
z3NDgNVqU1XEJHF0oy/AJBke/T9pisRH7BIiDn7f1rhjzSLH0iyA0mcOriF+dZQ+ZGrrUgYZbt0+
8Kaq/et9BXmxN1fSzirawW7MfhYsKqKvjP/tnS3xk8kvmszRGV0j7er4LB1F6+PHU89feVP5sQ3l
Bt0a1XK50j+NtJbwgkU5Dwlu192CYv6Vm0W1h9izJoEKozskyJB/G1vYsEecwPAI/vnsK4dRF03D
YN00YxdeW8DzXwTOA+VqwtxmzNHHp+u58dX+wSjt0/aAX21Jm9ZqT0Wqpc6+5zgLEt0wiR2ZZ0hQ
lPPrvte7NyTY1etbz6+NkEeL9E8hwW5RN3rO3MQY/BSDWQNbcjo7LUSfq1acLbva/LVA3LGKxeko
P0dsv7pR3Y8YgQW28jdgE3Uz6AQsrlwZtVWn7hLXIOOfsusVPylZYkpO4bW89AyAtdX8M9IyROoS
vLo+fGyrpDz2cYZItkQR9sWabE/IwfvBRDIVhNFpmv25inJgI6mWgKmj6tNM4dtY9/8aLf5ncytb
EGFUgnRtii4bgP5ksnod530cESWbPTeC7+uXqgQoMvXg8BU+1xZMwg/O0irhIVl7yz7t6oXFO4Yi
2e3NrEbvQqPe4W9vGJErkdxZuv3vfCvC0Bij7G9SMeLj/m7udB8Jeayy71bX+Iw9+mPgrD3IzoCh
34j+iCnPTmpT6V4Nodh6OaK95W2mcrIOG4UTOaai0EH1/kpPc+ge+GUO+2V1ehJc9nVhDLjlDK+H
dZ/yQ5DayIAr0qnwAMk1ikDD+Ji6zBo8G/KJZTq5zhlp8ky5s5Us1dYgYrtr2V0AGhXiKmoH87+T
08kUYUCqtAq37Y5BpvhanVLZ49MqyctKYrE7X7QTlYu4F5vsS3dSVIjSrzZaebxu95vE2Y+8apdQ
MDwTaPH0TdKYQ3L9KSBv/E2x7EKTh98MP/V1fmvfFeEPdDtXyqhKb7bLnn2VwWMYQjN7UapUjU1f
nMS/ofOyawd+oZ09gINwblRpigw5eWABE9EgEpnYinIuSNaBTS0VAL4sdC4nhe+H+4FOqJw1nsIq
m91/eeW1T7x0RkezLWYyPDY7tzugS1y0Ommv7z2mj2NvPdNg04knspA4AzxLFKIeSDWIEQJvyVx6
QDcaId9ek1fOVUQnAid6+c6vFI9tuTudfAwjxszu+jajC6g8z1uCNOyCkotqQmlww9Qr6OpHsi/v
NSF6pGiwRaFepBQjLdue24+7pRSG8URyM+AI2T6fWfjb0zn7UcLjvxREQhS1UT3eqotnzYU7GIZ8
DtByIGt8ln74UVY4U+WZf8VnUWYsITcKMnDZmVSwulaP1NvFFpKHhxy6tfcdOJxYpgATnMKF6OEf
HGp6dDIGDH/AF0RltV3wv9+CDRiB9pzhcSWHhcFG/GPXakwMPOw/L219ytA/ZCZ8ZF/c4vDWkGam
RK7eiswR2xmJPbLFkvaHWEX9k2YHJ4mSDISGYlQ+K7SiC4eQDrJ5EXh+gXweyEqwtt+n9Dp/iaF9
x8MycVF5FzhXhF/7c2DDxtkSZAac5atHTYcCAr386L5OizXyFwdGhf26/VhJczu/wUpY1UsvJzry
QbHaqSSBMAkLrkLxowXip89L/Qx3WJCr/isNqIWKW9j9cUlLZt60YB+Eq70PClWprgNLSImNvBDr
IfrIHd5QLohy01LRkotEGtCZFr57Q57Mw2lX/nULL7Nm18jEPWm1HeQWI8Gqn4mu4nJ1DvnGzDfj
vOdP8ITzmvqMFGzzMyh8whlK/yD8mbRHFsbIUCL7vmyt5Phzverum6JVqY4PM0txW7NXA0blfJ4g
H/3H9Z2de36ThUJBG7lzOWaj1TcyAT0NHY8/FXM/B5ueeO6bIgTXyLK3Ku4mNiXGsKor33kxL3Ix
szcE6Ut1CChyfFl/krY3+45flC6SmrE21+ja3UDymPzsEHlx9WMvnQ/7/UKvb9vms9ML8LSMZDLh
tGc/QDYU/a9Suf0DMu9gMVJ2cAA1IkuWvBHM8JEl+4rUGcdCmVoodZu9cj5lfykzC/nb8hDanrJq
I6+MjwqcrHPUyFqX/9O5UKkgk6PxMHrWh87FeW/7esdZbM/J2MnZhvkwbFgNfT0XSMGOD3fPvc1v
o6gkrdUJcStFjC8EovJubHSwJIrOTGPTWk/GhP/kIYmsL09PbBu67/javpeW0OktjRKk0WVGNK4f
bMbdPjIEFtFZckQz0k1wODZXMjG6PHaxIh2emjy/qFlS/3F5Qoa/43A0L/Wp1LeiGcaw5OGZX2fk
dbfUQI+kGF0c+r9zyKLPvhaAmCS3hs3a+lxOijwjTXdsYxYUBPq5BKm6m8di0Q9CF5OtjNCkwPmP
ewvqgJVNsoP2E2dcTNxeXPZ3icv6lF5ALz9xwbBVAxYZnn/25mFXKV31NXWxfKLj0j1myZ3pFxCM
UUcw5Ilx0BONOOPk51tzDHWRmA39P9j7pOJGopGH/aWleaRk36FxhkbngW5vgAJzcst5OSY9KzTL
J129tfkD9DYbtzNtCXelqJegBezbljahagbDPQVU4AajKO/6yCuhclwxpoRbVWLoX6DjLZPnWUKo
nUnXDkCy98jymufuKKKZEUypyYGPntYmPOpK5MHzdudIntRA50vVi5zkXbLwGbPLPHCdan0nBsgc
rZ08RZA9xrqfHMmsxh9+1LLaoMg5YMQpVFU4KQ8d93+Lypdv0kBYe8rphMuKJZwUJSAFe+5hYy3z
HHJZ65cvYV8489+nRSNEbcnNOSQPNH784A38r0M+whg/AIAioZfLzkj9CnL+tzHpl7YVgRMPbj43
P+oxQDhVRln7yNG2GR9n60NCV2cQYZTMsUjfx8VpYyTegW+O4bizCAXj8Swltgf9wkUQSIhTURkI
z9bPKJeMvEDHcUGKAuI86+eiWsgTnI3IUcYDqZEbuvzC5DUu2VLVGPcJQ20frqY1JVrSJkyuwD/V
35qoTsVjLml1bPs2aq+pD1Jc8ReiLS4wF/C7599Ra/6O9iU3E/Yvz2oGYJ565TbjVpq7LIacLbEt
D3TEY+8oYNkl9EjaDUb3cKjR+gY7RbMF9jO8SMoZpQ9yQTRUJyWJmka7g6RloNjS1EW6Msc3yUGU
hPKQYrZz6180WOoYdc70WpDp1q6BIjvazF6Lub0wLElLLL0pHo+aMsBGFUuGRfy0G1rBVPJFptPx
AITaPg5NZyJrXEaDqw3J7PycaDpCwV/brv7C9CiHp+x3zPRikSs/8+dyhDqHO5tKZgmGgh2jvncN
KnvT4nJ9IIZxUqdsslBnPEoNqOU+PdzpS3Yh+TAtPJdjgkQNmx/ztLZxhhsTkANAdh6y9ou/cXPR
XMz+hn9PYN3HaYtUlA0+9bUrp0j3/ldPNkBTMkkHVmKgDx7O1Nv6zEsGFn15lCy2q1PkECz32YHL
ZbAj9E9m0ODSqiEkb7x+e8is40KLzAHL4Hp3ZBnDHUq4Mdo7xyoOHgmW2od9byg/zIQ9KdodE7nR
/syxYGFk4zqueV5Jgg+gasDBmsvgoCnyNRiiDmSY8ok68lNoN2WNJt4X27j7yj8v7YakSI3QrT9O
fyWFP6Otz4Xh5cmHIGaQaDB8v4xWjy9Ytnsav227ETCqSWylw/i3KixyFHN7BqRjKlB1sKnb0j/+
h2L85OgCJ+vPP/lZ/t8chgfHdGULB/ZRFSDJvJMkIQb2qq5PpAlA6qiv8zPHPaUQaFcbntCY39Io
2PGJmnSFDBOyXlOog/5nT7BuyJ8MQqNXvPJ017QHtp8ccpHVlktgW3aTnCyuKEvMOZrqtLnupQ5f
eei8t0Pvv30k8arjTxyzd+dVKJ1Efvqa2uPhvXOGv70SURUBt9uizwctxplPMptP8aw9jKU0pj0q
lkw1kO0iHRHx1hH1VKFesxuNhcuI1FYGPqjWMeMF1gk2kYLnaihftAzp7MMIraAU87qEzGxFXtL4
H6P6Nm0VHzF1K/sAsI3jSsdbOAlr86ZenxvBNjUb8oQPC6TNad7Fv2NqciqJWmgaBQ2AlKGsWLGF
A3TioRCfAp8F2YYkJmvRpXADiD45O1tbqe9SOdrML+6gye01783Ilw5Zi8DRv67iT62Wvd2pvUU6
NcxVSQcbC4sBz1zDWzjTOrrdMtWNknRSqNNYguzj7CbaT6tAQaLJcHTf4oZJlXVdIYXrTvG2Cwme
t5eS6PMjssqbKOhOq92mX/4kIAEn7pTZul6NzgC19pI5wkjQ3gIKBDWrr9eUF4tZlNFaqDko7ipj
sBzV4O2CkUdk/zgDBx5hIXW5Z17Nltv+oTQox/954/3dvOzkPkhiLBxTOSxnzwp86xUBUNYMI9mS
OuCYu2t1KkPGLuQOfPtROGm75AMAhsh0yQf1qy4PTJW+YUeRgx52/AXQqurqWLSmB5utVrL7nBNw
rfN9TyLR6FiaqBsgiQ5PSIXS93plXkheqGfWUIi/Qo2tYdwANB18lgxmb0rzeRAHH6WdmEVZ/bDT
nrdgPKLMlES2vd0xcceN0Sh8Un1L1840snSsijPZcflv4vME5tduSm3NT8+wpIwuef6XmdmV1SGl
oSa9K2/3E1dHRsYQk7PJ+0pucRBX4SC59xLrc8yDe73iIgeH452xAVAkQKrwjd4LjyVwBvf7WpYn
Sa+zTclutvyNX+2ueWTAhwJ1+GtoLMHv4iG8Clb+mY+VmlGV01Hx5XHOU+9gonLYVBU4yZ4dICeo
WI8gdfwjCfFYQk+cQB9bgarGIrmvxVcqCyZJ7VP+sTfSZbca2z4hfZhJS2/HIwo4CWVLL6KilSzI
os0szTpQ3to4LnSb9hnPKb2WTTHXkRKVVWP+8To8TaYy1bX3AEsh8BfC5jLMU63JjQSDYDHpx62d
+sEXlQzVrZ1SjEznXEOMt+v7SAr8nOHnkDCRBBIaAE5g/yLhkzu4QKlr0XaTPrhIt5S4c7Ob0OUJ
Zu/ne/ZjZOxzMRyvekbMCnHLoyyDDFyMLMaQIYPhIyqxmb5qxtZrsQFka+X2U1abbhxwvutnLxJL
OIZ1u/srHEwtCk4fBJ6qfGcsHK6WvZeRvK0DBZEPLSagFTZGznkkQfPcpTn3HeZqwD3jvUyvChmp
odie7I8l/UcZ12SnMuZ01DjIYYfK70EjwjhEV/pg2Hz3+gPFvCjZAU61PQ/tJvHJsWo7L1YNceK4
ujju65SyoXr+WYuxGNJZgA07ro3FQLHuuVcbo5R6xnxbaQEMwKbTjrJL25BbK70jTDHzKjHxd2xK
ns9RMgtUSzn3+h6FPIcOA21VHoJnwGvj29C6x/0l8QgkVZucepyEIG5yB6vMFVAX9fVrj9zneIsO
PWGWd6FbS0lYvsbixhJlhvGbGs8aBhR6uNMGzwIM26zKnJz0ln4eUpb/0H0Mkw4l4PP68HjE4eDz
VDonwgwcpaCcVMeBAxfwJaz3vp+3iseTyTRgJe5vAQxSk3NIp+fiIZdH7lXaxsTLWUoknAagJq3B
QBvaRLxDGXs10CS5TXIYgh/MfKU8ndJuR61M+aK4W55njyVIoADuoEA+FwgUhTS/TXqe+l2bjqVi
Qa3tEIf4bLnGFw4kKS88z53aUK4Xbm9At8PwFGgMB26uBswJVsBGHGEox2cGirzwDlejdNvqF5y7
MqwhcId2U8wqpJk62W4+3drZo+8X3r+RUUXxuOFsuCx+Uij0y+eMoCSLTcLPmgJC5szeTEUSKL2G
5p8jNBC50ulzIoOBsZtz/xsXRGiWW2wTpzfBcCVaYZ333JJftkzJ/vR+CWBPYkrBfV4sJypQB3tH
ErWJb/UC7kdm3wlYZ6dZuTf+OZjUuGmnsfM9tfqurFkvIyW/vXbgLNocdEsmCTQm+QZvvwkU05en
BOCPB27f98tWbA9ZvBrr0TfEeEmA+Je67mggMdA53H8UdVULG0fITFdd741r7/md28ZLjmQb9/8R
KW09pQcB283bV4fTt1nCOhNEEAqYGgfvN8fZ45hzredrg41GKEmCYWFdjh2QT+XkSTRGmSyPLUEp
rTEokKidp/gyOCg91C1BnAjHuZ73RdhiH0WOcgDjecSk2zdczykBiMkuQHQX52E8HhWsaLl04o8B
ckxCA8QF3v4ppWMYvNljURr4tMfXv7jctEo9XpQXJml37OMy+6FNlpc6yU0zZc61C03PuGmcattM
TIIj+spaI453mPRC5fioykPrBVH2ndh8LaFtgevvVTKGIFO7FM+J76jnfIBANSG9EAbZz84n0Ymn
esXoCp5U4ogkYliZUlXpU/+5evTPaC1zUKko1PVVO5VCYLoSATYvHGZzHGWlPO4xBYwgGqdgJ13Y
anN7iIoN9RWITopU6chGG0a2damwbonnZOTa09j+ch/dmaShgiftwu7u0MXXEZjHShLH3dDpVi7W
zGG37BGy12Sr3ZPK4GluL94UyqGaaYTPcbCoDvHyn31tmt2OoeMlRT739VqRPc1MjjXVegBYMtjs
EpdpwGo8xTa2mf/9/pEO/E4p7LZAIM5g18Jq3RR35HXyrBcLbNHG4gB4/cbXC4DQGq6daunZM9zV
nbothDqk7kwAJwMft57u5/jQCnsLePcqujOr0C7suVzRVJ8zHUnAvKaBbjQY0NTcqaMY43gZZH7g
eeSHi0xbTorZtD1gD3lqYWwK3bwBrGl6PnnWfQbWKyvXTOWYVyS5dGng9kox+L8JlLEMFKjkxap7
Iw2Af3mZ7r9c5GSjT8xBANzA8nYvyn+52e73cRGDI23IOU0KFjJ82ruD0qiJPIMCdL06qC5NtII7
oSUppfPjt1NGvewZPUnj/pEcI5AFs/Qi9tVQ1G0Ak6NMek4WLfSl7AtaPfudPqKcc0EJq33zspxu
PRbfzD15DkTpXCl5ZG6PKMkzOSRT2Ea42JG7+mRn7ZA2wYjdrJToIqFCEzpuSUWXPknDtt/OTmiT
4yalFVUaKwidNWhVoKIwA6YqVp43OzrQcjryg+/KrCRfib/5YICS1iPH4LHcsBXwCRuD5jvcx1Us
aRi19AG0JpSuVKhiFublcuKWHMVXE3Q0rndDxBjdC2/ISvnQrmTNHUin3dLkDyVVu0giFjkFFK1u
jeJzRxB/tJBKt1myWhwohKGQOZ2rsFK7d/iQDfDV9OMIn6qTPdTXYsLNRAXhEiUlQqZIXQRVJaUn
lYwfNACRy0iUPBN9kMru2egq/6bsD36zNvMuO8+Hrx4IinMM+5wnBtJ8mt3YIM37uWgEcKMrZ/So
P1nPlkxztNw11kTjWzrpkioB8BVegN4J69n95p7RuvGFFbKVKFRWK87NggbukKtsTecb9FIRlRTq
BkEsYREVrfUEnaC2dFH3GGmSEi8G5CSGulMPbmw1gtqDgDOsLLcJ79ynCKsHLP0ofUBCrIspB5AU
4ll77Hxi89wbMNpm7H+xx9uzjMklviKqU5gZA+Ao/TSHKOIstBbrB9YuUTQncuaFF+qneFBB27hR
ZXULvDK3pl3x/yaeyeal6ZWJZdb9rh+6GL+KCuDddjQqHk9lTlsN6aAX7D8h82MGaF0+WIRiugIw
yAmxQ7t7w6YGGSD9oqdgnPCtEvmODGRyP28EqMcRnxlVVAoY7m6FyrMr56j5D9kyoZ19TAdqbUcS
TphcnOstmyRDEC2pccELkWqQc1IDz+tlTLOsHG2KolepxKnKttrm3uB055GbQCqyxg6/2K40y2C/
aqFdtC1jJ2R2C14K53ykF5VSFInBAmn4vrzcGHlf1NBOhLgnmNTb497q0ZKmUR87MO20GBWXOPhj
O8M2n3/5l3gCYzSet3R9yspf1OaCT9JCKYWA2iX6JgabcbIRTwWDtOB9qkKgEebK4JYuNnZHbL9+
eREUQmrvqXiLo6ECW+BWybBbJz1H49EvjUjJ4620X8Xs03i6QuFb/tM5YhPats+ZMLV6D5ty9FTW
diupBlomlHn/hw/50Wroz+803Fzj5jsmGpjrynr0yZqYL2KUPjgrAGByAlJ7bwZG+0FjuVAb/4z0
7fLOIqeNOt9rfqFVKYFPGZOdMb/fmUAdTjIkxR1cviKfqnSCfDGPMLuwuOa/45RYQo5NSNtFQ/j0
P6KLvjg22HAt6SDf6euUDjFHQJqioEt/iYP/KsvQOfU/YDTclo3ddBU6k7GXAioWzVBM1vh0t2AJ
GXPkmR0HvtyLxX0HqpSqgUcBQOTbJhVimujJCZ/dVf78xWSsbkHkmelTXBGlbk8y5dRdLsCfD76C
/qh+5LOKQEIXj9LzpE2t7Q4UOU5lJJ/krSbUMpzMrdxpQaVrnGD55f6HZJmW1r7/HcCu+FMSRCBn
BalOUDA309IDhsbYiSv7QJwsTsyAPIPxmHAcL3DP2Q81HL4EA5Xjp1xJmOTsM/CHLlWVzYONIT1H
79nswwYkWDMCHrQOt51k2TTOTNK+7ooHUDluOqfN/Z/Hv/1KQuJ2yfLzQ87Eu3NGrvBV0/5l75FP
J5HUBa7JYdCjXERisJlKbGzk47J68+0MlsZz7EGZ90cMRcZQ1LWlKMYFrvbuiKBhJEx/u8mQYVlZ
EbNvRJjFRDK8qL5Ts7ZVZLL4adN1Ll8C6SR1ffJ5aiMAoUkW/SoRJLKSFSGr/GS8DdVhmq2pisfg
9ZPtJPTlrlw7PMnPtzlABLX3ZyBDXEiaOmaocWSSoEwcUAc7AJZHwgKmXE5SJK7TeZ+Q3pryFQwX
AZjXvgPu1Vn7PUQyGtd/XprVv/AlqhZg7S+cELiG8OlmrrUgI7EseipU8alMpsXTb1letdMS8NT7
OCV0zZLNkPjstzUqnhCOMYh+dUDXTBWJYvtTekpRvNKxGz9T72xZ67QuMpEnd5b92/A0Di9EBAlS
AIS4RNn+3T4hGUDdeVTQ0+Dcn/esa294Ys2dAE8dMQI4FlQUfOxlI/J5+yW0EEeds8Rmo6wLBEoT
G7yzB7heOtheH3N6Twa2RbWi0lpkjjWmVZN9uZCRQVjbFYhMZjrs/FEg605yIIqAevbBV2JaQBkd
Y0kkVZJCm0RCGRDapgGdKTzbrpbqkmWs51A4f3kXeGoGQqBzB4kpUIbgI5vNdLQobuGngLkyhiVW
lS+b4yPW1hZnqwhOhuzUQ+S2kuQ3GxUi4jOB5/N06/nC4FLMnctPpKJZZHIiZwcV5phaMJ5l3uTp
HKWBiqVmG1c0gK+YAX/N9/cSiDIYAVCjwRqKzobGkIo1H2E6aWsR8OMzl02mwIPZQAjIlWDitryh
mthyi9BbU6SganGOCFoRKdY8S96STM+T0+S8D3vGerQpkIAza6TGWc0+nljka9xDRvbxuZdD6/nz
SgA2Yscl97RAdDBtHeJYYEIb4S+hpHvuBGVs8VhCeJuu/J/fxO5CTQoEfajWeA+aWJdp+knM293H
I9OoFtcxs1FNkp4V33/kyfQi4Y+B30K7CQSF0U/5g9+Q5IHmR+J16EzDAzByFd7+qBXQYvAdUwzg
DIxB5PvR0iCfg0bVbhs/zWL1JZ5gGw2/tt+wq9S52Ky+W3+j9fguMF5FLDslyFZuEP9ka7GDiQH9
lmxceIQ1cKQbKWOFbGQ6wrOzrQXWOTPEV505yktlX0IXmjg94t/ebUKj5ZVZU7V2lmjxnXfb3Qep
5cCVqO7pHTnx5EXfXO+YhPrjSB5Ygoo+rUEJN6cFamOUkr39AEhKhQ7Q1vdIvaavsuT5iasdUrXX
J7gibOia5bexrjp5CBD46TS7OfjDGKqtHKrotq4RQmJCX15B1biorxgAvy9fK1rimzyLtjU/Z14h
S0JfUjtK8CCXZOG4lVOT7OUKpyNkVh9yXJgGyMdweECNx5MO6xvAZDPUhdKZS2s02i4JLpNb6dSw
Bn580qbSJml+A09ZVlMpQwVF1BtSWbZBuUo3DuznLTTBIO4TLWficr6BSDdx7zCj/bdX2DSQN8I6
gijiCgnSOqponprGzOKemQc8TZMHP9/ekKqtOOKfmHQy9jJ27i/hSrwY8rSWtNNZE8Dr4xLd0MW+
hPwfNzgZt9ua8GUXj5P7sbvliWRSA6FFS8qPB/+RrIuPQrIl7pg8ff6jli57GsS3u8ZtRnGFR7oz
DJiZom9T1nhD/wR3FIaw3YWfaOPnXK/RzmqGzJYfpjJ6u1BQJBTfAT6paVnN1NQgrddX96dX8tC6
Z2oORWSysx8fzKmOBIZRMi2XMsXJ7+EIj95zxUlf8rNUcr09Nb08CYoFOOevWhKEC7Ejiod2bCYV
PjO8XS6wp/DtnL0VV5w5Zk02FjqoIXqAlE1q8rNGeUtBntpyQWnPkDAh8CCH3sBVvcw0oAgaxIqM
c//9VtZbjya5EFfN5NLDLFYXUdk9FGcfOai7M0VAfi3OuuLWhNcPJ1rx5QOee3grjxZayFkIP1Kg
8CLRiYxvXqpvlWGBOtyLOG+frMxYPFAeBPL6LApfIq/mBvZNAimkjjhLjPeAmSibS2FW/av+m/Lz
Ly3+l56lfPtYQtSSVGcH6rqmy8+j0GX491tPme7aet2EC+sqK92ErsPE/16HqswXhNa1DuOmqcKD
z3xwV5mJzanwkWIGKsS8eNfFBqi9ztRMZ7xIN3fnFtclC83XKFA2MP+Qlyu/R589C95j/NeaQePO
ztsRY+FrtxD0eaqxNRgoxNsPBicnHQgaHLlMqByRCqm6pAgiguQdP3Z9Sv3N3l2Uo71SVmXINeOs
Htj6EgCWdV5MYMzq5cA+Rqizj2LZKvARWOZek8p0rwRPjpJgVqZ2pw9tYdp7UsP3qru4aUbJhQix
ooGR/xkLthTf+p1mxCoSL/xNRhX/q53mDr4ZKtrZO7BrsPWo2FBLnhe7ou0OmNWfwUZWmFX9omL8
+8ba6Ze43xWR130zgZ3GQyvXNtPxk+W/b34BdcXHXKZLUVL4GVVhvCgb0PXdbIznx1SlG6PXhKQy
7aeh5MR846+XYBWf4WZqI/sRbfchoT3HK7E+YpAuLRy364b6tHByB9DDYBv2nADO0j5Ro4LyjWZG
BgFzALb9OkxHsu4TRTi7ULdatOccw0PopaoWeyP1XDBpQXaktBb6OF55F1bm/kb18uJgiyzvphUR
zLA0OeGKddMrPTVniNbBI2gozAgkmHRd85Q74A/AjAJeYCnR2LZNOA8oLpIR+Y5M5beggH3foMtX
0tfpYeY9xF1kJoxb4AjjY+mKCGDG0aqIZe6b6imHYoNd/YeehZEi+car6k/MCmVkoCr0stTDp1OV
7Q/IHGHvQfFmQZE6eLF5gJ7Yv50hF4hl4tD2UBUQM9/riL7t6q+Gwqe1XMLDs7Ix4MjJtPr5S/V/
M81RiLSasFacDvI8e1gaFNNjqVDP9xUmC5Hw2sugLYRfZZIFMbwc46mzi/UrM4VOKMr8KJ7gS/pV
ZmcgEox8fARaz2qGqY0ZFIsd5lMP+0TfWTg1N1MP3s7T9WkZDEDT/mtmEkOy/BX+nLcBkXOoDsNe
nC47UhAvAJiD7ofwGddDOukpq3iL+C6pCgACrbwHwRokcH95HgX1olinbQ1izKPkTm9W8ITPnpFR
wkz7+X87h2Q6WqhxLaE1WfhOMhd2jrKK9hqcWjczkb6guAXeNynvkswGw+x8/fioVIrEufYB7cpR
Lzyoikt8leTek6UqpEXVwurCRRgirjAePMhjUG0oL97ORI8LjuLti83OpGStA7t+asZGvng7YBwf
Fou4q5FmRsVQlPHk6yylPs/+yeOsmvAlbhJ3/8TBZf/qr3hXMfik+QJnBuGgXWqqafkI7h3XdG7o
MRttiGekA1EwFO/ARGfqN73pNZAbomAVINsh1KgjGyu84xxDQ6h/uMuEuSSCVXALrlQhfLipGcos
/usYaYCkzzVZ7KbdHymkcwLkA/eeMD/y0u9iFyZ3KgDzKf4tMsZA5gKYj99cxcotHV5Ri8czXNiP
twgnKk/V9CajQqfD5uUu1cvIShudYzD17iVVZE1sh3LSnVBmLmFhmSckbMoVDIVyjklfuggi1mLu
BcMlfYFPLSOdwT3NiK8PAds00nljy7rw5qoyOH130hn2LNlaUZUbxqPWz8HUqiUQUShEW/BEAy3k
tFItyQ5XhRq2BN991KghnJfti/AmfwZnnjjGQLeIef5FLGLy9Adq5Z/rbD4/oKVOlD8EPDmYP1tD
DQvtZVu3nuOOBbNFL/MT1Whox3AtA8iPnP/5Szy19+f0Jt5GBjadjjt2OY9Ojv/TflnDNN7pPYmp
2a2tw5ljrwd2zgZPcL0gUEEOGD/rAAi08UcRD5aqxK57QUColXQTzUmEOE+GnS2XRx52jm9xMxje
IdPTy5Vc4vcu6NqIFsP0gHqto9UEDktN7wsaY62Xb2Z5VSKeGhaZU2RKTZAIk0tR3GcL/PS2CdZP
qvo+Ji9BprAEBn98WLtyuI/8ke5e0hdErhVVKE7Fqe316k2wJKiJlZdVnENYaxCIureLmUcWYddv
h6JRksxTWP400H4Kp8CsKBzuEIFzaBoz7LTi1UbDYpPSFY5y9atH/ibKDZlUYTtoS3qzfI4mR8sZ
DKkGWZwU/ocwuaNLFWFRoqA8/gcPDyTuaENy/1At6M/Mw3gJP9W7zG+rEmoBc/1kH0atHGEoeIfl
lGuqU8CUI1N6dlCAC2kAHvszMOvSg0yIwdGuobDagAq3qjMaGA3wLqn8IwCEKB4SsdwNtnRpolN4
3D8QDGCpqwLgDXQJkojBNvUGRYei8+oYeP9AUoDDuNRZsNCfSBsbzziFNi5Mh1L2P9adqXL98tA8
flu5v/mVDOYC5sJ+M4x9HcaggM8CKMLCBBagB5qdmkjCBviVwrzVjezRFno2M+mz82vKcYFwT+sU
nKBbVXVayQLaJ5h7JYJgKt/jir/cGuW3w1Xu0qHeX5wejsB6Aa8RYK8gt+9sRZy1rEaw/Tfpz4iQ
USbit+ImDMY2aFeS36ItaPk1jLJW5uTRBp61AITHLE/Ed/A2YPO/bcdcib1IxIXcqdCj7XgPgjl5
ruV+BTJLpL1EgvmSVdaVJQvBXkXFBQrA8EWHA8daKur+ewQvYxEExMiceja+i7+N/GJTKPqV0t58
TQy2JQOtUCWuB5ST9MEU9CqNcF1YQUWCMgrvTY/Rs3CWxBUtncDmSCFFc+Y/i+zsOrtKRs+ju+44
sq9ZzBhK4QHsjSShDUte8oWZlkcfFYVUY6JOlsYq5HyE2kO9m3vKsWEkmVsBeiVU/m2wBsePJp9T
wRIkyCrbwPGNzGVpnBQbZCyjjAM6N1fvHzlJNJZMI2ruP//hp/RLJFLIiUm2mXKGD/2prGbLncFz
ln/I3cMVgkA1FoEdMG+lZooP3y4I+xpXZAxKNaH1I4wnEzhi2a2B7hVCvE9PXFnrYloWpa8bQzF2
KnN5zXXR5sL14G6Q5tYYc0QsyGq1ossWI3uJAs0s9/sbuNWy+rlhl9gQuVgYEHyLU6V+fIyQEqje
Dj1ajd77rdwfovxdb/FBont5n5J26h/Nfhfd2bf457gFU4W3/8ZZaIr33XT9QtWFN65xi46dk0zQ
UN6utASCraQNt4Gn5QVSJxAH1aD/7mlwpL/+D5OBHxAyHriYk2KsZs2UST/39OBinxR0fN/FOY8H
rndO7GzToY+FvTmkYctr5qW9CAHKBFMBYCu2S8FtXtC/MdCVWyhACP4UC0W8R1xqr+LyzMwa2QS/
reRtLJuo1PU/DXzTrJ5kEwzbdpfCo1PBS/yqMNLRfZ5Jvy8IvgokWs3STDPpD1EyS6X+DSyYA2E5
VRblDGUBKQwhArr+sXfeTYsXTSmji/fzuUf2izC6K8QQ86/N/S7hRy10mmu2pHyRSUVjXCkWlkE+
HZihCmXZB/ofDQoCtRwWpOxdk/sEUxs+u2Mx7Izz69ky4uTPyl9U+QlMyjwKyJ8ZWaFdFgYXmxas
gfmwp9Kt3ZFeMBHHBaXyFZVoj1qzri9EJeN6/cA7h1mPv+LwrVRg5Swkkb9gyCkl9Nh9ICIomU7R
ypJ513FgAVJ2zqqtfp4WAUvTjhlWTQgalwRJErYUJs1aOthJ5lqM4xVC7rlnGuvqRNLIiKh3FjwX
mpxfoaFwNmMQj4fSekR2f4SSjJjCWcyLcSWrvoRKmuItWQxXQXDKsUMlZpTHreL6b3OR55T73A1r
E0rlxHDNvg3BhPj4ZS304rOkgYedz8Cx6q9CWSjArsOKaRDrmY9xXAyXjzfwuBCtI7on/gpI6Vms
5vdW+Ga2d5UQ7ZSqZTm7q4T1k5RaVkDa5hc2VfjyST37efyrNVnYEgo2PTv/CraFp/hH3Wx7UQ65
7fCKjTGUWJIR4GvgpjJ+TCcjNA1mJ5nrsI9t34VwtBlHKJpa+RcAqZ2bw/SVl+yNe45jAz+4pMeC
mmcfy/+udgQjsSfhW/RynoO+qPpCXxt0EktHjbjBbx0+OD9FYUhBV0dpNxkQ4a9vQzKwyWOiegaX
6ylmKGL9b6o+NMA2BlmVmbWqlcLi5qmtf7t5AVTsYPD8IK4nJaYyfkOZcwoz0YmQAOrFjOpVR3Id
rkIy2Sbe3FR/8B1ZBLVQgrSCWkv4DsJFaroaOy4JQUJs2MX8Mycuz50VJY3As+t+ehIpd2XyV1f9
+RYylZchUyJRAhmuT5HfJQBTxD2GvzrmKDq1k/lg36/fepF99dNjNSCsi3R06TWoE12Jcq6nSAgu
ugK9zz1U2k13lnPL356JqlBl7hWb6BlhsBfe72ep1t57lVVkYCPcv+hCHeyDqGS/+kfp47STeWMJ
uS7Kmvytb/b/sUF0pOqyHtH1oYFxTGFjeOo+yLExhMw/sUbBfhZXIvtCXL0Ku2cfObegK93uRZ9B
gZB8Fkx+SvlyWgwUF3nVBFSeRnMq26CBQ/R0pGnFb//X/3BLARCqkYeaeuppmANy+mCweSvm5Wxq
Wh1AjLSPdE368VmZI1r0c8L31oMiSpiAKaaRawkQljd9QXUp2H+wsNXDkU7rUtEyhHoyfs0sIsPP
hOYpnRH31UkmWgV4fuW9GyjvoNbodr5U+8egSKKZWgEQFOPfaTcdrMCT4Caey3HGO2THGhlCqhVg
TLw9cMOP4uTK2sAQ2wwN/Aci485+Kuzh66QYlcnNZIlOJwiG63aIRwOHXfs/Xk0BMIKakZwkRRR0
EiUltQ6SCZHUedj3C7s+atqU55DQBMADaNSyksCNj5iXYvN2KR95JbSJHl/iOFQknvPr4sfVQq76
bYdzhZysAsrbXhgkAzxp1hTnkMyZhVgs4hQQ7E/RkXXJ8+FuOFBEGG1jMC4AuUiUyh43mx9L7+Xf
Y9YkdrfUfEwhhP5kHop4qrioq3ZuMwz6K9BwrSgiFSDBC3FmhLdEG+iQ95SqKox77wXCJBg5VyKJ
TDyzZgzaM/YNdYa0zWq4goZau+uq+zNbrfLJ4DVbZNxb7KxspHhAXi6I7sdJrQbw/eyT/5xvT2yf
ay+h2d1GdEwlrkaocV2z8NrX7JB/enoVqypYG5AL3IuU58ZsYKh+2GsEiy27ctP3x+8Ol7MzINXg
q3z6l9CME5q4P8iFYtiubO2XO525hyTZpV/hoYDPgf0sHoogEkJlrxA8hAh4Z9dLOIfQw8Zj3kaX
giO4Nxi2wSa3Cxi/WZvdLEcUuFaibdgRY+uK14AL+geTaOhNRjEU7sfZo9D6TcpHD12IK9R5Jppe
sWZ9m953SI5/2QzhU0mtt1qijtC5I/29esnMes2OE/I66bjTRKDVdbYO0apmF01AP+srHnkHhVny
74uz5554okdQbXhZuIdirD73bBXV50WbnxVOO5+CRH/sQtNCThPR1OWyT81N/9aEKaoiVoaTrePS
RJxn7UD5/3K9qw6cxIyTIPvqbvwwhFY65Ps9EaWONFH2et3pb3u9Ep20VHQabog/a6N7RGybvhyD
dSiATiKJt63jgODLN5sXkdVr5LHbqGL+Q9zSApRoqJCyvKEPolPaW8dOgNDEdBRV/VmgKLYHJs36
IvUDf1OpHq5OBs9G54jdZaHj3+WaRgt4kToaUZzAgCfoX0RqT9RoCNRUl35rS2N9EV8Kf4wCxGkD
IHg4E3Mg1azY0+KFiJk34RGSidM+HZ8fufVsUTedqph3zKBYFgG9xmOIHH8GJMINo4yUTWRL/LSx
lN5sHw213jsnFC2mR3HqwUWWKd6gBCJydEhZRQtRTcEEAlYAWGhqn3t1fbwnK/n/qd1ezMqspivp
cCrygWBSCNkoB9+nLn4fjVDJV4OEOAlGH36f+76VvhAZ2/jy9jV6gtJ7+yXSmXiGtmk6/99NWBXs
db501f7dXWgFN41blCo5u0ir/9OXyqsZaRnzP919c2r4DYraBnQQCCBH6lRaMCXFaAecq8aN+pzy
umJWc+gPNEEtbPi8eQhhb5Bt9D7qPGYDE5Hy2DCYdKOf+/HONEkcChO0cGq6HrXdyTfy0gZNPIiM
0NKMjlxd/LuB6c9AVlQl7MOaY35p73lAQPXqUloDPh67x5N3NAIIoGEztzkFcXWt6iG+uQkHdkuM
6vNEjps9DoHfGQi0Jlb3sYPnvdQTA01LB5xLocZIhdRhxhY/YMjfoTttVh8tjJUj0NseShanGJSm
XNO+AHvMa0kvhoFRsyqKXD03W1vuli+1y+oabh0XK12JiBJCDpWFXpQNAaP/9vmButVsvKo6lfz0
QRp69belH/ehnZAgAEiFUrsB7cc7hapqGZ/+Qt5tXeWJeptLjStclSaSG8+hfVMM60SukMv3yxec
Kx2ZeTPvT1g+z6WGAvJpVmqq6nCQXykqjLYkUfR7y9dfL4aC3ZpxQGo1adBqEU9uiRMchwWwbxAG
SnxqHWodUGgyV4adgKOGXZRvK+jNlens1WK+Sa/Bp9tk1bNzdqvGCCKxy/qiiMvX/Wo6rb+Nv6s4
Hjg/kCN8jSufE17IP1+1DVP63PN13wfDCAsM5VW2RBxeHs9Ho5AxBPiFxvP+XjyORRUEgLoLe/Rz
IFtwU/NWc/wC1yEXJ8hYvX+u06eDQFOMNlVMBBSfNKGjIURsxoyTDPYJJ0kBaSvx+fJiLCZZNnBL
efD3zSu7UG24BHXovl1vFNWdGTIcpYI24VgXvoL8tW9BoYCj+IIiGZQRt4EuMHNakh+yH52nGgnE
a9PaP8+TFBHDhNTQOYWIIAffCGsKEY70eb0ZTwa6dIVxGgpigDZv+dEz611kc7zT/vvF2jH/jS1E
l7nCQFvzk4VBddkJgX9gqPT7ZyTUEdc6WUJnD++xJxnoNhQLe8wdBev9idjs2mALNVmUMg3OsYbt
2E/1QiJI/yEMtrdVEMUzjrJ5K38J60/cqWm+qAtt3SMxfXVwxHSoMz6XPyY1q0p7GYTZQKXwHGB/
M2TWuzeGOEWHmKUdJzIIHsjkY2OEZ2m4tm6quQo033pwBddAhwo8bUtdySp920SwewsWFvkVhkTB
1HotMvi52jsn2+wsFEY/qF8lW/fgc/2We985Np1a23Ijw9Qg4q8PYjHbSgru+IyatYbFoRtcs82x
+Z344+iX9uyLUbMxxhGTXutIjnfh52W9hCg7yLaXZ19mcZkZ3vazqEgmZw1OiRSLl0x2kxu+Z4ym
C21lEEHzBcJVPD3OGrDcAZvR3qmDDD1MvaJqTHzc0VY0iyqITZhMw7u3++rVd7GEMJQ5Xm6zB/uY
UmZcR9HVkw+/LJoFVnNt3Gs5EhJyyGKiiwbO47rGvVbMqe1SMWF9vQQtJ/ca4vgxB04MHtu3Nz1+
ksWki2UdAzJTg1+rDNl3MpOzp2eCJ7phyBTIelEFVDqCoC3e1IE+x0THS0KcG+ZpE9veblWqX4YY
R++aJr9ujLmpzp8So5C8ZnFlfQoV5ZXiZxJxlBdLrOf9baStHIiPOra356E6yBaxioFVlZVXWkqM
vvqVdg3V58TTHzZGvM0XajxU493YVpAlCU663wKhmkmaxOVZ5HEKRbgMiBTu0vwyQb8KUC0iKyT6
zHwoFrFsnUwLlVuVprFlWBy0DUaH2MqBuc8Vp6uwxGFWiD+PHQbZ9l1Dc1lhyOJ4VVDq0b5BohkH
H1EjINCRF0vhM98cV03AzLctYfgpdJARL2uV5gTYC0/7BrFSvH+Dei1inuXh+4UeOTev21e6D6/c
RO5LN6g0t3AlJBiDkFuf5iQP5eKkv4J1YUACPk26PDz0jcZq6tIaDubM2mf/rjlpQpRDH7ewF6e5
/jZkhu8HklrYC5MWVBpoZ6S3KIXrpAjeVZn3+NU9pcylRlwlJTSQYf6981oW4GJ9P/GXzjZWjeDO
OPEzJWK8mS/uONPqC7aLWfC9C4hhFtSn/IN+7NWzsMkel3JfhvBFIEdKnlIAa6WNLZtPOKvsSPad
ok4Cuu40jOvF/xV+oDOd/6ppOml9H0oHik+km2SWUhVwIvAfXC73XIHfn2FnFsTZOBTj/E8u4JfS
kPeY2pxVdrNCngd8mSu5EKZXFqvJiZOuQYsKn2RjheHnmo0qoWURiPDK1PKg0qiWuzfNInCcO48s
z9CUQeyqWZC5iL0kF0y5uhakZhN++Y7cWaMjHaveLZpo/N6FAR4ghiSBy0SePhzspW1YwYzSfaSY
1Q+xJvsEQWyRNUpWJUg+RO1Wl14JbnerWELjd/eo4HHNTv/p8Ka4YUCO1/8HjORLJi0V7ctEZQ1U
iwLAxbrqeUqAjNiFVQ38yZ6/QN4TwWnKyRwbhsNww3pJHEF4OkOnTyMqy9smAUeKJRJVcaZaWspJ
kp+r7DVhkT/HYVnTCOZdQPF+J/piG1DHd/WDiIpxgV3Au7g1fzSEZlAVlhNWZUvNZYMg8NFUV7KJ
W1+LIKGuuZTLZp5xzR50P/MQyi+ddjFyNrV442LzFSRXq/39WAuwMyS8TOgS+4yFX5ICnmx9BT9r
j76rz3p5CappM4ZStxB8nkdJNYONQzq2UWhGi7bL4/OCCqszAPtcTmQSjarX3TyND4YXQquKT55/
7HfxItcAZ4GZoX2LPcQq+HFR0WDrUJmJxP72j66ecetfHRXoJhOY4p7/6qZ6WlPzHQ3ugYLudDF4
FmOEqV3xUOtnJqACKDh09BKw1gO9rrVR7ZGbOtpuvQGvfp++ztUEqaEvle3f0zaMWsZj5hLQNweM
X3BU5mAjyNJzZDihWUvdF9GOqgXkpyHSNq/8nq44W9N33JICU2UKazh9S8VT6308usXzl9c2buc1
dn957ZYCjmVlz4QHB9obubfzD3CEd4tVc2651Hk5lmsZQofPYm5MjWsgY+vOD89sWATKCDYzoywN
F9xk/779+P59CGfVl/u1NPnLnsA0iLowLwV8gdh8OiePUML5S2Tl6lAtev1XCqLv6IyFZndkteNi
sZnhlGsgdrsF6RaeSslo0QpHEvAzLJHVCJrm5wEb3+nL2Pvsp+F4Q99xUxlIJJNTjUoBinhHpUfF
N7X1T3PlyP9nEW7ZmVKwE0M5mfe9TsI8f9D7CbWcK1ip7o+5zYsYNGFWkcRjBL7rYsBIeWVPLYUn
Wcmfy1mxhgAiqPvp02IEHpO/gU53foaiCSju/M+jsHFQHsv77dL1uSIcQlP5jmkIqUnhP1wZ6ego
v2z4Mm2A3ks+wq8J9HhDhs3iq7wJyDJDBnk/qNcjmpBql/LzXC+Ft/XYtKtK3fwgwtdmcLlO9kKI
qbap0Aa1Vn48BP361hZZU0X6EzLqku9May6lqBR5rFnxfPLBMFf3AoegPMSdTIk8ymd+AKAYXr4f
bCMJUWcfx+6i536zDMasdJ1lXKXNXL/yacpvVjirg1yQhnhNOmMbACIREsVsAzMfwtjG+BogSy65
Y0AeVSPeV1aAJW5N5E2XDDNx8ZN5BH1jN1pZKfCAL+nBCSp7wgGCacE9ZZJumaVrfKV97MVkt6bV
xjTw1UVXmho68WZ47DQ5AIKySglK5ZVds+UG2Qn+crqVHp80ETxhTGzUWMdxiNdNXlZsEOYCdIX9
XRA2Y3krrNpWVsygaHaqxMwWP3U/blV0t8yoZAxxmnieJ1CGCdMB8I28A9GCDSumVou4rV8OlxYx
3Nnnqn3TX96JA7UP72oVcZ1JHcLy9ghl9ybtzlACFXfcHgC3xqckXVgHje+rcHvQ2OJmz5FJtiFQ
P2N0x/L71oRQ9QyJUROYyeuaCoG1DOOaZCMprIDlau74j+pLVTwXFmwhoJ6oXwIbcQHxhXTj7xOb
hHxsF0L/newseDJaD3pahwZ+sSejIQC4HfaOh4YMh5H5eqNDH+1UGuXetKCckpZtrsK+rkLRn/jx
vPFCx9gMljjlUiz43Dam1GFHUXYyacF0TxSG0YbDOOc2yLgyR5nQsPj1DBvtfOmTcBZPTys2RYWV
13ZdsMx+N6vLgTPyIdKMn1sjK0VTL+lEKEnAMQD/qESe0dFpjfeHFoLHvUdTWR24RyI6u4nA2J8W
qVPFA92l8eM+XlMdKcHYozjdTkRO0Cg+B3BIB8++19DBEMFEFKqopHsutrvzS/rt8OgK1+V/BuG4
oDMnEJiXHBEheCcqNY3nwLfDCI5MjbDu/PIOhACpmepaYtv54nPgqkDuqKxNAA09c7XICAiPH9kl
osotB7eidU0SqBXpb3YoeCLN+EcxxpW6xFxr3MhtOQxX1gxBlG/enxLtXN9VuCLjDgQcG5QbmTaN
wnyz0m0hNmdBp+wJOA0FHeuX1PqrSMibvsTMWRFdpT+VXU6avPiAMWdgHV3kVAlPaTq4xPEMyHr+
GcW83IWlDb8H3Dr0dK64TenHNXXgAC2q473PTp+L3Hnj6VnU1sdhIZHzm1JS0iKMdwTUh2DR6fkv
ljyXtswSWK4Il6R1c012HTBrhCiqZn4zmE6yXTjGD+Uekw3XSfubfLFg7vUsqKdcGsgOFUegdjOz
aXmelvv0q8oVlfZmzY1uWu/m4t5fAOgEn2Pahw3m/GmaVrWcDpBRGBRkdEHzXEzwtRxeYlXsWltk
iVfzTHTgBobUm20kAzkDbw/LbsrXxOaekzsV5lJl5EBl8v2vMs5pCC9pC/0Q2JJ/rydtX8rWEmRi
RFy7dz7dzXTe0GQx3pYDnCVaYB1Xh35eE7BUo9a0VnPSr7a/HtFKX2A6ZDKZZdtmxPBhWYchOQUK
AlwmJlyTOPbV3JUwNte+ZCyhmWON9oNyEiqG3JNrL1x8wy0XKXP331dUN2VfoyMUB5YfRUwwUZyI
Adobxc319PhZ/45NzV3KOAzbAm5WwdD80TiRUFnynQzqOD37gtKSkKGRO3WXMAdhqA3o3Va1uyK4
JcYT9glEpNQge4N0gDa8KF+KC0gZy+Qv+nHYnqHDRxB8RcdzdMMO5sTHSVeT5fjTNnZpcOo4rB1F
MxMtL3s1EjU7tcwS9yF+yK8M6ySAZMtYIs8C+6r9bjq7yDpP4HLbI3Cf3HbM3Zc5GrQXP0mcTDLH
E2P1/zNNW2aUOzNhMeFtl14KZqgSbz7XFtdnkEzQnLii1ia55E2jelQbeobp+ZaWUpBEQHmow87Q
KDtQSYFbyMde1BtIJhLl2pSEcsZIzQ4wgzc1HJi53mZwzHcNPpEPcj7lWCsfoaO+pYgblBGYFsGq
grUyv3EqE9rPFrYd17/0TrU6wbOhDT3DtSCd0qYxGHKwRcwlqIL4matGeb9we5mNZLueCQsxWx6n
Zy288DGlhRKG++nrLkznrYwaz3dFz9S1Y0+k/xzXlD4TINo2n9zxlaTmEe2Eyw+Q2hyLuCs+g+0D
A6Sm7+5p54otE2qOt6eLFs/qAli1767oRExCWEK//lQUPfvT/WyzpcG5ATjiQDERyp3mtG5Mfphb
RafZg8RADBeKYAffOZPnmkmQN/cuOnzOqhEX7VBIF0TKWdh1cZBxqxMeqNmAY75qB74XXWOMqalc
ZjkdaIOEwAHhCcwvtB1sJwgy/jRsomDIK87IvKpQuH1CSxIBh9Lp6SGPCwU5ZK1wQyfxGJkkuk+0
2PldSsgq7kcSTv7DZDcuJYTOfaJIYuijeYP95URyB97gREX57YyhGAk/ifsn+cFkzK5yzveJ18HX
WGvJYrheEWSQRQwqwWTniM0K3Olsx9h753QO+MvpMcx9dHdGuDzmcoLQCuOZaqL5DdpYx0BuM9mr
VLpsd4plFKL0oISyCsltUpQui++Uwy7aseSLxdDEMTz2judxnvM2587ronIvm6xsUjc7yrnypZwr
aLXu820WeUxJZpONAEXCkxzuEhiG0lcesuUkHTCrUQkbOjCr175AWBEeKcnOgrHLwxUAzOvqr0sA
L0cc8qXO0JrV0P8XtiOJqDRUb7BzreieVS4B4/e13PkGr2ojOB9O3iJubuYuJIGEGX/MbAwDoaAr
ne2oOWwYLffXStj+lPRITSeTMakQ6AMh4l86lcH71SU5peLn1CFZFLzXyQxk0dxcAwoP0/F0Ua+0
BohfXUiSwLmvCFHO8N+Zs4pjmfEPACVcmmYDhqBn6fpNG85bsNUPmSnQjHJDj0ZaB5LErkDELM86
1JeLYX7PVmrdAmmM3JRegZayb5Ck4Dl8QqcqMAnKIDUMfMAyEl8HFPcMgZ04//FfIwr/Yo5o8MiX
ZW8ZVRpauVNYPiDd11FVSMqT3ib2nNPb62YkSlGsPfNPONb/N9sRNo6pYi8Y2+BKonbBEmanp9/O
TeS59mDNaygxUOzbymD+X3M+MK0E1kwxqChOsaH6GRppb6e/13hERGHbU675YMOXBEentgyKlwzm
DOsu+mz95lGn3/4kcxL6pD6wGmVFJbpmI2Hn9PQqqtBfOc/vQKga2nlLTaSYYSq96TQXfhOAIKUw
GSof8HZPCGIOzkaTlCoa5oH+1CfUapvXWK1z11W4CqM+8Kl2U4ndM77+BXeNy5oSN25UiLzX2aqV
wtl3pAJB6nuRKmHckCVXwBdGl0XoU+y16noJnLmVPw2Lf8nFHaJ7UfpLdtczzYA4IdnA5v49CkJW
aj96d+jZx085R2ApueOB1E/sFUf04UJaKhr4hQLftOeT4Pxsmowarh/4KzTu5UChpVOzMCD77cvS
FYczx4zkYp5xiwzH363GECDom3Fyp7lQ6+4ILWnWn+EY/vjxcCDdunu2HgTo32p9InQR9zdEHjBs
TU94lAsXnLX+bCpfbqS/IbBG3zNoITwgJ74sHqJyxFjUrpV7tsaLnF6S5PXdqTxApoDi5g3nZg+d
cJDm6GNzYIAYZPi8K9Q8i22RxJmsJzWCtlxohBIfZd5875T6xpgmNirMspqdfuJtyCFfWHkoJ+nk
nJ7vy95vQABwjmtLsqx+DDzlRKUtqbKyDypd2tjoKUmDmibjJMM3SbT9QIG4oqAsgk8a9KrG6mJ3
Z5qVN2kOnlrp73XLq2+j92/8AblTh4Xkt2G+Q4Msq3eHTOcy69Bvy0YPfIIbj+andTywcWn6GyPH
7WkYZ8Kt52kFxzcGWGspIEja2mNGgh7XrLnscm1IpW8QLRebcpJzV4oSqbqRGt/LAoR1Mmvm6irc
V0hcWMst2IvANwUBhqPFkDYvOGPu6qAINf/GitCmHEgwsPBYbufpDcPYwKi9QugnQMh3Vk2vW+6i
p6vRo8IgXRhxknov21YRZ2IaziAdRtIIMCnsKTyDKSikdYpdoIpk/MIDC4j2nHLfnW2fn6ogi6Nf
KPMsiAFs/qeEnt1934q3YHzVhn+Q9gZkYWxGXMxlMFYrZ1+uhGdRFFTIYxLpd4HXw0CvhCw1B2/Y
bbXe2Acmogp+p2wYh2qWLM3n6mtbCSG7XmgUVVKs1Yp+21TfRQXFcDNwJVkdttc+rhOZPWhDZKKU
e69ryyNgqfutBsJAMu+0Ieeo1tX8M7Ly2bv1K+IMvLW9UtbKFqH6EFt3PJTJYLBKmqtpWVY2g5eL
1Fh2KGUNZ7SyObieV+JOqBQjd01q93fn0DpqMphzwbl+wmZSQD5EjIR1bH6MoBYRQtgYdOOtUPng
3NnvKqfb8COsXWE0nx//Vt+ajoldoiqHLhszTwu89DELvheGq9lKGJASGJ7lk0ABuhsCi3tTOvVr
I3CQsZjRoe4F5J6P8c439Gn00JabTFP/jxYN7PMLwYVhhrUcVMK6llbtSkSl+sLEsILioEmjLnC3
eeMmBgOR/O2b/t8cLuTejdlSsxI21JFCN+Ta+JBlQF2vIiB1UbOSnEexH5GxrGB3bcAZi3clXPKD
JU1p8q41WGunAAcAPI8gRZLrDNLyecgOn+NdVncqKPz4rDBRwNkoNAZEpjyMKnovqycfftQsPs5V
nli1Y1pmMKFUz/4IIZKYs1iLO49lrjNKM5e6CknwyFFq7lv1/NNuBrxOvZUwxoeI17kUYIQS7dMh
Ps9eNLQ6FGm+HXlcXjBbSh+xcnzJpvGbvyG9qauSNs64V7TH04ifdYXyXxZTsEL5mzhtSzZ0LJeC
lM3nIm4KS7Jsk2a+gPtR7qh3ifpHRuNBzJCpjB7wFRGiRxLPai9uwI/L/Za+F/z9UwVL51pUekPk
7rM74ptuK3BwkTD4u0WaAbLafszx6GvZHj1F0O3jiMDliBe74iLKJ2bXyEQCzc12QqC2ELe73v3N
XIBF3nFmvZPXmJYmRGsnZhN55Z6fIVQQ2z9Kx3k8GJY+UhELLwn90ejJcV2B5tUWthwXWOhLqGDb
cu5AvnfkDvYHEpYp9a6haDy/mVptALZQd76Hk4gsttlVHEmxMafBAb/hmvM9RLLX8CzamtSWSgzk
mbE2gx0jATC5pRGatEIzdadkerh0PjC0hsl7tUe1vpIlu7CcmLfV9V2UtyBhHy8DLH/BxrokTla6
2YmgUSiKZJ/MamUyCnFFiGMKO0IaJbE1V6bzt71mkLleYcrJQqdkSJg52nCx3ca7HSVdpV2AHafT
SrfQeeFsOBD5z9EppNyrwkM4ZvDiW8A4CPQ16K50VsuelqsGAVlcERIY1BbXdIvJPi2m/PSbuV4c
h9H/EjR7/7NvSlEr68AWQe1TmnXmfSbuaTby5x7bWgz/7GEdl6RPWsqgEjmhsJmOrNU9IviEcwoI
+izb9euQGm3JlaD+7rm2SZ0atytjyEsrLoxcBBVyucLucb7LPINboAHZZcuWKUCIb6586mbp/HZ6
EU16LLAnbZPUspiBWuDiTTHkIK3zYQwnuOu+Kix0728T/nkCv6J8Pz5nqeY2uoiyndIOFSRV8Lzy
5WX4OPm7pjCrx4WRYJLzLcfQjZJJZKwK0sJYyY/ZRWWbi8GLl8WxzK1PcWcwGcTIAXQsu16g/2zo
7SqxtHk8BzeNbJFW1au9FfV4SAe7J4a54jlybcK8Y1dThoY6sSpt2apUqRFUGvCtQigqfJiKpg6G
MFb/AbmDIbaUZ8w5vBLZ/u1KgGyKY9Egf4EZNjvNdnb8d1c+laTrT1en81jbb9I1KzTsHu30yM9L
nyENYxopVccFBHkkZSofWmM0Og3r7AwsbyHjXDhtXKJHOW3N5Vjgvz5K2onvmCB+gIgiTp1eCXyx
IFVWa083ql/1INnvqi8qzykjSHqs711i2vyRCAqS7WF3/tXmvK0WliwvYFhqUaiRdYb4X/ZwrRT1
gHTB+b1x8gPG6HnV24JGYnqHKLvD7YhqPvYgURW8dFtQ6VCDc7bXkJifezzP6bf3Pc2I0soV35g/
TIss9fOqyt1J2XDFtuxH7iCIrCgulZ3tOTcbuhm1lrriNm0nw6ukkdror+M2cRC1JeKIGHCkc2QI
mUhoKihWkN3uf21VyJx0vbxV+DNEnbyKbIHNwo/1fDdtoXbF5FNIjR+4Imw//z5BvAHzhnbZ0Zl/
0366Xoqg8C2vXOE1Z1nn9ytdNWIjhuXZ3Pibbzw8/MbKt6/us+sLia6OHMQOXdDGDbq2LdgZoa3O
ZZoHVnuvqik2MaDcSIoj5+C0vEPopQuXvgGUasVzHgpQC3Q3nS9AXHvLoNEpLYf0ILeE8/XzeGh4
bjlyHbAyxv6dfhBfQT05hnkZ6cCNuHxUzngK6+RPBkpRxtxvVmLf9ujdg6IvyXPeXIaORPqUkrf2
xR0nLkFsxdPN/ZQkn/UymOyob7q2lfcuqclMgdXUZvJY/6bZ2EyKpjjnYUBTQRY0eeas7+IbrCL1
BlYb2XKOoHNhYo53PQ5YYco6A74DpN/Ih+uN7rFoqJYRs+Iqg1YScV1aRlm4ERoBbINL057t/lY9
6jEspUi3PSCy/KLOFgSVAN5zJFba4RrKuoeqGqarc5q3qPizmLznY405s3oC9vnMLyxfd4hwRnV2
AXEULuU3MKphTjhrQUUwTQiJQlMBNWiXEiaTj+1P53OBKqQS1QbC8m3+KChk4Fs8RKJWhuLhEi+L
WudJRAu0Qrj4xuHj3h1jinl0nhV7LJhiLXWuLXTsQNvW0a0UoIkmtHr9abZ3rotcIF2gKl9ff/Yd
XRsJ7mTau1BYH9ldOd56TgfD+GHCTwcsaEQYnP+WowmlzYsFUqiydtuPdLRxPIip44VrXBDQvDZY
rCqmpRnd2MlCCMLSPjxz6+oBQXLxUEgtZRry7uA/poMi5RlbrNrcWcPmasai8m4l8UviO4rTMDpA
CMZzLhRfwrvcXrMu9xAgvBB6VhVfu+9GeJ70ObnF3A2GUC/fy4FttvY56ltJ/8unbk+uOEFtA8A8
WDTRlg77BSFxC23yLDNkYY6o7lILJUXMZI6FChtA8qWhPt3OMsvL0D2Fa+GAJ/pt982bIkrMg8b1
3PpsgnWf2OleuxGDaMW/G/fYy8j/k19lb1oR9+MmfG6KCFq4k36Hxx3RSoPFnhutYzt3U/jYsUmc
Vn9WVd/08Xq3Xn1rMnX7cDQhhoxh6wky+JfN8IXVaqu7DFvMHHu7zYHsE6sidp6rt0ApUsHE2qB/
ccmZqh80vj+HSQmYxQ1JZevcSHiPQTFEfOWnJOnNHy6n1yRaxVToIAq8qe/d8CVHNqysEETG9BaL
gZxP4SfXBPaRbvlNxbjXBMMuriuANx0Yt2TB8nxRrhILdnCSnmFB+2Se3N7R/zJa/ZsK2WHvqwph
9/dL9oTcWU1JIE9WoaPucbo3JHaTaCUzlBHnJXLlc0NqUeSAcKdM7gxCGZsedOjPr5SSdVu+Olwj
pb5gGOUoVkItqHw/cRyXKKQWARojPcfrBK64m8+9I5414FfWfQoWeFjqs3eyNf3+kc7U+Bxt92a2
LTyYbc7pDPEIOa39EMrXLgjfGoL6Iog0iK14YywpM3j1SXNTFTSANIndimLWvnG6VpyWm+L3mYMx
e4fnCQ7314hDTheSiWA3GR/R+JewjfNJTqy3gFK41cueO4GygYtZXueKcAyRfjm942LpgkEBYIOC
8/oHBsJuI++6N1Do4ewyz6RCWClmOLbf/A5Pj3yWTtnE2VVGEg3+1v6YTHYVAn607cX9lvmiZliO
F2R7NxITSqgmrNKeCFGxSe6HDQVnpLAwsINLof7JwDRbcky1O9bpDSxGnbQ2n5y5Ko8kEF01szTH
ZuqQYuxkHrYGKcH5Ad8DMC3cIsdJVwyUtP46ueOTeNrDYYOkuGM6+cJkOseIsaY14kEtHgYHmtQv
dUzE7ZOSVpKfGe7s3pe85U4cYV7Mi4KY8gnMMzeGzBAelVByqSuWH2wX1KIlWOIyBMhi/Ll4M0y6
vbSvaRbvfIroS+NRBIQgJ2frWWPsjStU0FNRbqNmGznw7Arb55GNVMlp+rrYnDw2wk/f4EWY79Kd
AdVkLjxAsLXR4/+vxG8Nez/aHKeIVicONgL60SFV3UA56WMql/bKT8a6rNFp317FP0dKXmEAl5ww
KL0M2M+qlOlsW0wnZ8tRZoQfLCOgtkrIbaHTAMJE4gGrnDG+ER80Q2ntSRg6XEzYh/yA/8H+j6YE
WkckADaBYH6epX3ohJBeLs+nSTuJ1ftJbkCiYDkQTeV/CiLgfvgW/E0BcJRrjKVGBQtDsh1NExav
ucsYS+yu6AaNOQHgX7VkbbxUTHEgH2hLLF4+zS9OpUGtlhcoirDqple9crC9YozGjoFk4Ac49ivR
C1yc83WPypqAhFq1GUxoq+0V8FCPTMXF7jBaNE6Hi22gRTmL2JENTAtaxb2nHQLING98JJ3o+Rq1
lSShDdqGE30jascfqahIRmDzvpVYvSxDDfRl5xixQT6bCzJ0uxjyaEB/U04ZxzZVip7oimjeHe0l
xOX0ba2mtkD/p3uXKuLCjlwLadRIpYO42GNI2StK2Dn6Bz9rAvpmDv5R1/qrq6SUo6U8Er/d5SBe
KrGcx51KN0AmPhsyPe4aJTumR8dVV6efFlfYzbmb6sQ+o+jpKrCvSRYNLh6PplSMx0je0KTt5wYf
WRDZPECrFt59eqYvv9ChhJ6809JeRCMD3c3Z4Y6A0w5qxat7GoXGvRCnlVbpvkEkCEizqV3sf7Er
XfVeEyGKN0VryvocNRC7aylfG7aifU/BAkYT/0t8+bjpeXctcv+hIdo2SdjXNyyyVAoPGRSo1ta0
dZSw/iWlVughZmdxCcdnJReulE5Zo+S7R7khau3A90frekEqMq8E/Q3pROLhdNFbOVLiuTjcI1eX
KQRoUicFt4eoFxS4xjc9dPY551H7uiy5Gc17aZE+C/iHewUcpRLlq9EfsXteo3o1x+1jQLlky6Jt
cwZxUodF2tYNhoAe2okztUtbwRHeTdPX3lzE52YDNK1LjvzGwnUZD1KYu9yIw8zWFBCV3owRtkZ9
8SAg1Q8ft39RTDJxWRi92YYFQMyG7b0agbwDesmWv4vMVuqgDVZo1rwQz/kcFw2kBg56yimwC96q
JRyy/TprDKLaKGf4o/fHYh6zLlmcqitVykZqLhEV9iJjnUdLl1AKa6WyEY4l4358EP6BF0DBnkzc
A5Pi+GRHvrwj0RD4Iuxfu/oMURoC9zxYAwNjYh3GxpuJ+A43g4qvwB2tzPoZJqSehhtsYQsviAbd
eZugb/fihyt0VwbPGi7xqp5hD0eqanCj0n7gQAiVPcfbOqD8x9qekZQ789PMoxZS3PqYta0Sx/SF
qImeEjaTOi8SgX1W9KXQ7m5Hz5J9xl/0yP+WopA4Qz8oywEB5RNEL3e/gUrcwlPi0aoOQ4WK1Mi0
j6ovptq8MNqSfvJlh+90sxRakS78rCWOBzE9DVnx7HS9kQwkYcgxt+Ca+UllvpScT00c2fiaHUMm
V9VAaeBmpaT6P5DIHdAgBGI2wyfmQoCut0Se1PQB69zoXvc0MbCmqe8S4mzASSBKzUgocA9a7YNc
7Mmf4bpAHNlg1axRZh+bSqqJw9BP3PxS/raO2RyOf8dBKJhjVOZyRGDHCskRdNE+s5xER5ux6dg1
CP7M/nUlkKsvoz0akoIMRFHMQ2vIQlOVt1Kn5/OHpBlXYh3rnDggi+YzEY6vMMjX5Fs4+4asFvZA
eDywxqUP8WU2kqwJ+FYEaozksZzndGJR/kT76ohwEVQztRmuE1at0uGrLtW+uXPRWdSFieeFNRjI
NjFBe4k0o6Cid8KUmQRu7UKQUE1i37zuLbqtlkFAimrHT8zFHCL8G0GcFgZ065quRzGg/jxP1RNp
t1LOL1kHPe7AIR7NCO1mDcQpIbSlf7agld6u6Sr0zKM2c3G7dETpBoJZSuYyGUPutP8d9LXCPS1I
foadpkO5VBxKP/eA+3C7koYX50gRwE6q7BhkAbvggO9R064WA1FQ6f0wg0lQRPWG+Do3ISQmtWjU
Cqet4yXpnrGVihl16gZZHbDPbzIoV1pWtEIzNqn0MaLxnU913s9cwEJuZqobWCJHN/do792D+El+
jwjsfO543iWtjfJFLu5DBw2Qip+Jbs4EZimZhNWSKSqdpzaEFLB4PkL1kEHn2SqL5lPijJA1GiX8
gnkqm6/9eN7VWOqwqh967TWG06CVnKpYlk4nskglrd329WEXPzRkLhndt3hzkZ+d9mIc9qHwZ8AI
ThYgmZD8aRlNXy3QFxn3naTdHb3wg8/poP3vuFYTrAJfJYfo5wcTgDTKpXZgYVfZGsrWkjbLza7E
xHHXhAmbHD6Z09MlCkozYKKAQt65NhaUNGvzZJsdugzYxUL7hu50HUofVdfV2djlddDaBChS8GVU
NXXARMOK/hz8ZH+Fb0KgVINFZjQ/+70D8WuFbXU8djCMoi29ATC38HXAt1R75QrDtT43ae5bSRi3
lwa52pCoZ5W9FxpBYuytewaJ89MIbdqmDLe/keeQa037unmK7ATKZZTIrdNVkaWDV2yNzcYnHdcy
UQeSlxQIGuVbSXhYWi2dpXyZiinJkn+FwZ9OteGC0KGkK0zZ0oehoWQ4wcbnsL82OT4WUue+gao2
g3Srpwqh97Jtim4JwxyTWQ0J8V8wQWw4os1qwfHgvCbJP0UEEFOKccor0JzNZ+BVsKHSiw6POhgh
SSGBnGSqspVRxQt9arMPaKQi4jMMepzj6V99+FBeIgOxGjXMb1RJRVWUEkigI3HkwbPgYM6bC9Ar
9nehu0vKtdAPwibjaT/ZgVowIMkTgGdM/8dpSk61bx8Hwkqihx+F/RTlFb5emAqeawN4o/AJpFkM
lJAxgqjFJ+j7vOx9i0jbl/2Ql5qlZAHdovGuKhTLVVjT5/o7l2qd1I+mgxaT4J8LY9kPWD7tzDgf
rYaqFyXJmEJtLMVLWzFIwgExonWruyFBoOxEcfhRy97UOyiANsb/RoaKH/fFDqp9QkcL8UU7dG8f
tPlUMo98pPi6yPGuU/NJ4C1dTRsZ2kYmxZ9Ma8fiit673xqtR4xjx/4+FXvI6qSrOG/l4Cf1OHlT
gZGuzfU3HoEblgKZ/JJBhe1TTVjNxGFwDG8Po2FJS9KrJIN28O9HQjXcnLcNvSSlWNy7pTcQW7CR
p35hXf1BWC5GQ8WjBbTgR+yeWuePqjvZvqtLU/piMFBHG6+ARFuhaCYNLa0/snnpFEt2WH04oxSX
uTchhZLa2alIogq1dxTKUsXU9OuPm2cQT1XUNWPbiGouxSLFrPJD7OiHHkpFz9tYAXInHvip+VOL
j3tZfN++YvqkS2mf2jjOrHm2WookS4zmzHwKQj+NILjpFx1bNBeF4JlKgKj4EGAWIi5CPBZoFOSU
yBDR6k/LRMnNCd22KqFJOwhfco2fMg2n6yBF5BSAsZQIcSQ6PZCFA+xR3yy3PIWgzsGSMrRirnD3
5KcPm/+e/5mS1zWMSBwpKOA+kHYdYcuDfGwIDBVvUt5LCeQaM1gwz8hXKTrQ2FyaAr1FBDCEdR1C
1kLPCMADo0Oa89f3/mkfn19G150TD4u5HDgIopl6vhvkGufbJM2jA54hWiSnU1EseCniiAnyHZmP
ksnc0eMCl62gSDZhoYQp6WGuCQ0GUxGDnAdWCqCp4RXfKHr0Es5vDUMDZYzbdKckcGIgjc3IFsPL
vZYnCCQgZ45mRKVE3cCTm4Vaz8Jq5R+kDp+WyGUxdlivG0DlRwckBECERB80KDvnQPpXuoU6pf3T
SAkeyfzWTmd2Hb6ikYyQfw8qT55z+GR+TPImFTbv1O5yE6nadBfxMjWtZ5F1A0sQWs95vefNttkA
5CsljFCVquzi6vfacpNT4vf3xpoy5us/bVERHzFawpgeaLxHsKXmJAL3/b9K7GJN5P6Tn8aKJMGC
Ji3V1xUx/tfiqzsUw8O09AX7+K00W4nisa0PBPaHMJ62q2Bba5QDIjSFupffqUGxU1qLSUAuk9IQ
66idn4eZsaEf5xt34P7jFswDkewlam8c4iu/UZLb/nV+geIsDFkMJYF+cwGZ61+FDBKU3rvuGFKe
/JTAR6ttfGUUZ88l3/TLu51dQpW5TtRPSQcLZQ0TmdVVWUWCNvq5JgfzMtsfeZBINyhkljYrKT1c
7UTWISMIIO6I6ajj18rTCxcqIihRNSX+xfzcXDep5PIkqGXfO9WHEyRiArNX5m4jGGnJqRa+z2Vt
la4bEfSQMLbeDtVAVnhEUjly3AVotfXiHPfl2F9uMPuwf/K1NGbZTDdmlszt/A22RP7lWfFBs6T3
ZRGlo+gxxrUuUe8L/PJevh9GN0alEA0WfcdDV8v2k9YoaWxcgKyVR5xnQkAr+VTgMJWZplc5FyX7
TlLD1228Wf7U04m/aEcqAGXHDK9yxdjIXtq4xUqfYGx493xrGRtZg/Y3Gj+I1k9LRS1DuOj8420X
zOkcyaVOUe0VAzANtpPorMmGpFy7D5jBMvx+pwhbWvq1BROIWI+nHGbg8vDpJjlRv6YKXBpyM9UW
FDMyzBD2a3KBxLAz3DjKxs0gLWNIj7QXbiS6nK/xUjB372K8xZ2/D4kgZrAklyv0ERFgMp1y8dOg
8GO2BnnaZcQRRj8GFM44G5QyphqV/UFKZvJjvSMyA6GiSaD0/hrZTgoNfFaai65O24F16+/zetMk
HQRYM+4EvLqPc0oQxtv2aI1OvL+hRa4MOheqjOR/z7K7rg1I5jqieuGlQq8Zxv9Ts00VzRjqrxbX
1lbmYJ9mEWHHWj7IW1LI0Ghy7bfxE6K7RE63LsE4/TtW8lckZxtgJ5pXkhGvAhDoukjYGPELpZBw
FH3fvZb3VNEmKrV2pnp/kV3B5SHk7arD0y5ZBT7xzog4RThN0ftMbzZYsTPLq4oz65/1nlBLesW5
C2cCtODM/hRbuESGhvO0fGuDKAuIN7H3NgUtWzSXaFtl7qiHJgyxM8m07pG2GZzJYqVrpkcv13pK
dDom6VxgFRollQ7+O/tt7QI/JuzxK27Fmoxs450kmyRPMf/ZG2gDYL4jn/vgUnJ1K3PPJznp6tJn
7C/xwo3adEZ9nlFcInZzucYZPW0fAzeKmDZyJlmoF8S1B5r0weQKO4wCwgGwtexPXffvsh6HDBiN
XPApUzx+m885gStaSZTMWOyKYbotEpi5pGyEL/UW56KvHGsx3KSMq+AwdgsO7D5o1sioB+g7uH3O
6Xx4a3X6ADCHal9+qmYxLslKqx3nyPIs4vdL2txrKm6h+6KJzUqYtu2TBURgNYQ1jcsqre4Iiu9j
8sTRLbQLTK2xdaZTMH0uxG1BqqRax0Gl7DVd4kmQN5CpQIqekCTIY3aG8piNqsA11D1ui52jjRIW
kQ3l1cC/y2LbziIE1HnvAhWs/FyxkfDT/in65S2aH5aQMPlpER4nOHsHTxCj93AGxMit19IE5nkB
rVY6muMGb+2D104omsHfk329NHEPVDfmQmosYnzANiM9KhrNsjXlqfMZNidJ7hTXlwp8lHSxAFtf
fliP0R3BoO4TJIy7Pc4b58JAJXTpYkYwq6V2Zy4AY/v2w7GxQavHJTSYmYBEsBHUtBoF9egOYLJR
DkdBtOXGb4sgaFADF/cKjFX0VqWIVVeM9lSIQ4VR8vDMRpiOKSQXJHtNmH+A9N6R91zkB9g0G9Fe
2qNMxa1FgY7xivmNTzmK9eTbp0KqkLIdCMSmXLOsizCy4uaonzF90bUO4BXLnv8SvGDNGUrBhJtO
iTKuyuh0EZkzSOO/lX8dHNEKP1opwOkViQ1nWmx2DF//ZjqhlqP71XLWkb0JSsp5PvtQr4tu6VJL
SoFI8s1JleCrCJp2764shTlnUQri6LNYRqqviGvnRi1blGvRSIU4I9B0gmQIDNHR1QxR6Jfcf7zz
5aCKYdYqroKFZqtL973PrE80ca7DV7Lct1oStNFgU21oOoy4A62squT/RFgo86PiWgEh0UnFdIeT
9DS1kdcJgXrV9Ms+M9Uxlk+/tQrpznrXRgkXIjg2MhUnz1X/9ElMfkjTc+aRFI9Dy4MRr1q4ygoC
ypHQWFzTCEUgBK47gE/YbIweJCNXJJ4Am6XYWMksOqTHvUJgLrWYnnpGIXZNj27ShYMN3lyIGpTk
yzIf+avgKD/xbg4n6OfkFeltXMIGkURGFQuK04KkH/Xl1+9VC+/+HFo7rypwqspC9SE4uMP10d2A
MRqLIzqPdj6WzjWATmG7/78Rt9pcT/Fh7b6lB7hChyl6XBn0/eeGZFIStm39VygjVg3GMY+gro54
/+QoV1wEnEViLrtycMDZlzQX6j3O0ZYx1dHbW0MSqE8JEY0IGF6CR7/kfdWDNSUG979PSctlDOc6
nECVk3XX9Gu5pxZC7cBe8SRKhEM1HThJg5s5hcjAKcPT8ml5KhbrIyWbhzJ7M890uMBYYNWIT1MR
RCg/V5BGLlD5JWnAfh7e7NoLwzhAy11rw1yJ3523RRmtvvX2XEra8qTY7vb777caaKE1HmgK/OMP
QE33XuassOmxjg1DP6wHEFcK62btAmirZm0s5G5Hqrhtej3FALA5NaOOA6J2gxRbsdwQAKMDtYv4
xoDaNyigP2ly+/hNxTwez0CSDghnrSmbqqbs92zlJwaQM7xhhrkbkoaPNi9g08/2xKBDNmDZDkXu
YML5dE9wPeF14ST1tPXGVIFLCmXWljM4sNMQtKhYeFmbiy0wQaVGYJPNY+mxhC12H6R6j/FLB5Ch
CiG/y7hEBCMO/1DI00wLzmD705KZU1e5JoDktSrQ6xKkRXBWBz+EddtXY9aioyKUuwvWED3D3N7x
H5RNnoPd8wzAnHy1G9DXd6gGLAHCEfHFkFclT6EVxBOaIL9KBQio4WfqTpdT/6D3yQr/LP777I0u
VtiEwqLQ0m0ilGbqXEPIFMv9Y6xYF0DK1uEe9oNLEOwF7bzOmSIzMPGdwoRwpaTPA89QyF5R5S3q
9OhAsETxnMjhgiKmhQHVTgQP5ILItIcKLA/jZWbzuNuONXlLqjRoajrJrk+XIyU3QC1/uiMcTbhd
Q/3a18C+N7FY5aL6xrYTUmnP8fNXakIPdNG30Dnh076+Jerm/hwQxOG5aHyGewzgrK1AQZuRGEGB
TAvkrMfqHayHkhAnsxOyq2mj9MUJwelEFJ6h/FculNgRVFJCNDHx8nqt1QV8r0x/2U3Yy3vPZUk4
VP8SNoFibkEhZrvtdC60Xx1Q4R801UlZ7nLNoe0Brjjg89Yy4iUUo8stF06VlPoK/q+8wUABqbl+
hYEBT0gZe6cTDx3c2YULULrb1vdHa3edfmDhGpO/Qa3+O3wM46XyPaTesjXv5hr/lbcdPVAGtOOT
E9zLWSq6p235eFZ0olRAWhc0oz/9CT4NYA939BBw1pqL8Zc79Izu3vkzQgGqqIKQXOc0tkhP5N1N
rLGhncp5T3LYWH39QI7iMlODfAUWexM6Nb10gx51P08fRF52ARtcAUh15wbhRwaAXdyJVbkEHFIW
4di0DPa79VM0C8rXiah5lHrTT7RFEevgOA4mqL8+8SDYycjTbbUfRFlMTJRWjqh+eGgYjYAAdztT
qJYYUrGmT1CDxNnB2j74l2iMNNsQXw8v4fEV/Vmm2XGMPt6TacqrxY9iYVRy4hr5Q9VQSe2s9b3u
W9ybUr0/Hor7iATot/0TZPYVY7IjvErjjmHbxa9YWsZkVtUC30nMhuoBOkkhcNdg6uOOD9MhEe3o
jWt2YlNubgNHBYp6w1e8NYPBK6Ub7xO+0a2qfRMfzSFNFJmNFwgr7S1f1StBvUSXqY8xoGaNAISL
ICQtqpz1QOykIEXlOdio0kErZQNFYaFaUlsxRpGyiiHmv1G72vN5cnyG8B4qO0Xnw6fjMTesb9zK
yrUWApGIcHEjn6TroEb4lTwXN+2q2jmCuhQKRWKLoHVEpsruyHfJkt7eI3U428pZqv3I7KP6svWd
EGB2HMvDEknJ6kiL9BwPBQnld6Mcvij8ZKULrQZrvNfUcZbUz/cLWMxX1ACEUUbOT7as+dBTa7Yb
RPHw6swMYc27pxHKhnET+rdgbcU9LD9AN7xf78KGvt0aYHEmxmwXFLaFYT1UHMSOeltZ59FW+vzn
W5O5dpTON5jeQ+B81WbUYar4PY2m12KiNbrFhDzUF+eLx25dglEtHxKuX7nDajSrHGkFmLBy4cx4
OY3EVPCfMHNqcfbKRzizeDdu2nRCIVmkeEObqWvpz0R1AD2ftF/tYTR0aPAlDrNAMgyGLuMtn/fz
SgmuxdCXN2smFCzvQbGjbHVbJkCua3RNcr2naX9xNNrpa2yOi8yL+wDSwHMQwpE9f+khQ6F5+/LH
vDfnDFeNnE3dAjtS/m7u5TrLlw7ISqXjvZbmbgO8+NpEwCwycyV0WrFmOmEfH3AyMvF1e11evlM3
kLElQZYWGRPIx1zkDcCVZUbqV9DZvp/IZQqi1Da8djEGWHOJI5u6EZGP/0CtBe8PcrOPuq4n3pw0
5ZN3LBiJg1EPWQLd/7UTgVb+PXk+PJNmWe/Emxj2Yb8okYzoUrCBwMZxNx+6joXlUelfIOeDfQ1B
HZI/RClVGI/3rpw6IwuKzCawzGqMv2oxdS7A1KGbGgfksPTLmgZ08kdBgWlGfDZ1IItcKNhjuzDf
pDDwbnHHccxeh19rmrZbsOge+RjLh0jFTSrIgf8X6SL2MCUUKAVbi2LJxczvk42TZbWsqUa/6SuR
wnUDWU3TTbqYj7jUmqraHMyMmexl0fHNrNitw9AM5sLys9gBj3rLrW7EzoWe3fl07JxWXyYbwDsn
R873OP2j6QOb06DOw21Ctp6E3+KI6hc7gmaeJ0qqsxSGjgceplK8NjQPX+0ByJ6mqwOBUW3hyyVS
bAktN/zZn5PkrZ5SXqXWtw9ihmyL1lAalKBbG6Kax5M8nA7u1iNLlpSEUrZ6cH0ZGADDAU0kj53X
Kg9m2RhRuSBxpuccX5fs8vIKktiIGZHD1QIdcTrMcbCH0X3XvHQAVIyjdURIJEKMKWZspxL34ICV
FOAUTyo5ZL+x9nbWynwEo2iYGWO9RBBrczWpNUcsmEvD3WySY4YO18YjzoQW5Lvh19F5UJ+geplS
Q/nrbQlVv0VdMEMNHP6/AeI961AidQMZ8De57+r6ql8MCv5Yzj1QUNoscixEIJISXzWhL2E39UM1
PfHt0ZkJCNEORwvrqTa+N3vRw8oSYoITzzJT9353Y/0ao77GqPg2pBluDsIbDfWcG29JP6Clwx2E
S9kA0k3yilimjU8dpiGQPJ1omOd+HnKqPO9S93mHPpes4B9vy8iXBYfGeOSqDEq+mek9ThUHyVSv
Ktot0MLB9mT/gg8uRPLQr1R9T7+qyFxnZUux5tVg5LSD8pfNcqryHttICnYtzYVfPhUcn8I+WkTP
9O8hn4oebOqfdn7IFb9Ky6hUhpGcHUEl31xn536JbiX6vatMYiNEAKuBgjM5cfy027Q6iVltJedQ
oBEI7mLftdihH+F6KQAbLOL7U6c0e07bVoSNH0hWMqdKlfErkmmvm7wAuyb2l3nZOEm69uiBgkE4
1JS+9zNS3DNNffglMzhOhHSIKt/+mXR76/c/mnF/+Yi3e6zm7ovKGI9SbrDZ6WunjNRlnPCQYXY8
yvmYKZp03PQ8KhD3OdaF0/fRLLkMx5TY3K/igFBvgROwl+TVATmloU0lMuOCT5p3Wmau/xrjBjiH
cXMcgMGk3JlYZcJAzwXyuWjHgjGalGOYTU0XSye7cXFPYTA/HicxcJxCzYnesWG7JeTde2F2VTw1
PBeW9fS3yo9dZ8I6/uhwwRvSV6O6rm6CaLOqysxRbY4jbGmwJd5WaaWCY8vPCNk1AhNlubSF+6L/
Smt9gpd1lLvJcXn5md7RiHUFzqS0QFgtvLI+/OSG3cbkuHHQsOw8fkR4DOBmeDjeELWI/YL4R2yR
yEf5+7F2YOfTpc3b6ub79F3U1hMZB4h3lULEWZKhvfy4vKNl9QKwVb5mdUIs9kX89Gyjy++zQe4L
LT9J7giDtW5ykGaiJ6HKh4usP/zZvYXVMIY6vp5Fn2FSOTH6oZ+UBuAPg4ayKWgdmc/3sXIreags
Jr/WjH/uh7MG8cXPF7xCiN11yD6384BzPLTDY+5LwRDiCUApxtXZS6hD+xCP+o0yqfD/V7vHSNrE
UPgtqtChgOFgGoLuUmfoNKw723tE77iL/LM1cOpcvGTf8IjRe1BHMcoi4V9bTa1LXdd0IspbGiPS
Yjd9mVMW//VDQqWdUOnEhzKJCkMzU6y0fAqPvezQP1kZW3f6vADqbV0SM8vLa96mWdGKhBpYcpgk
nSrru67dVVKWp8nWiM6m80c13vhzobY5nDs64NI9YYmR5kkrHfQOI/irBESu74wQc0CDRYLTVzJw
DsNY3o7GrqcQ0eEu9q+X8N+eOXNDzplitZHmb3Bera/abn6PUxh0ojVbhtsNHGJZn5qYtdM7hTRG
m9rPhnVEybN6kZJ94MY1LfJThy6Yl9efLhJfCM66ZhIXiTSEk3Faa19Lm/OuKChORtYvefy9EFNT
IgK3NhmHOKz9mZhSh1XEiIwaeeVQODiW76trIkhm/qAEjy+8deR5G3+/mBtI9LN8ESEDlBY8in4C
X5UdxSoqdXewA3XNdwHe6pwbaw3+rtPP7OUCH22qgMhN32cWQnS+SzI7stxXHE+o22DK4lp+9Sxl
lL+hWFMFvCpSCPPIvvMfq4HAxPQPLc4k5p5aPDpiwBaOaPjGR3Lxe+W1HO1IuoVbvodyk9iAkZly
JcJC+kAvWcyXI+MjCIQkrsBM1Bil2KUGeipbfQhXpjFWMail5r1Pj6QRUx5kRvvW10rLoAp7XVss
KWovuJnYl9IBbzsMwMJGxtK4s94nhKlhOcIBrbPLh9OpWAarH624Yx5K9F/d8N2UwqfeDOaG9F/k
hmGh/6ICMGSHxb5AMPrztMxCsYbZy3ljWuLK+1T0QrkqZUNo2U1sIIXwrh5gbeMcw2MM29Kh+/M0
F9hYZBVRJIi9wan4tTe5kK+BgSRt6rFQADh/5juqaBEcoGwQiAvKzPOx1PTH3NEwfsZY6eTTUkli
WnJQDM1LW3L7zobSt5McToMRGWi0CgplDo1oUuCFv49g7BMND13uj0KW8cRglsI/fDtwTXzHnC/u
1mWg9Jkk6AuK1nJlHtrCxxA+7Ga2cZikFd65l1tRRgqxjj6bOUNgiAPhsSG7I2qg00GnUFzWvg71
s8s+hhWYdIndQdZQER1zb3imjntP6hvcTcUkfFTbfzi88eCwjDY3gocpzDyt8dYbVo2rqIPv40Nt
vM3HRuSvTUoh/wF/CV8IJsf/7NHdx8Gn+ALjOuE+f+S7DzJwXoDIUcmViaCkdJdGqzpwGX++XXnR
z9ndI6/WG20nDEvDR54Y8kzckDu377COK4VtfZiHfwgBn6wQB28jH/mWClhHaZO2/dIIYmIfwg3/
wvMr3Zf0psTZJ8RK+VmZz2bVP97SsgdeY95yFe9OWVOHw+6kCgL7H1UqnhugPGrxtJ3F5lFCZIq3
PmbsRxcXMLu4GkKMrRQHpRmm9TFfYRuYHLH9w6/2S0CURyjPFBtSb7j18zTnwm4CLHRrsudMaMzN
uG4JQyarYqzNUuL7ZC84NxiabRnDC4lnyQQdIqWNGilptlnU6S2Mv3DGu734Yhl0hmKXLhDhUz62
hpGxUdVHb/R4yg/A2/KkasaUwT++PfIxKViWyfaBgguY/XCM6xlvU9ckvYptKN3NBsAdYCqoHT4i
FV9VepIMTDzhutxK81b9pzbn9CtD/567bTHoFSegQkHMQ0MG56P6zUxi4kbvHRRhusJLfeLKP61S
99oIZ4u/vl7QHTfKhXa9g3mm5W3DxBPV6kpuWrL+Ouqh78Dkq9VSCxxptYeLWn0MUegjG7QYGqkx
T+rN2tLxSpQKEIBwa3sxq/YdjDpM6NhWIaum5Ydi/+aAqjeC1vKdmyhyt3wyIMtUkAcDZn4sjiqH
/NfgsGbfxAdiJ3A9qi+kjm8MIVz46jc+gHxFmbbwOsFWpqeT2ULmMgoCynCWO/FNAQqxPqFU/Gtb
qA98fq1d0o2+IvpNX5pm9Sds+u1NBUDybkSjsEOanPOPFF1+5uODcTDR4esVCV1sZeoEOo2rzyDp
y2E/v+AQ8Y3vUed+0cEjiu8k9Dz3Wae2pG/QzJuXI+PuikReSuGSoD0KYltge0IMpqazK/QKlP1j
AeO9EZ+GKoXJqGpzuBZ4X9ZU3epSDtk9WhoRJB110mlo3S4+75nV/ds3TS6TJ/nSAuv5tm4hR1Lm
n5A6SCMBkY9T1dQUvaPOzEN6RnC/a9zrMKj8z89DcGqoID4Pw3PqL21xwPr3RP/n9ozyLQFxanCp
cd9vYeSFcCRG5/sXvNdtNjEw5tfQD55vcbtu0ncw5B1A84gHbJK2r5bCYeQO7I9cesEPGJKaDp8i
HftOdsNMhvRzi9kjXbamgwOnl2Hvmlpm2DIm2q1nOnosMVEOXxxm1x1L9qoDVh3X6Bt3q3CgPYT8
+eBfoqBuZjI8QPriru9cSGq1l8FVicYjYZSmsIB3GcztUgUJM0jaUrje0N4TfrzcPLl40qHU4tZn
zU/6W8kgyZrOcYdNUyVBVOakjMnyv2kf5yqEo2xPCbfQ2UiVaTf3ubbsXwXIWLzaHB7xr488NEpA
+tZmSZGtrzbXIBdNUq2YN91Q1RWReVUY2jVHEMkd1sNcXJnhOVVn2yGjeUQctU23e83vUn0WubF9
EWwzARiERYtchf0kpA4UDexqW0qCDA6gGo0iwQBXd436I55PvHAXY5K5vT4N+ajohXctgHSL3l2s
zXgDQWQ8VpAbfw1F6b2UbnZtbu8OsunuQikWr1Z+RouWUXSERvW3dxS/axiw9RLCjmMQxyPoJYxo
sgu79E6adrkzz/kYgtu61FxmDF8BgxG4Kmpi6VBYmdCi4zwMktD0NNl8qBGxeyG9/FDKyE0d7xbf
z2qbATAryTzBECqGBoKlAKTIV+RNoEnR6fmXRIesqgzaD9RS9QHgpzPrZagFW+a4rrCLT3Nazu9d
mSu1XHeiA+dMdhw7KxosQOS51FBfiUWfRmWbM+EUng6a6rXYXFtTNiGSoCYrt9E05T5Z3KfMBIby
PwzEerQfljZMRZuFYqMioy/ZCSXnzMnujAzZs1wGxrU/hI3HpkU/EQ1b9sH4GX0JGVBBOHXau4AL
aX5M21CvuAWZNud90IhPWEXmmnTXCy7OFUcXqoiUjwrG0fscCjtTb2+Eq8bZMNdP1hxBAkSYXcnK
LATD6PQf4AMu4yMmrUB/spvWvEESpuRbdiU96e17gOUC3vJSvf9cRWHcI8+D0QDD+DSMyB9KuScF
Vig2m79RFjGPRDs0hHJB9iUYfmmK8cA3Mb/koiRD5Bo6QU7Qnfnb9FsMsjEeUtb5+nKjrZzUX2mc
RTiPK6idhMD1rje1YbZSqqrUTy06gRiALR7f1ddxmzH9VEfQEry4f83XG+O2EDhMzkYdjhUdqfQY
JbTLNnxY+I7ggU0GIrtSKZnJZtykKvecy12qkMlElYqXKE270AVQTJZ/6OXS+7g7GWtHKvZC7kJ5
e5vNZkie7K2I+WopGVjbfyyDclDwqKo9W8tTME/5spliaGdt4OCzss0oPgwxdm/4cu3H/w/H7sIY
DLZ9imI5Y6SfpeMWSrxCXXG3+KnIB1GxhgtFbKHh+M5N4Gl4rZ4rFBnlH4Jp5+OIDAqSHxwy9vk8
+hLe+WD++Btpi/y7IuVxMS+UHsdfzbEpJb7j9ffH6IfeAlekzfw/Kq9XSyJpWMwOj98dwoOIqizc
c7S51IWE+XUNNk2MTRhBJaeqhFWUDKKmXru+s+3JSi4jQBYjtb5IcErBUigZv9+v2bOtDn4nIHvj
gp8BgI+OyjMO6LP7nLgLam84CufaxnwWt1q/pvKFW6C9L7ehm3mhq4cSmsHkc8JmPgqlff7EuSCY
ZaUVVcXUD2TEYSNQ0PlWD46jrUnlAx29JOgjYLnxRIlMHV1O4aCIPrpgr1NYE/A/qoHRtnRbOS7O
dQTdNWnzOPGERfekA4Q8ZJRYjFuEaRnzyrXk3F/zHk7nisTb42veXUpvB8+6uXOsf/SvaQ4sYxae
RA4GCSYf7IIXPfu9FnLHxndO1KwP8fhEVY6Rf3gIR7EUXsf4r4q+7iYRpZglV7RPCni1sxuMJbUE
I42jEFFqngm1U9VmyC7Lneyn5wJtn6WNWx0Ak76/ezglnTR41GKMs9Tvkvh1O2C/9me9b1s4tGM7
CWix8v6qvhUDqcAoWx+4bFgFcvMr6BYHahm7gy35rE1q6DQlwpYPYx9GjaIno7pGp2C4hzhEb3wm
NzPzlbLU5es28wrnD2+VQrobPPVa2B2n0P+dbyQGCRZys9FC2p/IRYAWgpGOVO37VuQ5U4gYGbPB
pF3OOvK+L1N9n10pHvx7mjdjVl1dqduayCwAw/L1SsS9I4QFfbWsKBTweXEXXXhGuvdXgCdIC8L+
h4vur3LlWQ/4CPYGF8WiDsX1iKXYT8+zG7v/LFzYnSTZMJ9hy7Id50hff7jakPACz2+XaGTar7xE
9s7QwVOGe9hEo2t9Em/O5+Kj5Bqf20X4dKNRK1DEPAWKxpHe70ealMq8tNH5SASDPZwxAbNc8Xcn
gCYmWJKJhX7cKQq4/UdOORh99T5NAOC9sps2v9VZMqTvsfA6AvaT69ucFjfT5X0zj40NmRRSdnZn
G16900I4yph5PV6ufw56TZ3g9/WxNTTlpld00hmrRVAFfmBR3uxs+PSkWw/u0dpFDurSOSgDsJtC
2NXDeHIUFmkfEVZoIL24nLkNdX18KdDkq0+Osq8ed0el+2K0mgcOJXyp8fv6bIvAw/MEsoJx//Td
xk/tUGIt8+qczSk5uhnaH7OR3coWh/0bCux5F4waOa4MojnLvGGjsYAonY0S6qkndsa9+qhZsT1s
zLBd5ad/plTLLy5QfSWb5LcYnCw1IqR+S8G6Hj1Ky+7J6um3gr1W4K0DYUogjMdhmb4bP+CXGsb2
puyMWmtfWOGhQWFndd40CGskWY86y9Oue1HlxY2jC8/Ezs6OPl91BIKh/ckYUdlX54Zd1p6WYnxj
fVjZM0DyuQFN4aiVrPD6PPgI0s/vOwvdDVYgRUQXY42eiHi+jtKxT33KLn2mpfAW4a/xk6uA2eMV
L/uIfol1U2JQsryMWSHn953gHUOEAgC1S6pZeGk8wEG4aPwdhwO3nJ9EfnD+FKAzmuk/ko2AhP20
WhGm/nbrjVx44N9pPN8fsQ+m9kg4Son2cDNd8RXoAemYzqJujZym6JJN1Q6kAz2qLOt2kG92gyHv
ysxDvnt99wjCHLtAvfaxgDEuUUBZYU6FkMld/Zqvj8TilvQY24/rtHeAYZaVKUmOjboRh3XeryxW
NrVfF8TEBBeWJHxxkxrmoZfph2m6tRuJY1DFt9D362xDwDXZFBdumXOOPR1hfjUqXG2F8a+/hDcG
iGTWX4k400Yv/TZuW9IulpUMpam4WBKlCNevFzY3+C+wC5ETG+C6gEJ19Htt39LZxhpVlOIeCArI
rcczCdkFJjs1KK7wqJfcYHdfaMeNSWnmkX6TNp2+uYybLyLQGoBeM7TzJSEFX6WK6n8WlkfjIcHD
AUrExRzMeO9N5DYFM/Dut8qE79f6MYfyK9v18v8eS5GSTuMkwmKmfZg+bK56h88DhIzaGSCNIvFC
0ARUmXA4qFueHZQ5MRca8HaahqjdIRMaZGQFJc9nz8YhvbXr38ht+3VqEC1cGSvjsVNTuwHIPo7F
kETpMe6yPoGeAOMTguGteBg4bhAoDDYDMJ4O+6TtjHpERZtXQT9MKwWaADnfoJXpWTmG4FgzzaDT
c7xpZF4p4LS10SI3WWR7aU/ZweEJwUtnqV4ijK2VGx8y278gC642VUagV3f5S6I7ryFIkpfiGsnn
/+v3CWiSnKyK1go7lvr59VtLb82HN3kWmu/t0X4S4oA1ka3pbgzqtOD/bKc10fPueOvCowEb8nJR
RkMvvKGcdkN8UoibM0gwJgz+jzsLcRYhys5k/IO5hFUfrGDElyPquTzpeILFcUZy1rHS0Jk9LMie
Xg18sFOVcaoJec0tmaFXeCZtL21jCpgiSnqy3nJddb8XAfVxvINSmxS+CqoJ5Z2dpGBRAePzyvwv
aouqRM/yOs1DLv3oYAcF965yADWuTT1ffKN1lbKbmyTx8Su3jLAyEeC4AbFW0mE8C1F6QXCXet5A
GrsEDnDIXXmBja15PN7V/8gNyBarDVtC37vAc5vk530M1Jm0vW7XP7s6YDKIl/oJp45NqssriCrM
1zMxgXhYCAiz34hb1A2HpMwdExcUn8wM8M6hxDm76UueIg4AaTDkE1kwC5kaDDDnc/+fMOsEUkmv
GfG94CMY9Z7axmvAxXJs2dzA2JUPh0mBELrD2fm5WB5B2ieo9p9gtgO7S9+UMKYdGTAOlWmKMeSF
VBX82uwWk81XVjvFWIKKEebUThMsoJuxRoH3ctWNAZpW9fn9LzcoHisPFz9Lp+F6ihIGAKw0TKNO
U5xfSbMDxeniV9IuEkGovZ4TCV1UPUYN7frEojrYmN6D127mI7dXcS8N53dbNIQFwNY+e3VTq+XW
Pl3v+MKMyYBBAkgoJLYCRf8a+UeozV7D7rLNc/5pqVV2dzJUGquNUbrJY7BZIRvcc73/mfHB7GSG
03Xiowg0XSYpr8XU0lztQjgx9awXH4+gU5hNg4ktPxENitRIhwyEFAOrQ6PyIXtCTGdXtv7dJFBz
9qwh8aRI8j3NoL6BIzaVWDcA9gFslkr8UheyazVk1udQyYt7Py1SZoKNzcfYTY8GHzJyCi9jr76K
U4Cn+uIJ7k2Yovu2rlpGnOfz6iwFXzANdhzWA46hu1+2CIwQzOZ2bZjzoO09Hjeop+uOD/SZkg2p
tejk0ScJee1ahsGM3buAYlayslftY5WB6IuE4vFHjfJqg722xSacx3XYJ5sYxnp0RQKmoV0or9Aw
6N1L+g/buZneJLAc3GPN8s1rSnfnlhQkRkj0KkygZDlu5iE2/Wz/Yds0auQUdFmZ3dhdiKItIKXu
4qdY+2o0nIRNyAsvCjsuqGq0aR7B/ixjpSdrG9G5/YewyGptpjRsPbXDTrN5Sre4Uujn3CrhLCNv
SjH6WQkTEprjNTXJHzHPZ+zYJ4lnMILyLbk4St4+TIubYHcaHR5sR2GAbxI9IpT86yqtBIt2YQNv
cWVDHJTVDAgC+qbxduhXCJo7eA0QnJ07qlLXgD3Mn6HVg7VabstWlRw54Bwl+2PM/E8iWs6UwcxS
OspDcCsNyb9xYWsTO/DBUnRm7c4YGkAYIG6GQOLDIneXdnmRXax03UH4KkP/sIxVt9g/rQFjPUsK
2RHKjQckqi57xdHC/OnBLezfW6VY35AF68RSr7tyqUxco0LHtJAA+qM/B+IPUXj/g0Wk9vMn98cr
mG59tf7kxWXtqxW+32kFc6f45envsC4dn0D2WnLgAiyMz5HuRrMxXcBTsIBs3rCu9yyTCeRWRNU4
BDQcs/XB8Swn3zh7hX2QEQBtKYcv6xNzzcj/CG7zDZW0OKH70PBVECbbt6xOppXKAF+rnuB859oZ
CxrFuPLKPlGtk4/9reolv3ECkV8bpIj2WNBxGfZu7K2uQYkRj3ze+5TeOvAnNYQgroiSZg/0UoSy
iwRv8HSu777EZwXWwYT+zTwvj4H0Y4UgD/vWpG/vED94MkZQS/YieWGNcd+G/QsNE0UN9pLORoak
6UM3LeA7UfH03bzCpS8uvx6Nhnk2Pkd2XunjyL+6X5qcdT5eA+aTqn13jDCOu5ikSMYGPXvW08Ve
hbYolsL8WwaFLPbreE3TWrM4Y8oHIEKVH9YODcMUBSf3JIw2L7oVz2RJeZ/hvNbQnZmslkshA8fo
cm76LnOtGVMqg+Ha0N5cSGFdnz19stk/TOtFquQgzS0gHpBcKI7kURqdfEN9mgWnxcPYHWrC92mE
X+4IUyd6I+Ccb1cQ6sek0nhRIsbanqolZ9GoSKk45yaVW8ZTD21ZKFVQ3zOthO6G8ENcoj5N7Cuq
NKo06BlVxGTMBN284j/9qeItOhVA/1uUel5tNkjlskgIqKiFuHW6s7uRKKxWsdKb6PGSPGcoYazl
XYSCkg4+Y3+CNsOUGODQgL1dhDRJDR0Sn27G2pmSk0yTPGroIq+GM53xUHv3IHTVVTEyQhL9R1KM
+rrjl9DNVLUBatPLziTZJXBpFC5MToIjAL5SSMsbu3hKHj7FWwgX3WVwzQp0azLRIvtgOexJ1oEz
ETyp+v6fP7IkSA0er9DT1YfzXFZRA46KG/mrXWmxAnwIQuTCJvYjIDcRBOfyaItZ2qeGbxFuSDKn
/RDiFUo4RF7fGQmQ6haKuq9XdD2BCA0i+OXzJp1QG65zeY6Yu1s3TR68dDG6Ryil2K4vwcygQu3F
OvQq3pgm5HYpxsXLTxhbkSfsO1xy/25QTiDQDawEA9+QkVzbFISkfYZSkA/soazWD9oTmUnQfA79
R+zInFgJ/PUNguFQMvmd2823s8jKIa447EqxGrOAqBasueoZTVGTzl3NybSUag1cPVGa8UQH/LRO
ZHSdE2FGLUs0zjHldNQdgDHq6xb1q1zQBxTqELtkj8ToNtTgMbykbFUam/o+tseBaXKXDTBG0bZx
73UIxR/IEuVAkOEe0Z+fw+6IEy+zQCUjvbJb8fXk2TlMNTWtsZyBBrfc+G50Bo/G+UKK02VzafcL
pEZDQD/aIRlV5Mb4PMeW0Uo+zWtDY1CM5EwneADuDAs70ySagSaAr1C01Zv32lxlJfHaSDm0bqd3
hBsZeGfjtBsb7QmioA9hlDryHJAR+yQFBaEbQH5MMYZYzf7p34OopvO0r+BH71M6vRFXSOcZgDUQ
TwxRABwHqi+Eugwn61h4VbVzQt0DbzhMqDBm6Suq+yeoAgCaJUfiOvBHQh43w9YJnJk/DH3K66ML
Ux+VKcr6fKvSGiQB7mhNH9EpWEOCFk38u33oZ1XRuDj93YVzLK54XojAGJjKqh0D5jALoH3CYBpk
CuNLJ1HgNSJeCtiH8iSP1SEc/YWZZEkOyGLP39dpw47kdmKNg4z7CxpiW3cN3aXSGsmr+H5zVpXQ
Avn83rKuv1hCRKHwHVaFThcqS8Y+2xhkZNAmAw7GQSPYFM5hc5U6qrOR30XrMkkjIAePxxJiaE+I
npaUBKGxOgEQjlzTQ9eZFECfLCvymP7muX+NPCu2G+zfjo3MDpqLmMhYg5SyGM24PNU7k9KTAHqe
CBecGhNBsN9ir+TodFqVPF34Q+WxhSLZYSVdJLpFUyTbwp0gpYJtPSZ2NTxSkjfEYGiVwIN3kRNn
M+IMRT6bKAHw4gNdP8ofebeUq/zR5SgS+HmZ/PxJWyUItip8pjB/fEhOw4pFSMr10c0Nk/qO/ItO
zGhY6Bk2DwCjktmRGI+tbX7UBm5n0lATFWTdtep6T1eXs2esaxwJi9C/tmjSQVsQtLkOGXO18tnW
KimnPVK7HJ28+i7sjQAhBLuVsDrlEAO9wAjvTRkO/ul4s69R86z+50O3hBJoG2KijGOc0UkbGPKa
em+bGbnSWuVRPgnjJB8gLdmuaB29p6j9uGO+PYI0vsBAh483nlgT6PyZwtXqRA63kzZr7L484GNh
bDYVyjwso/eXnqJzmb9KTyKi2sctF19k6bkUfg2T447JSqplh4mJwjsMq7PCXcL8SZcYUxaE0gH5
rdbMAAlzASxUtL9LfcUMpuWGqFwxUPKyYmKHXPpcpxK9NM3T3VlQrsnsH9AAqAPDMzkrhN/9meV6
vmA6jAWc2MmyHxJshp+qqch9jEv/aF/GRQVY0Tf+L7Txz5f+VuIsWcTgfj9dYvvWYDgZSZ3kBKPT
T+b/2yC4NXFJnu8zS48iSHGn97Eck7cAfOFDbIQXPzke4ju+C21vLdK8YJVJ1idtQhosy3xXUKcS
ityXJwj2vRDJtzm7AGWrdYfOBuaghqW4vbzT+ZqihKPd/sR1uvhjb8zYA5pQ8pbx3qjLS8z2lkVL
I/9vpw2oZtxDqJWiiuvhtgrhgNWVK9lUSfJyEUrsgliIklvYQXAmz/a8IboCMErZ7s76sF7r7g4Z
oCnDIaMYLexhMBpDhXySAq1wOgmjNLRsuIL51nPz9z5V4a7WZu2Cyj0DwmTlMQ8W9w24C4oEz4KI
tgVki7TK2lgFezqRptgCjvY5O941b/v7D0PtvP29kr7bJSmbAG34VF5qQZs2iJLvqmXl0BI39CrH
mAt92xotQYuQV16aOBE3s06TdPRvIeW2vI9EtbvGDNu1jDehk5vApNgxhBrUiPpd0ICe//+49AZv
e2zNQwlK9dnU0I6Q6VdxmdEEd7IVvW8SQwM/1wFEQtboR2PmBONQDXqLo1bP9CfPZy5etm6qrwxi
hcOpy4jlZ8AQKGVgoFXqfa4DQx4+cClyIFWt3lGIeoHtNQbg4BVA80PBRkhxgLPaEYtPQbXU3YYn
x+93OvY09aGQ+V73Mn6hGQEEkMxdhfxly9SGL+Ty/a2K/7unGuqG+mqwxVwn/WtiMWvXvKoY2qfI
t2PeLMjHoRprpT8gDlFhQTk/1JQ7V1rK9AHFpDFC1gcxMKscQVLL/9oNVYu/dmUyfLkyUGN7MSiN
MUDifIwlC5gSnnidjixS66xUiaj80eLqMN3lNthz1hihW6dFnVAij3R/QOVpV2duoBqyyl3dCK6s
lJQNCeCs5yDL/I7HTYGvY7AKLiL85EsOHpP9dguu8i3CNTQWr+AFmo1yXPCJcpzKEsnkKyNkcjZb
FMGgugcI8iYnzoyWgsyKZbzcN4ODOJVOhg0+YDABSklr84koBVx2VEayEsIhKHyaWV1qt4hwvY3X
FuQPJTddM6hFbJ2INZGT4pJlxPEeUlb926bDzV1nfeGeedYno1kPkTiTPQE20k9OavvW0McdgTLO
7R5Yvz9M3EJEDZYpaJ6SiTUIS2twi5TXPNZZLc8dcvd7Ws0QYNsQLjM2xw/jPPniZOsdtIEpXQ/Q
vQwg73B3CFJTScU4L5NXGbdJrHNQlnHVyfBnANIkzbPY5L9h8PK0mcOrZKqRArZ/Ga1XThvd91/E
UbNvieK69/vi5wMZu4avXVFLewBL7hSr3EuuqpvbXOQmsLBHLYxIbTM/XaklmAbbxWZkg+nRUc04
H6VJKTlwAb0vWPFUYdwELjQunS/LdiC2GsS9LS6o47YoInBkBHkRW6upSgjqTqU4tvdcs8kLooC3
9IEuANVvfpuTpgwuGHaiALlXAOqD5WcM9i9XJ8ynff9o1GxsimuECE1OPsok1dv1W8eAZ7BM07g9
Npi5PyLMhEyoBVZP3HWFZFibKPPU3UN9JejeDuOeCFOC6S/6AOqlAXxbb5dffSNYGlJ9tevSpM0P
6CrI9NQM5kmlNOI7AFx8axRf+u6l5Bmt/SbOHE35d1cVHQaUESdT2fPwZiKk7QGT72rsx24bdQbF
ejKi6oj2TjI8ycs9LfAfZIDaZ7dbll9yRs/VCcgI5IOiJH5dJYmvaNXXtXEyomrPc7T+StpBJTHq
cY0RDvTwcrDArofE1rPypG3x9sP0w4QI07SC3xx9mT8YpTTNNA4RTm8eEPO31jctGPIF7BIiB7Nk
f2+wIQ86sQuze+BnQcKfc95aNmUou+wbTd+mazQf7lhAhf6yRQVE4+LW/MKAtw+v7hsjO6vkyMb1
/z7eR/aANV2OkhSiwrvg2r+zP2MKT2DiO59yNC/ZE6D55EfGkojzX5nizPN1dq3TGU+IV5U3x7AD
NqS4k7q5mnDgl5c/IDxjNfBmilhTvwx94Vk9yRoRMbMt8G5eGG0Svsm1hD48nx0oPaM+VxzzEQQl
hF5kI946g/0SWp+mpMb+xEnU3TkTJLyoQRyZbLbzR9m/sFu/y5FgiLEAt+JSCWBFs5x+mkGLTg+f
9Whp2Vvj5LXzW5/urRuvjf03Px23dTmn9jj44XB7HWKxoWbEUXGDmMleBvXvcGxtJH54sZ4eWIwO
5fC+9Sv/2AvtoJMw0m2bDHTUBldA00UYc8NoAjRruYPXA8pWZDF0eKXAm2YI5drkDd2yvTqu9KeQ
uzkRIK5p5U4G9cMmxmRVu/8CiuUbUou8aRkql6JLEcCPSF6A2IHpQH8yDwLc1asPGiTkcCTUgJSl
WY2rlgezpOKVPynrABMUYpFajbytoB16Y0L8Aeq4lSWA/02uxsS8dvLbqrzIM7RKm0jUs6TYo4GD
v9irZudOQULh2anudYCWhiDzi0Ll3T28r1rM4tliB2KQwVtETzDjGwEjW98O8j38hRbcsj5yhoVc
lisc8ThBuCRJ7qpS1EEij/5wEuIsMp/gy9YPFNkKf8zvhB6+8BslfOJefVx/HcrpIIdoNzAxrRRs
cegZEpB/7BNe3Ogg2wdbONA4yQTOF2luE0FVWY35+vgaq8+Ux5gChpDCbhMDSU9OqEijZszOj2dd
ol96ne58TT0lFYJkUE86bKZc7I6GAd5dwwnZsy/bno+oEyr/Lp/aCT5QJL7Hp6QbsPP6WNAkUoFC
EPP5Gzf1cZSnNA9M3nWkRh2LDjnPrg6JSR0fKV0RfQ8Xw+mBwQ3ObTgyx3ju2A05nMJZxbQfwK63
x1xyE6O5O6pqzfCfvlMx8fODIir67yZNl1+/AQ0YUldMSZpCPn9drwiL1HxNHdXtr7oM44iS9Omm
Yo6cY1Ft/uP2f5UrW/bNjTikxDHSsYUaEOODClpMA2VaHUzrHtDUydJr31QiqpFi4kmhpj9nvBZH
agmbhz27oRoRERlbF5XqIZJNUGLdDd7eP3/wVfLeO1GbPTvQd+Sc2KagIzrlcw2j9lOmc+mMCj9g
YZvcYdKNTMVdcxWbqfjfmmgNfpHGs40Aa21Fd57V6LTR2lCsA8GiHUp5/zYQauBq6hJ4t61BRVxA
zOuqv5YBQIhP7g3Sap6zXtE0ddLcSJVcKFNhBjZoAeA0hXl21Al2zcwklZh/LdG9+Wa4eUkca05I
lhGr3oI3RMGjhzF1qvh/OMjw878T6AQAzldxWG+ggJ1sMhQYwh4Ab1GfqIP2kwQJIYzyj2t5RfeM
sQJG7ZTa/iLpHLZxTxHUTFolsJcGnFgQAWE1ucwLvRiaKTlODEzu8PeVoB1M2wjxQDpdgPjXpBX3
n4XgFdnTy7TBGRzH3yXHQl4/6lBFLFaWuHBUjw1sHgY9NS/Y50ceCRZCElcIbgv09wpsSwhIO/hB
HVYwMaKqMc2HFGHGxqxNCuFvErZAzQfAURcDueBiVhSlCsrAeNMHJaJ+7hMrY0Z6e5y3v91MHL63
yoHTIr3qg8vkS09QuuZqHwEdjKIMlLZaJOXDSGODloi5wkABEmwYeATFSGkB7R7RY+ObF+WN69E/
0ivABTJTIA9116FLhT6Kc5iScxJJyhG8holWT87IakqJQt2tUXykHegUXPvRjjIxcg1uu0dY/PnW
YlP8aX7EHKJsp+UddSnU5BxgygnkS1FGoqgPTux9taE3iNL3lUbavr4KTgvznkqAb5SCQAKIX4s8
urc+qms1fHRjd3KQhKHoDyihP3RZGrHPhS7lNWTmfFJ3c7w4jvmsEE66XZOjGUyt/fc0LNSiamEU
Q8Z+bvxbaQCSg00Fn3hh5BqWkByhVUGuEvCKL1Fx5+M3f+bAvIkP83aAYrtLL0fLzoTrz72yX90Y
RDvckDH1itjuQo/EJhjywu85yPXxjsO89+Gu4tXPUdYj54nQc6kkdsy0wrvZDu7SGdQZKmlxj/a5
ajY0m0qQ8dp9XU+qe1XfrHQX4ZO5zGTa2y1mblzg4zV26I3TDMySVcD+w0csS8fr6JAyPHCtY6wk
zOf6F45kflAvVbwVhCyzUsgX21g9O1/nXhWKz6s9UxiC2/Jme8sVqdRJB0C0gbl6Z7m2bQh0tFO6
67PEE7+c3/PBdGow0GrtgP/r72vCp3qAhLce5wN65c0nLGelk3gy4rwpu5jpghDssjpRAlU4JXfL
SjKaW/Swu414J4dCJAM/my6BKgkjutwwkdKdJ85Jim0iILLDdHHp6x+BmLimDg9v0zT1cB6lFZsi
yfEC7CdhdOCeTuU4M5hNnR7dRrb5QWTbr8rRSEsZlbnXzb0CZxnXml3CutsD/zHnS8SNchGKcn5w
n/O7DKt37XBOTkDVAVOPcAGNma8arMrl2Lu+HWjePpSI6KjwnDm4aaWJ7MDoiO2WeQ9s3XBCaZbi
XvPh0DcudKakUNPg3cC7brbkTapw+/Dil3vSGj81xiOMCIFNvNqq1a//1d9JPv041wskmb8FKSxF
l2jjj6y8tFFT6co0Y+VU5/KF9S5gFyVYGzYeOxOJyOYjRkqWGpLG1eJqkvzoPcyCPvkVG9vaUWVd
83FAoTHDogUsokoJGVZgAYbawKBAz2f6+P8wmGyBFYgsz4/cFy9ueXaGbotPirYJGWZG+Z1TXig3
TpdeuV1TMveRqWg/w1UeI7a4m8wu10p+J4KcNxHGgK7mZC816iJDWljRcue+xWsMu3hPni6lgXku
9QHb1nm9RTZeOIiyC+fnURkY+SXAz+0FmS6xmVu3/nREZlLqyqfjMvQ/8srTABChZXaX7qNBpWyU
rov5KKHt5Oc7vnFRfGoRGSfdLL3f4rDMXSa+qhJmq0zGCRYQhzBDj43dhdFSsuo6KIV9cn2RB/f5
tuAhnPLfP/4aHKysXE50sz71DgZmQsQ3QzOdP9FPBhh4KrcpDTcq0aTHogNTt6tTehDL2P5jsHEg
2kTPppES1qyYdxCrM84oHpQ1C6VjYUNpVtSUb3FEqRm3G1jQMVP4t8m7N473fu515XW08M2FRb7s
fr9jHEIb0ZrWAqD1hDjpFlGMcpMSKsSUn1mZltKut+48nAKMQJQEeSt2Pm9rL7DJWbpppX3KCriR
TZMzrWpw7beLmBUfVih8ZyUcI127fU0RiDS22Uj3UWY/K1pm0DWndU1a7276D7uMVr+xnW39TNXL
Rumj8onNiTiNdFRhOlWojTqwozxxbAv+P3WQuhHDU7FYGLx4kGrbdMNyCHtsRmoKJiQwEPoH3r0o
Y1mvLjfG651jx/N/u87JFHxQUC9Ip85xFujXxO4rs06S7Z2Ob0Sd61m3KktC9Yuw7D15qIN6cquA
205sfl5swQhUOCgWhGox2zqvzgINBEYBsMDjilk05xG56gxww7d2NlLIPNsuiglacwuiMrtXkRAk
xFyh0dRwhHiXERDu8kLXcmFqlfvJQmtitgyN9kPgxgDQ6sgOy4TVW8DFc4IwA33+8bJwUEpd1VfW
4curpVF60C8Y6OEfu+vyS6NufE4b2vzFRISK86BO7Y4sXuAwqgfkLp/6xWEBQX2U4R5lXrT5FRYs
PmeP76EHEgmUSQQK2gODNeKh2w7/RNuliITnhemHcsviRECDaJ4US6ZovcWuLtAhWOOBuUPxFt1n
n8C0AsHzCr0qbODs6Hbiv99VCw6in+6RRf6s/pCU0pQROU7XsG1hyBUmTCiEHwfC1lQI5jEJUKax
4vmBZppUFcurF4UgPDnK7Mwfz2I7wyfsy8xF7ySgHpHoyR8sdMjCoioy9i3rALD87E1e1Dv2qjgo
0LwCpZxNg4dsjk1UNOA5LID9MsxoY+cDFlc7mdG8iBafrVAXx9RMbKqCc2FXZHI656FhDYm4oB7R
WSMi23QdbBwqGE0bvyQwMjn0D3jeuGi9f6h5I6NN4WXRn79gXREv8VkAHQa+1aVwutQHyY7O1z0I
eYUye7bthD8yDcmxQYVjhQaKdLhwzezU+SEh14Qreea8xlgAB588vzLTi2zMlu9IaRAsC/HMHQHY
CxuwFgRfaWTVyItDbfjmP7nOCYKfhCwmyD0mB/pzQ4OUW9N3ptfsMMX/WsaeORK5cImWaHxokO7x
7Lwp6eHPlkB5gnEK2LTluu57Fz3HWSdpPfW6OTKnhEo4BO9KL9C2ZRN4OyqzKwMADBpkCByDSkks
ieevrV1lK90M2KTUeCcLalRhifXvG7MaUriz44fyxhpWxGpDkRnxySYWggzLe3q0lFS2N4z2hymD
owKBOkwBFrwE46BboSMPK7tb76jYLhc0SnOuTRQ29t/YAXjaqwMh1lu//5da/NQmMzJs+51t9ygw
g8S8/pZpbhSHbi4tS2hzdJVGIqn5xMyaNG742KAAmFxbfo463I47U+VDhihwMPqcu41KvKieEAI2
ET+dLY79OMlS0foOfn6UmsyNcgs7GtyEmyscdVuTNUejqyOr9OQQpG9L9BjGhMgaeBbvDV1MoUEY
x9TjcfzwktKEi28dI8tTz0EN7wM9zqzwSGkfnzUSF/0myW0Y5N5lQR6FQ0ffjyd6cgqnEBoIGgBl
Pqh8CFbTWSyndjR1F3WT2rVCy6wTd0hsko0mVgPCwOS5a+LPban8KbrPvfyqUPZm3gZfrlyFDMM1
hP9sSjSRHtdJrlKO7NGESmerwdXiqZzoduYfLPwufZv123mvV0uPKMrzo17i3kZO44+KtWihTffg
FzKqFPTIXSTE5DBAeyEw5jtUsHcqQkN+z+W9eD1jL9hHflAle4oXLqP6QlWQfIJn/MXBUgrsbZsV
gsEGDpt0ZrYhyOIiLBSAF2QR4Fpar4WuSCQ12/WkO/ME9UsGLdadSkjiHIB9mCyOXYq6WSBvc9yV
t9w90lPtnlcSYlwmgyof9bBMIbOKAHpTtFmfL+rdZHgcI/XNzAOEVWQWbzgdmxg34OckeNKggxFt
SLTGiUcb10nbyqqTeeCH1MT0qvjIpNRsJ6PZUUsHGE+kW+Wfitz8/jD7fLoe2KNbQTRzX4wYcEfK
Yn9OsQc/kwnxtFelWyYpK/rrHoNYaHKeV8ADSNCHgvP3SnuoHCF7Fl5ddDxMvup+VaMEhWvTpOTJ
jobK+gKuaILnwWBOHxyqmZPI+H1GZF5bPyt2QcW+iJ1zKkK8e0/UTsJhmnR6CBbeeg1R8WR9CIvt
KccSoH5RpWJ+8uALinHsk2Wa0NpW3e/gco+pY0l9uKIVfzwH4rfu2DR5hgHXF3v5yqoKYF+PLImo
NQ4qi1UV/pUrg27MIiUFwWm/kPPtwGY/0xIk8BSo3+eHreNZRpy3VwUKdjKaITu/RVD/4sgbV18o
scPs2/mO80uMlqoVWu02zNhSeO2q4lVBZ1O5AizysHOjwvsOdhYJcel4dKVuEcc10C5Il2AgBOTJ
aShT5VkhdCj0gILnLIbYzLbtutTVO+eZgMjN3a3swcPoc0l+9UW0897fb7+m5C1Cojebb6wSD6zi
0Jl5Gwta5jF8QJSkdtPfdL4hUa85fwctTBJke9MK+6LW3W69lpY2cX5Bkgf/AdJV0vwagv3NxZex
R36O8YqP0kVb5SscPz7MxWgrWgjcYyZAY71IMTs6KbAOW9ecAe+Qpm2GV9SllKu30wMVmfjuTK0G
HqzvDDgDDg7Bam+dVU3p6dKwBLXCgBnpCqv/uHn4joQNZVhzPGwTNI1+hB4q+Zr4pn3tOQs9vrAd
/WhthgUQSRSeHrj3nWgZjwjvXs9kBIsKhG0zrzvr0BRFPcNDS0SciA9F+8XvnlCFLToaaMUg50jR
WJbdUHg1v/aHBO/+1BCHNHvPnZnsm7uXFci9Jtu8RNUanHeTIB9v/W5aJKqoEHr9JPOqYrJyTgJP
LEdqB6LpyLFhD4qhRBFIWcPnyBXnkvXdmOrI3gLsACH6DFxVZ0UcKszW3HUeREhV5Vjegf4F15St
30OJBPL+pHoXN57KkP50gcMHyhMRw7mGTNJc7JeEbxoUH2bUV9RZx6lIhu4nH0J2Afbv4nyQRUVT
WSic2P/fE/64ffeteEv03rSgHTeb/kKm6pvAZrUZATQeMkjgGkReWogP7mB2arqijQPybAJP2vqy
EB9vOGOSIvwAMlAufWQQvaPKbE7p8bETpypVfSicZ43/rr4MXQxgggnVe19qi3WNWu/SBXytDE2d
pvHHmZO3MBia4A96yIZp/TSDDzykbeH64rgZQLcnAPh9MAvnOqSfwohLP4biSZlTWN5TF8X9RTNE
AuiLGuycS82yxV8sP598k9PbKddFHOZGNJrTlQ9sonnvmVxYc6olK/4x2zFu4tMBGFqOy8Gl2VWK
WBeoR3LI7vA3qxttEVlfit0nIaX/ucaGE5fPfW5nMLUbchHSAqmLNSAJ1cahNHjDVXFFCbEZo7Xy
RZ2pW7qkH9T513qkVuSC3S13c6QZPADoKIgoLwyMETcroogrgMJafft0bW8D1CaKSSGkMfdjIuej
Ks/qu6c/1YJsxuleMGvxmcYSCUbVunxgWagRFz3PbpzJmye0gcMYc4YduVYmgNjTx6On/ICWa4RW
Y+LujDaEtxm5PDCwypUeVGanaaF/mNVK98PjO9iVPSYu874sFtaAIQq3cwFFob1DDisrMberBK42
WgyQOqIn0YMZ+M+wrR0U1J5yzlyn+9SQ1i5aE24ajc2868TYFaiZeyyrNH6zwrPDVzQZzbXvJnS0
leAeAsP2DLSjBOW5CS1sttlDMEGmSwl2VYUiHWDGTbHppcmGgrKzNrnZQBPyNza+L/U31fZBvnU4
NlIlzn23lEGgVcI0+IRAqY0xrb0LevfDCXE8vH5wW5OfzOgT79Bydq2nzHv0Hu5Et1rON4EJeWHx
lnudjSFK3H60zLaxhO9i95ZWu3n/KaRKxsf6jPr6SIEiVBJ3hNdQ/uj4ltxfOyDZbRBn7Q7sEOQ3
cgOud2sa47iiQodBj/NrecZRd4Y1jOCEPH0blT5zblZO8TWHP58GxJw6EayJYg/4KSCn0TRFt48u
2NWrGlYHgwB5UJV5eDVSEFrVR5jdUvfXVyPchEkiEQrj/xaaFQmC6O9WA4kEo+nNdoFRhhaLiHqk
rBkoWDySt63CjAMvyhyEzC5fCQcVCZK+4f1eqwM+O3M4NzjkMUjQwpB7cHahnrn0XSV1JFuqMOMs
RqIRIdSrMTowkmgZqUyu52D6Dni39FZqrw7TaZ+OryIC7UNncmqomnmyMCVZYh3LmYP9/VxOTbGx
qtYwtzAIpqbU74Q59YzHe7jCRa2YUS/8QCKqQsC9TYsBTKwmtScRnjrcXG1xONVMgQPw+C24Zh8g
2vRFjhiK7lB+LVOjnMm4d1TIKWcSobDDaJO8klcH/EXn3XEgQrYk45CvdqcrHWiUBb28EZ/Rl7AJ
XrkacXzVpRaxIEcrfryY0jB1XVjDNecSFC7zlgKsSF965aB0HKo7pSKKW2UlFDunfKqYrrRT8utf
LDkg/wEORwEHbZ/ui3XSdDGeShZlbv97c37+fPDG8y5osU/0rQ5foHjjE6BMNTVOePGgJy3k3VgO
EgJ7wzvL8GdXoyOySInr6bpV4eCXhWlAi5ssZdMjzM3rfjvzWjkuujK3Foc9vZ19udwKEln0f+oT
+FmIUuWL2XxkLFj7y8G1eohoOMZ0Q2AkexJhxvhT6MwhVi/oMveKlGvYLX06opTlfPVyBscdoc19
xO3O2EbFI2Yq5HK+hhoGwhasYCQXor1lNaPWZMwxSSBqFwtma77ABCtjKly5vF1Rd3uo4TgiXf2+
rQ9o965EwARmmGugqL5ZY2UDV8Z79mQteTvwac2wDS7V5YXprn88YrO6pEBI+KKIvMSgZkHWDQ04
1HoGsOc3+D99nu1FvrcmQCYj09ai2ykkj/2BlKVdflMrPrBoQHY5ybhuAcsa4lTwStwBV1jJhNzI
0Y5YWw5MFagFDCoCPqBGOVc0ytas5FZDZ5/u5GVm8SKntHLSNzv2TdeKvGta8/eEJD1xoai4mcyr
qQ0FlKkYucFRpC83UjE+IsNZi6T0DdXjn9vo66ClJkQbclt3tK+4sjrJwLxT+iBzFtVoiA5IlVpe
8AYkOAVIH3e6flSsOGe/9R5tTpL33edAu17FFxnyLYjkyCA6gQXoXjmGw+npKzV8xaxzrnCMm0FY
btNqI3DhsKGn167icfXYyLXAScDbH7Pk4Pn1Do7YRz3QkezMGsfZwRSgRypsdje9U+9XHrjkyJof
S+5GGv3DYCzWF1B3yJHtOK9BrMXNE0DMmea5tL41QFZDjhgE+cvWq5JaOy4VohQFc2Yzma3wCdXe
wgVoXz1/pWHUv6nBepNTspsndRnQknA8XtxIWqc/t55KVCbjMvDiz8QLyBuSKSxBYMF/BuJKnVvt
H8vYfa8LzfBTHu/XO+90TQl7IGddX7yjhDFMuCUnvxUR+UIrpq2wQ7OW8qh6S4u1QLcz57fc7jD6
tYWNhw17OVfNSd/fM8buvqBz8DiT2V+LhpSbR/qsB74VcxEMjvpHtqFvnlUx6uP1qwBjBddU4F4a
3ZgdexXbhepE5zPpag+OWtQC9KbtC8CxgEEeK1AQUpDIglpcy1jN0er1gYHn8uS/oY8J/QJNhBEj
x5L1bLR/gjq2Mp0iAYegMyBriK86mXios2s6QB74HYH40UvIUp5sfa2dOUyDXoLFKt3Wgf/LGTrZ
E5SNkxlh5kVxOtcInPQGVwyegjhyEpvk3Tru4oSh9ohsmtD7l1A6lnEMQfamyl53rZG1j6uTCPgN
HUMVClTIh0pGEHOyqjkyMs8I4V1LJdkDMBpbVpQQclsDAj7tafDkNwSOojgfr/GSduCOJtdbV8Di
cfz8oakBFTNKXG2YXCj2IXUpXlnLSMUzEy+MlBEa3aBpY6H+i7EQMP8JDr1+cnBjpDtqTuk/nnpt
IPjT0ANN6R/IFtUbvdLjFzd0dBTFOU+OZ1XYPEJUByHad+iXF4M9kO2PumKKRHyA0yjBC28w1mXx
6mIwDAghR6DYb/FAHoTw4Jft41mEln4xvSJje1KH30rIBVV0R8D50wCEm0XSgiT6em3R0NnYEK8m
NRmolHimeHYy3o4QYD1Ak3S1mCkj/BzxlTaKcMlppeej+0HS/C+xC7n19dwFh0bXg9aniSk3x+H0
mEtoo8lh+9nm5NEDcDcjPT1xKHGgB+3jbaw32kvf4tXiizcwWIr1diOXKNnl+kjRUXlaXIbs8+H1
aNBePlHjx9knq+C1YXhx/WfIvIy4iaaOyee1EhFg7L8UiROtOZUKMk8ywN1yb8uhLECv2QLpNPqi
siiYWI82vYC62A3aI++3QBbCpGU+fwkiBUL2RbtcQvs2Piw7cxgRxY18rftzq+DQGcWG5/e/+i3x
FR2ktNpqav0ChmRnzTzngFc8u5IqqXlRTTRfbY/QYDFnHemeTh0vBsRXgG55pST16Tqma3mCgpHQ
1ZgDoIBo2MhHdtsKIEM6ub+Byl9ApNpt5JbJV2t8Bw1m85iS+rKkL9G6/zUFCM9u76bp6uR6f3Dg
a9LuadnD4Bo1c27r3nqu/gtvr6eJ4KUloMxy+UBODP406+U9xYzeply3i79dCa3Y0anVcGMrcG6L
9wRYprlQE/Wmzkq253ondhG0+00UW9YppM++M0qbjd4fnQhz4OQ6lEV3bCuJmpoddkID1sItL0zH
RZlqcNkrRDnOpS1rrteJmjrLrdSsM6lrnzwvh1EX2F4pTql7SqOQwmRTRM2yrE86RAO1T1I7UpYP
Po6zjD28DFqCcB1IhXTfh6IshQsS5Bm6+w7zbEqda+8DLAl/+zGHyCHu17jpEVe8cVbP269v+TFB
LySlJcxDoxIsvy7MoXmom7xSqQLoJ27L9He6VY2vN7jBQI9DOdViBz9aUIjLw6hYWRN1QM2tas8j
VSVRtSnCc1bFKdJktyOhCkNOMJLQpfSqqPf5HCs0KOYwvcSC4GmDN2GNq3XbMr/STa9Cf94SPHn2
cZFo9yq6h6Kyu4uuMqecLYuTGvmWjBYYsbbp1o3uvYrc9vbrpPkj43VHzp+5fJniL0+DmW9htYFi
DRRFK9YCIzi1Cko1IfNX9rjREDErmjhhsBsr9BhS7B+/JL/uc5oFIv9bNYuYYLQsKTeGQ9M4na8C
fIrv4SNYDYYjCNkSqek7b5aI+e79ehwixMbwbCDG3LxhRWioIC7LSQsPHzvmxMrDZoZP/c7N/pOP
OrR+PkFza4i8HmVxSX10s+AMtSxjWmjNHLQwO4eZNBz7N8dL5B4bVs+gXo2op/ER0L+elk2XsQnI
0xdcGlE8kPP/4ohFl8d2iiAoFEyVddB1k8YzXcrsTDaf65WVqEwTpxcXJbB5uv4B0P+30Wd9WCbs
Cy6yoWnL1foNK6Bg/YnP9Jo80GMHF+woZVCBNbKjIUSmYDFz+LzMigdeISjp3SXl8hjdyVxvNgU9
xQmplWorKayh3iakX7KXguQLYsAk7GIc/Uuu0LCxEvAAhamzhp2gu+Lu4Cefp2+GFmm42asmBsZO
lcHEFn+40eE/7hLdLMCIYs59C9T6OA/Y7QV39Kqnon8v4hz0E3vaCposWForTBuKI+epumA5npUB
LvZFxM5TnlH4oh/9ySFQxzmchmafuvIs4SbiHZ9b9ejtH9oi9YPyMRAAmtsihtfDjECNcbgXDDJY
/1uo8TkER7r8idFW/eU2meQ9eeq/MF1jhZlgiSmiOmq6mYoZhBjH+wm3NtBWmeUe64JmYjmJpeUm
lxAivbred5WeS3MdOLrvQ+35WARLaXGjkS5CMCSfi2l9M37OvL6S9G92G5A4fBMDyREz+iyrkC/K
X5ABUXN58m5kXYMd0J8eBOz3d3vCcLs8rxLcg4RIvXHeBgLVT45hrShGTBEuobVe6cIUR72U3A54
1nNqmpbBztkwhHQTtIkg/nTTPNthS2pMOSd9hHph5bGt4nrsbWumMLg2wMs5JNTKEo/xyQxgp0hE
C8PBH5OfMND+Kbz/1rPotQSkwRJ32yyJbjFiL+aKNVMYfKW4mC4LlyYCq0BjCedWi8cWjJBNXX7o
bHuaBOJK1XufrlMLnzhnEd+StUpv/hhiiiVlXxA49CGE1DHkP+2PqRqu1ElgGlXqaquKIc7uoDTP
V8ahAFgFjZy45dDLXo6wzago0genwEao9RZXJ5QalHlcarFldqXj0AFEgs55ZxTCsYqDDsabLKFf
HwbL5gIziioF2uwLCayPoqTXbIbLnz3sM6h2Tn6ff7ezPhQhBNLraBhXiLrmpkYa5NbXuCSY/W0T
hsTM/7f79bKHPaXDh9Hg/c0iWQDgTwGQlg4FuLsUS5HV4Pfyf6fd09cjA8rm0aoTeApUhD7V9U8N
P+SgynbRn8zgXtf+Z3seIjS+FGxqwWaqHtLX/qa2ZEmsJW+GAG7Y6Ca+IBNLCFXXl3dVPwk3icJT
QeM2mucTeahrSBwpBk7Xsej0uZIaHY4ZvvX1foc9gi/jm+c+WfDTw/GdZEmBrER9yyDacIcpP0fi
EhVNovPv8TmD+IJOssr+Pktc/OT0jRZP2+R/rAYBMYfnhM2A+Q/TyP2YINZovl1jkOB/bP7dts21
u5LfIflvrsz1Rb12sRZgAoQyA8kJ/Nrv2vdew4v1F3dVxmojWnJV7JGctYeEfvrLdGa2MUbqe9OG
v+HxooDnroUzIwpPl/v4tddfCBcDEZ8XGMeiPUQZZR40zubhVGyfsofNyobR8epd9rDKQeEZ9VHA
xYDGDxzbRqAQXKDXtTxir2n8ikTOfiNM6qruvK2ksIfVIJwiN9bD5xm6VTQEVqskYzCxUq2BlfqE
UvIdtSrKXqI89biR8GF5obQaQqr25GqwHYt9Jw4hCHQuyTIdMXx6bex+b03X6d/p7gV1ZjpMlnaq
vxRuxs+Ojz15UoTfhmWdcMJeMTrgkUQDfOuS6Fsh1AKpAa6uLBMIFvXmR0fIrj+MsUVm2rgWwJVi
eRMSfU+QujsCpEoTnROQqNDVd5exvtaiZzE/JGGNy3UtKMD8/fysmMSaec7CXFFX0M8C5/Y3wbnI
G2EfHEAGX5aA7Md1nyCUoUEWns4UgPXfcn4Qu/r1iNRgCngt3QVOTBFh9MWjb/WFJPpf+NC6AHgi
ZCKnjxl2EDnkFH1D2jgF/AqHaEwIHs8Wn+Ak0Oswgwwdsd4lDIN/K8yeQwZYwm2qfMeMTvegyalb
5Ud5g44MY+qwExA0/Szl2yqr8EK2g7n4VrwB15keDZ84VJmsAnt7xCqlLTgbRgnbOOclkXg59dtn
OpNtNBpBATf3r8j0cpt1EbZeeumC0ozMLMUEHc3uGBX7kOfY6YxQ7HrUJCkTpAbaVShJaClhkNIx
OnW7+Mitbs73n2+h3UmXnDvPPKajMoK+dneSsW/74r2DzMkWMG1HlS/lAFvXIAu7D9k7Co1yqk4e
dindMgkEuR5ku5/z/kclKj8QRYQi5s/RPpLEOAH6Sza1yFNFcjXNBYNMHR7C+JdljNJArWNGHUhb
2TGJTMUV1k4ilZPAHNRveTm77TcLpIh6KOyKq6FDqOdQCLAuVsDuRLpjtjxjfgHzNfd5s1N6taHv
AoGQCzkE/J1XS6IBfyqkNV7oiZPZtuSKLzYrOGmr/vfwBaWFFR2IiyhYuivAoSiYcjiGbzcB26eJ
yaJjigmljAGi128Zbbx+fpENYlg7ENjKFV4rdug3JGrukCTxYGom3WhrOTVu0Pr8RvjGVCCmuNws
CbMTg2bj70R/hmuRoBRr3g8g6/mxjH2igCw/9mvNgRJGxaNgm3mFM/q1oiy231f+djYca1pgquKF
Asdy0m97tM7BxVWD4DCTnVzW4KbGVodKE/4Ikuj+EFMuWMeRR7pXNrLVsDpUtSTHcFch8CFck364
rXYscS8hs0verH9Syubzq2ovpZQmIgMk8A9KX/dPbaHJEMB9X/e+/Bu4+L6sQkorvDF9nkcUC0kQ
PZLfnUr9ulyQx/UKmeDtUup1Gi9yGq3QbsBQ2qhHpfplTqCIbcT0MZ+zSfokUhqZgxKtYm/ovSfA
n0p0ciNP39lYMj91HgWdG2HJTp9bKM6ZlJ4JiYMZzk47TBtKH9W8VyIcNNNozq9lVB9wkTQF0gKA
qt08KBYsxjMrfKqaln9e5vvaLbCp2t6RMMnp1Uvwfz/F9feZVyndJRgdG4kX1V3pHpwvcjgEEGHg
Uo9VaArSIS45Fz0AyPPdmo6mK8omJiuJ8WU0N2MtnMUlmVZkGzObef0rn4w4bCRXLPNEPL5WzznM
R+8n9XIuInOAgMkNhNxKBbfPp8BITbD3FRjJprMeERQIQE5eeLH/BTbvTiMZoM8soCETBMlT33RW
V8Rlxn82KhlJQ4k3ufdSTyQSWCNQpnNZfMFy+YpRP5JF04QC9ro6mGs+AnNw10R+UgBRXOTRnCIF
bh38RnNod5//NiRAFPH4gOhPXnOhmpk0xFvC5xatKZnpYTyUmLco7mFwWQ0RPGCe7EFHGOwVkCn2
5g+BAc9xUJbuPbth/BjTslpkVrwcL5Ld0u5e5P+Sq/jEyK+L1XzRbs0re4I71VVk974TIwujypU4
Ca/FLn4hebit3FZJabjWFKPtnsdw9X5lbRsvOAKNK615JTIo3nMzmAIPUsNPw9Yj1hTAITIqVsTk
nfaaOB6mUBqKgzCm/xlrTUjzK5qN+7LFarXBnSvAOC04/JIa9znPhTvDVC6R7N5dsxP3WjmeONw1
oDdQkZJ+6AT7vJjWOOg+O8RvVa/S9UH4CPO/aI2axo5HJkNaw4fl5AoM2N3S/uLdgrUlj2BXn/OH
pDv/DY8jtP3/OVBSr81a7eOG18L8F5bD//n2OgP2SZLnGQ5H7SzNExFYKW1DG8ENnKrSyHzOqGv2
R7h1LuCmeHgIDQyJ1pU4gJG90hownFFfbv8ZYxjAMD6zGTPhnYRLxgnOYX0CqI87aK54qYQ6b2a9
OzGK+xsj/Qq+hpzLM2iybwOK7tf6ZhaaonJj/PqcIWpYkYbUFsbKEUC+7UdIaI+QkVVYzP9ohHaq
EHFWAxe7uwzSnlrv4Bgx2l/7lZ3SluNOYFiUlS4Dn0rgPOcIUTq2o18+qxsB9c+Q1l+n7iATggdr
ZXZpLLQAb8ZW5K1jPToaRMjdesuBpdwvX5rvNX+1tq+uJ5wyIqZR2rVoQPw7v+bmNkgkIm9sKBjx
oC/vImLiPPaBVRDH/3S5dRLTv2JBWrEvd5NJlKjLuQ/w7TGETv9p75Ual/XcB7lA9+8BYSrFoX2W
U8i+FI3/TlO01ASPfJvCrTMr47Dn17ewjLr3jFc0TwT0uMbgiSKW6bxawTBp3F1FMiHYJLBk88JK
tc9o8Et7HS3WMu5qyHEvFtiLr+kkjCOWDbPWXHFu5TX1ZP6KtPldmIuJGvoyR8LXUFk0WZqJV481
U4LhHDRX7d8/7R/sUBdkXs6FsbjdZd4EFDkkl6IqVPh2Cl7WYC4FLPhltKJZC5AVh3YGzsgdFDyB
ARUGkz3nXDkXVGHOTJrNy0qqT8F0WChizQF935BZjpgQRXm4D40352THHdJ/5MpdsEGHiqYdIoXH
F/pKaPSMvh44ajwItfafGpS2HZ/U/8eJggb+ZOaDkIBXVeQ3OjHpMFlGnofA8X49nz10dTdlFUEJ
rLjhWAwvNCGh7txjKcCbkLiMtE1imvTNjbht3/wVaVMhAEvLqlf/pSWuOR97ISfhOVWcPXxmUGGY
DO/Zs0aDdDW5/rFRP+ssqZm24m17Z8Nrp7zI6hXi931M+fNlIXoIRa0xMA/uWeVa/zeETg24UiJg
EtzspqcbyE/K2RRPYp3CGK6VF/YwF8aLKEf8lW7C7K6yRwZzE3Aw5ORiN1TtaBkUuoEHKexQG2+v
AgpbIpGrEArbFaDKBYtePNQCoDkUPOI1EyZp3/wmqymDIwGQ5b/Oont3D3ohcDnZ92dwN5svFETW
PgKgKuyq+OJ/BWU/rVYl0YagVPl3kbEQrAaGXe6QfYYSWgNcwzpJGDBogn9HBkCy+6jtrUWxFLYX
O2K7pDIP6TkgAR0CGSzD0IKh2+t1MJtSkRzHIeua87W5eGq2oDxMWGzoVwWLm+vRYUqf4tY2NFhC
PiLXmuEY1lEWcv26J06rujxLKsFMhGjQnZJwbG5bsuMCpOCvgue/SqDIMzo5pqyy1T8cJ0isDC2x
m8kNgAVXL2WsNPAOcTVnccqdIWYq7zO5QbPGgZTkEiMmwOISczKYJK1ya+asbq2UA7SEkdq9L2iq
XesmCwTPgAfYThVobx12U0KxYmMHiX+DuVZst/q0e/F5IiCOCtnrZyQMW+2HgmXjyJiIcwBBZVQc
h9zLRvB4+coYCYJSTSKaAPoMES8LEIK9iuzjddATEm0JVOgW/kQIsep9bcQ2JNhmpK60LylDew9h
sEL22XRjnUgr9oNUEn+DKExwkQZ28O1+nu06auXaZ1jblx0PY0i63h18W8B1GU5U1chamkxL8f5U
4FdJAvTKKgMfR6D31PeSScZLedquLgmD4tG/8I12qONWb24KEWoTVvINlS4JuZ+mYv0XNHvLK8sY
aci3k5+s85efaC/DeHJ6zDgU4f4tkOl9MmFFn1sfkq8LtgesDoC9P+9J/BhhqFsnYhey/AGWDmcC
gM4VXE1USqmuOp7boyZQJ7ifIb+Yoctj6+9kbowEqRdNjRHSjvV490jVZRPd3ou+2SzwlNc7Ruj8
dMWTLWhncsWj2DhJhFM81N7UfGePcyHjwRh1J7bZYPlNKPrQiX/OvS16MFeQ+gPrzl2uYo/iHrNt
ckAB0GH+hf1uIJSpr1IOYpEf+cg+aOz63LqHf87cdTCH8qJsy2x27IoSlGpRpF74QABZAptYL47Q
r/gXhaTbSZl7ABniE5U9NJ6PGbVJLittNO/aqx3QN5N5umiMycmp4cNgQOf8ysdqOqkEisIbmyy9
nudwuzFmtadKCqCfMzlVOksEZ4b03A0ejnJCzJ3b2vqR7Vse00m+7amnZmG1UFR2h5lEe5kiTOcN
Yz2daZ9he2TbfrDj/PLEXLD+nX+VFQdVs/nGRnjSeagLZ3j4xr735furVsUgwp4/1QWHB/JA9ikm
NOm5r2SFrHh1Bp9px+cfLo/PDNJaSDpfc7BEnPRVew76I5v8RifnSpqtIX7dAf5HzOqXu9fZOEcF
+DgW5b0IL+q56K0VUEg6+dEqjUZZtaQ2eaMje6KbE+feOcvfDJqYk7seLnTNCJtXB8p/JYuVk1uv
+Ja5zH8MRhgCup4nS5p38GXak1s7xJc40jVbiolLjJwQm9NmXgAe5y4p2oo4CFtp7YQDx7pK6gD8
q60SbO82RiyK+/oyD7etdes0HWPE8VGjXtIr/fSpcXP9hijd0ukK/tkdO9+f1p3tLNMCqOs/JYKq
76FFj23iZYSIZp5EJmIx8ntcsxDcIltq/tiesPjKbWZTdyuO6uDro72O8ChuyYlE4WUlEIJqW750
DP8QtfXaJpAn0tj96i5FS522mJlxPbkbOQNhtPoH4w/fcQ5lzDvuHJztVjNwtZX4rapaJIxe+R8D
Hp/IFgb/tZ2DRmbNKJxUCW6Til/PUy+Y+HPRyTHPycU6kIa+34qqY+sBPJQlXlFXRPVYdAr1+lVV
aWry0J9zQYFad/GCR6WVQT2BIVS9HstPDxLFsmipQRvy/Gqf55j8WbjlYacZRSPmozGcRQ6YYb6R
0MdRxBj1lEDY8jkRcFBVfWW/CJCQH11BBs/lB0DcLQigpXm3A5o1pLYdy+7KsLcxJDi2BOA26WMK
5nI/d5hvBRwmzyvR4jw6r/yDvgvDcBJfxOYvcix4lS9EZc5BwaCN/VffYlVQ4td7rTQL6vafbCSy
WhorKHle5mNk8Ox2kfkflVBc/BT4jfq4kBfjrdqMYC3F9f0NZOlbJl4smA15A0fPK3aYKV4MwmGv
XXbRRQSeFP5dbpy8ETJmptIGgW6Vcl62R9nbfjMTnhF/p146m6epxZCl5FL0/w0VVFc2Q4NPF3Mc
5QQ6AWfAg+JpaV2F61VURqA65+pWyEpPyXn3aVOF+LgTX8RoE6SHtQ9xJ61sG8FylCgdbEl8BGyQ
thqVeEXgTjT2CPmVNw7Y7b+6Fbx03z6hM/DnFQAziS8LLHbyMf3HJ6ZaxhxcfU33G8ZHKtXxVwWB
FmExwznyGeU+C+0B2vwZRWrdiTlReY+D4t+KSbmTf0j2X9DVZXItw5ULiD3+DBcALR6zeC+BOQKe
PjdYscTfNfDquMZafRfCMYt4hTQZBcAYLfFUbScBc3L7zFAtcbuHoUMh34iry/wMeLqmwnoa7pdO
jaZhFKE/vDWxHi2AQemgXGDbUlr+YBkAueRdDiJMRp3zfEz3gkOInz5qOCtABQXpBEmNRk/DSPOL
HZY2jIF9p76+j8BDTsPtjjmmevQkbDIggvruTmWG+ym4w6tpmVKQqmQs0xQ1+m41DMpzPVd5tuE9
tGRq2GlR6KraSc/dMuRsIAlFP+2a1+7KRStmYDLgtCCK969ryKvRJWPNeneASkjCD9I8qQsnxxK5
9ElMMk7FW1oH70zEShgkd49oJjgWR1gGb8h+1uBi7eirDOvLlo9OCUQ875LPHdrtmh4INcM9jRQq
75IO+V/e/E/MkO14N0JVrjMyiUQ8UQbe3LqBuL9GuLgyZLWRw/lf1G4qlCICxcdy4VCCzRYTdZkr
L+itv4YJsuG7boHSoRKWbdKSQ1bR5wGk9V5MH4h9eV/16eS/F0OBEQeBZuuf33j6LPckbhzVfl7P
aDYzPzszG5msJIYxLta3bb+Mf+vKFU3CkRblHKWLeOLJgDK4qUJL1L10rQqxsJyc+LfnurY1iRXG
B/OY+JNWs8k2coNSP3Bv3ApPSeDJswRSgjSeUoTMFPCf10q2Ewn/kZLad0OYft4o0uGG9eLA0g0t
humsKxd5fdRJJcEa2rynf7GdrYbGXa5/JnxPgHsmm6PgerL06stXwkzebhWp2tqqUTAN328I/DQI
af16VGJOc8+2IlBiCkUf7lPllDkl3fONL95rFHTuVZCKb9npWhtESb7Ds4P6wz9tp0f7FI8MJARA
O8Rw8C6rQLdpYpv7gxuC8Kg8gUOVwlA8CiRXGf/n4/Mf0JJxzkm1iARj7SHWm9ZPKMu9yhA4v7cI
L+AU5HJjpt6WdB8NFQh0mbqnbiuv3UgWWdpJg5cI8pauTxWXmcPu+O9R8D/KO3frB0Fh8CPwGZxW
8nLsG932+guEfin1gN9PhXse0cdT+Ax/lZrXGq6/tubE0UhmFpjyrn0y+F5PR0YZcoihBzwDObno
vgqAQIFAQfehkTJ7APZJ+R4wQqP6nyNry79XVmF3SAG6WqxA8LGDAV4Vr09cw2olwy56I5XjEvm3
LISgGQ/UU2BmS0kyW1oBFI6/R3LetPJRS5g/ElL/4E8hsANJffDjrnXhBIsWbSwzzA1TZpUBjgCs
mKOVC7JWcQp12rIz1GDT7a10SRB/EaJuVozObQ2BonJOaOc2WJVBIcQA5rk9L57hjmnvVTf84VR5
3OWzyEZhFZdd92KEjt8ykkYlRWHPoyjjCkEz/xC9NdyYmWNIbP4TwyITkp8XV7yhDL6ZxHo/rvh8
hks7e67WArLg5zveu1pN5AvlJPCBTjQbp3Kv5N2n3RqBVLhye95lEA03d8H8QU6qFkk3Ii2owLy4
XNGFMqJFcdAzVG1CDr96PiUKnUitpl+RNBOn+F7PxNT/WBZayPzGhPZ0DWdb/NWYyLI1L5pd0594
XISrhmT+ZO+n0QgpTDwK3gSeeTMazJmJckzWOfuJ8RehqhIGMJIs4WV1ljd0mP4u+RYKorvZnsXv
c5MyHmOiP3crHymgHyBARIT92Lz5hdW2HKomlhHN58mLxd7v8YSaFN3KiTvqU6I7dvY7kX4UnYzw
snxF6zLLYvWsb8QJx3MHsKQFOo3w4lhRr3gu3qUTycIzS4jfE5v9ztVo7L2gcdFG/nhxwhaBMnjS
fRtOASjfVoiPh7Ut8JJ4kxhghg23UeC9O87RuK1GDlvMEIyktamGr55D2N3Duxjfj03sAENhTSjZ
VUeicAS6xURS8vGBygatmkBV8g9t1QSoq3pXa9sS2eqFQ5BLeiQfJzakO4NSybZkIWw8bRvXf68f
PXvB+pnbAwYkxwLY2NgmvFBl3gneQ0KlrSjBSR6QLRL+aKXNFx8srrUXXcZuTzIluAu4Eu/epQEd
TcgBw53VJ44OoslVdGNFYluFQENFx2cR0vqwcEROpQPkrX+FmgqRbmAErgn/NZIV+onxGnKxD4zJ
91riAX3Z2zrABEnu0AfXACFUwlDgx+7JJNWhsTv7PsWTW8Zws8GKZnMteb3sdS5wTdMQa4LcmlAD
dPOtAYRbmsfFk1fuEFckv9saKWVpSbwue0SNtDBVgQHKsNnkeJm6KKnBQ7o3JfJXK2Jt/OHdmFsK
e+GUIQhyRPEbpwndKZ89zUFKq64tFt8CtOYmdS7h/VLx2MPUhPSBu4/Lkg6PH2KhrTVqiIZXC3Y8
h04yiLxo1/QXbIZrgJVGGfcdKMDKUsQtYmtqB2Fgo6sU7suatCjtBzMojS978SRhBiqX7J6gBrct
dowm6/9iE0VMH1hQawuuXU6HtKxOKKnKkEkV65J7HZDLXv6S7BuFCIU1n4iLUvyNPDPN6HNSDh0d
ah7HxHkpbeIvy9hanKDQSWNx23HJHR7njb2lcSACk/rPK6Zvcqsw7XAwIuYlTicZ1ZRF50Oo6gLC
9mV+GXjtyBwEHcQaPE4yVku1ZAN8oHEYp5ApaiA6svo0/uPdrZFkKl+g/Ybj2V9lhvOzFPUNNOY3
V78CuaL4LRMVwVkSEA39u9IXeVbozTt2wF9cYAlGI2V2afyrv6cnb1QFB6/MK2A2gD7QOU/2TLuy
/AruKktYgDenPAgx8//6uH7bHZSOLTGi9bz9og4Re2blsREKaMMQ0yJTp8Q9dD24Gh3kiYVN+A/e
U3HxGSKaZEeqq48mdYfiN+/wRfeu0Ehup+Ap/uwLQ5cI0qyl4JilMoK902np/3BYUEarDtyWIOd1
jHH3d1fbhLz8H+BB6hbs+RWIfGS2q0JtC8b9MXcGwPQ2lAIgws9GVWyFMeZZmKgvijauXpE1Zs/U
aRw8BkUY/dZQ78XnXgveQjScF/GRI7Vo4sRgQY+KYD4JFx+og/XoLBu/P39p67xfMF85f6YifE1V
qDrZsrkWkLgO5b9US+HdW9LbYO4SKy5ApKwHXz0ZT95qwXljlgG5320BdvUECARG9D8ESUqcLGBW
XmacMqc56AvW418K9piMqR0PFx9u2mGdM6KcjwZ3YSnC6+yddjuy0DO26WIXAfUsB4aeybX4tTBz
ijI+3x2E9dVN4GMs91mC/S2sN72N3zj7j8foNXEy2fl7WFfUzKtYx6Ek+RdJngUnMXfNHcGSbxAf
H264wV1SWbevX9qk8jF6gJH7G3HMFEXXfmiTel1EWRt8XhvPInUg6Cezooxk3A4uLAVcAng0wTTA
EMyOl9v5JJMZnaDSTDTdxaHxEY2g3MVRbgtLacEjLs0QOcPWHz8OMOzLlGAZxjxMYUZ/5sjMFgHr
3GhqMzTzpIR2UeHmmgGi3kuMvMYhUp0q5EsBWTSxovZqRNO7FFkf2USy6dZ//bNAfOTVN9vGkFJK
4SeLUY9w3Vs11KVIsmfl6as32xuwQnsFxpujWrNs40HIz8EMGSH039zSIwkvBWZM29gVHU9F/njD
X5/ntuRK8Ab64xS4NBJAS16ZRxTphT9QG/koNPB8XFFpQxvYt/tTRCkdxADzJK7ZHJO8DnjFO1IU
40CqWLLvrK5sOMXvpQGN9Cv8utC0pqY5AigjaP/Ez2u3X6Q0aK900DAf49ava8NekLTkiv+QqnIu
/Rm3mh53DBuWW+nlFZQmCeDUDBveCQnWvtrUCsTPmk35XTB1oHY6numT/XMP9SRo/mhChisYPgzX
1WvudVxjPvwz9gUwbXtEZ8NIdvgtZsS4D+U8PnGgE3YdqkaqyVAmFm4kzlX7ZRkpWVqCizDOwLv2
tH+T7op3zJdOEiikik7dLFpDkxtQJxc7o4IrpP5NNJL1fUp0WHV4rB5oOncUFhLp7dQArLWrgtiB
zf9KeNglyvFGEAkNEPuV2PMjYxc/hCas3dGjQT+4zDY52zBDTOGmZBxSZyACrRBJAtLc002NlnQc
XLa7tNvxB9KKz6jfa2WdBKg67TAI7/wV/1UBxNXSgZtnj0XMZIlq8uc5vvL1DtSQJA3bhhf+GtAo
66Cz1B/EZTtfzIigW0OF84c6jB/JeyVNtMcPwcnertIfs3EMxBWv+3jV/01zbX4XTT+0HKCyf6MG
Iz+nQN7CV4n0C7YWSQ73/iMMUe4pSDAefZrzo8CI6Urr1gOeNCq7lytHYZ97w7fIj5Hjj5IeBnBk
xZHDFHRi5o3x1B5WZuGQ1QDnOGXfLzzk5EN+EWqxxlTp78X209bi6nWo/WSj7UxO9wApp1VTskaZ
SIXnsp/nEDXWMdvtMtVi7d7Gc2++R2T6qtSLqEtVWn50gVogXY0rLkisyKnHEZQRTj0w1Qt5a1Dr
9du5gHaKoAi1QyobhCY3toiLmVCVbEPAJgKnfLN5sybQ6VBdByPtX8/j4EatNxfahGOQpdjwKkg3
dXjtnVYew5P9/9zUGVhHRyRaxs50UYCLLcDynBnQ6LPWPn8pjZMCX02yDfsqWyv1OP9KS0aN88Ay
a9fieQx4N34HPAnqJjeaUaXrA+i1bk3TjYEBu/WBkVtqkuQFqF53KCRsO3eHIw67pLyjtiH2ZP5o
uo8g1d+QZqGcmbk8rZML/yGqvQ6XsR/9GhG98KpkONNbgI51NK8UDRatNvf/ES7ayuZ6UGIuA9dn
0mA1H+EF8iOByKUzJyXnaIA2b82jm21FUu3i0lWz5/ZRbK3t37iZmeGmIJQsmN6naki3yRupYxib
Fsz3ymFVVOz4/xdd5AhFDdUA1xMBb0j4H0eWWsRJzXb+KYjyzDVquu2N/VodnPISc0tqhk3rMuUV
ecPgu2WxmweN0xqRwF1aMqC7BXPOlKJQMtAV895tY/J5HTAQ19pOONHettZ9L0NFVk+rn9V4HBQc
a+B8bRIKSnr8codjs81EJ4xlJNymh5XKlCBh+nXFTzsZ1VLk4Y08VSDznjjfo4WbFe9f7Q0iIsuB
RAsxPMYfustymz5tGt4BjfiYz0O3AjdpQBx+NrrB8x1rwXqVdiox4VA4sivvMSFatzjX+YHVfOdT
oV44cCsWCxlAcwtYPzcRWg5TOktA6XBKgup4I1ndb55q8J6JOvsrsTqzxbpS48O5fFk6krGzN/7b
hxP2dhefzKksnwf1lLf1HDh3J+x/eyvCMx5y8Y3VmeocFNiCYSJ3UChvdOOFWQXLte3EhPw1ztoZ
iPPhrQ653ltYW/k6t69rKuy47kp8QEtC9AkCo1SPaa0E+KgfFLgDhzZ5vsf+mVi8jGawATB0SRNQ
WQ+mUNxN1QQrap+xDYUyCGU7xF/xvHLaP+WZuZlEGYIBCByq2++2vZb9xReGBQj4HkCSq7GKqjO8
mI44Xomb9zAJxQ/xcylpkZeXkUjLtvWuYsO/dkRnjGkYsPVjLUCV55efZuq4mXOCTepEtHzlHUuw
cEaATlnub1FFxK6PYOcK9y/pts0p5jOqSH3cckewkewM0VgJQJUP932xQMlcI/aIBau1wKp+hvaF
KiOf1D3YB+OqXT4Up4culW/g62E2ckXGnN9kNDCuBd++8Vdps2kS0LOt5FOkWRrNVdiTlMrviWvU
6zXbCKy0o2kSyPzhzD1qD+RMpDB+zmUqeb6tYiAeLo60gRp5f9T3+Tj/hE48jaPZ8zkFHfiLz9DA
K2tfbxOgnnXYeJUM/9A5uL5BgzwwgjK/q4++/YpIqsTt3iu3LNMXnBj0pJSz27ZvO7bxR/FP0oaA
4Ccp2b8beBPEEN0XzTxBnPIcD9O+e0roOwR7Wu7eJ8nIPy4CemwPMVoD3E8QrMX+yImycMb2yuov
UonK4rMpZi+4BrzqWUQ9lTIoNnjmUhhYxUUu0MZzgUpaTSDHKFuxtarx9SXww1omMs0meKVwp/rB
dXUo9TW8ed9NEZBiOMc13a9PAHWSNj0pSle4hqy9kaO69qe8wxdtCkG+0OdNAqLeADzYULdV3LZd
YtXY5+SLXVIVvdT4UezK94q3/PxiWa4VqQlWQCjjDjUxdws9yLRXSG8HsfBJOI/lq9HSN0RjDpwU
q27gXqb1KtMH2pykVHCyyodf/1rw0drbvrBWPMiArNpTGEs6elyXQhDt9e6gGa/nCaVLuk3C9fJl
Iw5TaysIggXPq+ekE9TjmB04iBouOznMaaSrUDPAY+x4bTlFVC98O7veJ7JqiGMnunT6wN466xlL
LEP5dQf8mk5UkSq/bxwNMxpUhSSAAdpVwI9r44wJ3Y338FpngnjmZCAl0V7pmXriYTFLtdcNcNec
VPYYU83MESHn0IlUTsTLtOvJHjaQRNzCnz36JLkwg8JcqgD2ZL6A0xvY98XbFefQdnN69MqmFnST
xovEYI0Gf2WrjU7ltzvpQeFytdc3UOnmjaLUnmTUt9M1qrreWDtGgla9lyQjjHDx/biYa/A454Cq
dC1L2FyZNGpdcyqj+bePYw0zc4Md0nyOEZtoEh8Tq4vuQD4mk1S4U5ALH5KMtOzpHqXxYVrd7u+d
yKkgIVjiJw5dn8gtu+MvKURCNatUoCqLsWRXwp+VrzTrLx9kl25hvVDzWoDPpHk5AkJMiXiU+enO
p0moRCmqtFFbGFA9NfRdJD1aVOiZVEty+R6ye/efLJX4kilrVxJlbzMTSD6pXSbtbe5OMFrHH2ol
fCVv2sw7OzXTBOP6KMApxwXUjpV/hipm94Ey8LY3ZZ6llk7sFaDYXlVVi7pMG32Gx9EQ5UlXTJoV
YleT4bRo0MOD6EaJ2KanVsgebae20jKTAfdx4mMoXkmWXtgN6RMQq60eJvoor83Nwd5xN8cZ8mqz
CPbyguF8F4EIHA5X/sTGmlLIpqZiVCgUWJvB68fsH6jtPBP89eaVXt2ezv8V145iksLXQR6dpz34
J1fG6bJam8bsonnd00+i61h28SH+26/V3gLLDc9wTbixVHFoVmLTjFLiUr43GqASsGdPiFTNZCB4
HIXubRy4qVUfmApvsoWnh2zN2I6+cMv++aaVIBM0Upx1h6TtEVcAXV7lm4Gg1JMQoC5h41S+bU4y
/UlZF7nwJJKiQiODlZLaSU/su0//0WLxNgh9e8zx7cu3Y/LTE06jtUDt3HOfEaKMLktiwNXaRaEK
ZmosFDv/zgKx0IhwwrpMzFpTAuX+qP/p9vwQs7LhW5zwYHoC3Rk7FS/+Jeqwic0NvZtFypWH+On/
epqh3tSbaNz0vTq9Z8Gw0kliUBPl/ikqoBSNulxOCokH5JrtmhbcjuWjlVI4O9nGhiWwkOVYwdra
I79KjHzXCajvlTnkBdO1DWFnYNKVp5cEFn2WpvEJeqHFnmEybaBTDyu0ETJVnJwCKV/EeBQSlbhL
ud4/PT8dq7q1e/ieMgquWkYyvDSmT57aoesqejLP4GpFACVo/e/ciu2u8OEKApHRMSzPovpQ53WK
J8O+2XWA9c+BtZxObzqP09fBc+HUGAjqNbjF1HkU/eKtWpS8Jyq8N0FEq3uqg+gKgiLnijbXEoQK
rJW/dzNdE3rJ8xbMEF9iZEVfYGDz3wnkH/6u3kJP+q7PKOFJqJcU7Ia647d9CLQ8BywgknOL9xeY
rVCUzf6WKokQOQWKR7xtAXEp/4onIdO+vfemhlPh74sOwB9u6Cgg8lTuoOwGecaZ456iiF9cz9dP
wDD+Uxl6Rn9LU053WuXxhGAtyTizfiGac2EUHU/4UgrcoEZS6+N/wmMQHKmb/u7CQe7wskoBNbiZ
prMpRYkzt8ETx/A5t/z2F72PCrsnlB6GHDAyiMklBourEQ93tq6qXNaiGVL3p91cX5f35s+nk/9j
ct7/teTXdRqYqjTSaun6DvjczShDN8JUt/I5pd+fcAyISGL2Xp3Oo59mMnRHrOMe2QQi6EzbkTRq
t2Uzg6mVhO1CmC95blSbPLIdcheValoi4GvoKZGDi4M/N4HQEzDbaP1UmvYIBAJCfx6WjM1nloI+
noHYJlxpEXUdftv4eu+Y0y7BXnWQqaxbueifTedtDpACrEhu948X9wfEQY5vWsjDN3Bdzs1jxrT1
/kag41j7SWtxhUYFQUjHIEzIQ89aA9udXTbx8KSXu00IN2V3kf1Rfd0KMaXICOkvq0UO7eJJuZQh
12yc557evvS/CpD7DpfZRf5suF6KqnQMTLQynAmXxCuoq5c3RPttKxzB35k+pTrJsPIJi+2B5GWU
pMyBt4BCOXiLhCWB5lO8GAfvj1qRQnn075/NZLBq9uZulWQNIOlho6yTWcvjQzyaImqGecc7Ub1s
MO8uD9q9c/mNqdGVOvgh2VBIEl1WRrdvh8T8CIdYhWVEGHBXtoVOpFWevWpHEF9grBYmQi1ebIjt
deWLQS4kTOMb5F/bXqp2kiEp9FsXdSmtIgjNzIxHAmSEgT3xdRNJ8EPrUOdXfaPeXQ8QWoWVm5Cf
lVz8p36Lmm6wLJdMWm+ZqQ83Zs/YG88GvfJ3ltLoS+B3yI538iSLLZswjDtqsGtihFZQxUk4eQM1
akVSY/PT4RSxckxl/ZcBBeSlNacaYQ93hzC/O2YXdKek7vxj/82uPOm22Gut+gh5wFrdW+HboAe0
ISMu7Ex1CCUBq0kE5c6e4+Smh4g9xbdLOuJt0pxyQX65Jg6Xsw2CNOFALeZOROZ6RfANFC01Cfia
1Ys1b9PijbyswJ5iErelZzUAH9izGf1fj5nez60ElqX7islBN6Akp3+akZqDI8lBULsOA9j7i3c4
VikDGkNqZJs69wnGhxGbON65oHJ5+r79DztyZZc1nWDUN68cDLC5tZTYBZyIJ9xkr3NNrKaOTvRX
BKG0dnh7Pvh1hfE4tKnYzM3ZMkDvuoDrAlEmfa1riJGmllg66X/056Kl7z1UhMXAVcYDl/epgnxK
2CGkpk5fweXMLDPp9HPSTK7WZDX0W/S3YLyqFzCJvkYqoTWGB34QFUhvXyUR3QV7kI7YTFsG8oRV
c6ouXVkhxk7RoHhxHWjtX/STgi2mMeu9hARCWGMg0t8GSHkBVmetS24PYelW5Y/QvB6msQQaXbSs
zY+IG14B9yzeGh0lxcqK5Qk7+rOVwpzGivDtwEZrnAciFqo6Jdip4QC7o7cz1hCo3nptUqpAiyeZ
DtKCaapA9IyBskt+5VzJD4UUAOcy+1GkUHnt81V6jgQVcwuQb5EVBjL40z581ZTLojA7Z1PnxTcR
BKkquD6LVJCJVYy7aR8Vi4+CgfjItGckXf3Y5IaCKHPiKlLC7GJQOpyJ7UOMmqjqGWzqSkcSU9D3
KIOvhQXprB/Nx/ddNtTb4PKCWY7UQlGATsmGEL66Dxq1YIai32ogdzTiWNl/2R6edOPXy68xjIUv
GP/VuzJF127dXGvYnKlav+EyIaeUTPlabGcsmJiHFN2dzLgP4pgZZ0EAE0JDWbB6hyFlLAQv397i
F2Wh4YeQnMJrVaFMHefrZvUiKZGFLCw9wbGEXII7oHRoZ4iEif1C4Dme3ogWq+uuBcpPdmak9Dqy
ZZU0JZBq3UOJ++VsJfCAE0oO22ORu+zJPQq+pIPVgKisoK/lEGMWhUHgE3SQNTNrJEFP6KNj51mW
uyIfEUs9Fn6tobXR31wkWsfZwhzc+W6dMvMV28WohpO79ZiVzr9wZy7ZvmfwYBQhi6ZQZZbfsS2J
mUmSBgvor5Dar3D86zh+NGbbsqZKYwmkCctLlpPNueoVEc1Rjmf7KsdJUHfQ7f3ghKDlyVdDwy6B
K4bjkwB6JzI0cgtIbMpib/y8Uafj4NGP0HhL7g7ao4nipb9R6wqA7ECp/iXmbiKTG+42064YLe4u
Tr8vrSmu3jkT9ZjAspTeuIngffaoKWuI/pAvVIJixf8goo5cnwPsgIII4OVPHvfCTZRzSQXSXaZO
5bT0b71Dg52MFZCn3sIpQlHc02LYcYoO35t4ahJHqJhwNHHcNS++GS1em1gE+7PjK97BGyxn+iif
NJzfVM6kLicoXUcp8AV4QjlKXuv8owB6n6TSfL9+5hWTb00Qsev8b0RLcXdBjIxf2CG7xnANJOHr
ePxBQroNJkBy5ItFrzetpMQ9v6IC2xGJl46j0C3oPHYpYhvKVNTpyolGZyjG5qdnVRhttOWSukpl
pOeBANvtocOHJ/B9xWwZMAsLp7HivgB8aCDdTGNPea+Ingky7Ps2UZ/fhsZhEJSJEHh5kd/g5uIL
c/XTX6O5uZ/bgGBsih9g7pcNO+xmAcK3/kbcAT6ywcFu9SVvbWS02dVUnXEzcz+sJ2+MyrIep3ub
qGO/uWZC0FCo2ojocDMaiKYMQdoBu8RdzxV50b12lnDJCMJpKEVa4hmdoTAfmN13ylWqLfgelwOK
l+8tu4bYvZk8aTscFo5lWmaQE7MQxgFYjKzeNMXL1Qo6wVaT1bXf6OE6raUYwnsL8dfAbmrmySaZ
WG3K+ioIfOGWy0xYW6ZI+FCartONjAVG3pzU/TJ3N6qzP9TpmAbuXjcAVP6UDzY71CZWM9XytCzC
5ioq+P6BTstBeTuNUxMTtlQc3nfeI8j5FAEf3hJSAyQrJFXNr3YHJdBNB6c+Hmo6oevVTqpkfxKQ
SQZmK5S3h6fSemJykTZFd0Xz98v64Aox5i8MUUf9F9hxJJfWR8w+u9f001+CEQUEN2o/hFQWdVBp
3rA7oAwReis9JfV1d0E9W1/BPKt/n8iAHpDyiVzmoxJNhDY1Bjw8Vuk9rYi5aZeQvkGjXsvEgE1D
QESkjwqao2Dm3OUZ620I3yvkGaKnpec83GchhxWcWb2wL+T1tpJmM0aJUjZU7WyEgzBjLNBNfV9q
dNLSirHvsfIhI0TkaE8Fw1HHEu1ToBPOu8ZdUyjFvya89dyYhrlyZi4s/DUbfJDNLmP/DH7ItHNd
Iv/RvJ//+orZvAhkrOcw3IVmCVj9oukv3OV2BJOHPvDJKhIARg5T2mpkiMUIQZi5Cp+M6hth2Vr8
bHpp6BNYAvk+BVjAQcsv8gvUUVLIT9QDYHglca6N/rzf8ZgsxRNihbu4v/a6NX7YIWeumAZVHc+v
DYe8xIWdU5+aCG9r3D9gzgKXmKm7gQ9Gu5RJUFHq7rW86Ffuf1WVfzmtvhoEO+BSp2I+9yDqxKdk
JK4TXIY3ui9QLipGMXEXPwvH97c0FgaGchVhBoP8NrF6nz6sz503JXl8uDBhx7lHSBomNakPpdhL
RsU5Zbgs7iL6+M8uHmwcha5rF/Aa2yyJRtrLsiP/JxVqypF+EYhpR9dR0j5OOlNKHiTPbfLAX2/n
NUsWiXgfB09gEaCP4J7jiUpK32pRgSYgSOEs3XlFBujrb6ZzZMxn/rKPuSagkS6U+EE/GiD/AZ34
UV3/ORbPUC05GVUn2JFuhcjUM295tSvaASdJsuCTAG0UpPx5gEBNwGC8rtz093CTYCmpTMz4RNZh
czFiIUcnMtiuk/x2nosdHO73cBCPrV6xJzybfGWkvPsxSjaTRg062iAHEE727D36M3/YFMCbmlqE
KpoxT48zv3jjedI2PAr+32Oaw3UpqWTopQox2ZQMg9bUCGbI8fXssU468dzDbiYDSedc7maZZl5h
yWppEI/EpwVIWb+JYBwmXJSshqnjchvxGCE3V3Xmh/p6BLccloBynaBkf4txeq43TKYS9JutXxCa
immf72dgyGnBVIu1vrQaCKYZ+ANkxbETTz3ack5Tf3JBA8g33R0Iy0Z2M5RS7YbTlS4Rq38DRPdA
XOJJkxZkCf9vEFi9AFsLEa9TEY1ychANIvBDfhu/FYeVGhXxbd0o60/zC28c9HcIhrXqUWlaUbww
8cq4VRj4rASu+WwaVUuUi9o48sbNxwpJf46Tq9NT/T3Rsz2Qe2HdFmQ52Kcv4eGACrqYmmypDPnN
kwfCurq6ZyeLv5Zqj/nc1KVO+rXCKug7O0XJ1c3bsUI+R7dF1oKIa2jRIiIeFfNoN4d9CCa19W6v
/0FHS2yPcCCJ/1J5/GUu3jizau2gs+cgjnqnqbQf/tlHbAfzJ8O1manekFwPfGsTc4KEoII5JaBQ
GjeCJS7OTkNRr3yeMpD/0JvXW07Bqz/YXlC4BlJeI3dHR+50bwzuPjxk9H4vxR053YVzggtVuKX3
fXL2Rq8EbJDqg44vnQxPe4w5NZjjp7FttGp4yNpMGsV019lcScJjNVGJnOqOtAe4Ag08u65zqLJB
vwzBC1icC7snClf1U84omptbXub2X+uUixIH8SxSvWSuzzM7NMrbvdSgD0saqx3Yd1fyXf9Yj0Kh
cOLAdIy+UTqYE9vUOaSmQo1n6S0RLMmfc5yGtdaHa6DiYIEW8Y4xG/LWxGW1APVkyCl8MIaviK9h
uAvedI3x8inN0zE+BnwYYBRQUjr4hu3VfzKJtHOeYnRNl58cZPSOn9b/JN7oZt9TCI8S7NpmZMzz
0OtBzPq24HhGSsBjD7jbKmcmOPYkj9DDWzoR+PhuPT95vGj5p7shxq+jI4EozSlIarWelmKORthG
qTY4vUTZDFF9zv2dheYAtjV4VLK/KTvz9L25dNHfCwI2PfdGpmFUczcaqhewEtGv4N5k8yCZbwJn
WZSdnJtRt3rdNKZhnGXisMZV7e0dKxo/c74/tAWZvoP59v/W7phCJ+ir+rhr63caSh+5ShEqE6Bv
/S8ImcMmcvLRuK6/QzXi6ndc/G99mbtODuZFHkTN6vJhgDoity+XBBANfpf9UQbi/aorKH1urNyT
//AqXX3OJankPDAhml2iHupBwuNvM8fXT4Yn3DwCyurBMwVQhNP1dey4iu1iRh21dUEAgH1ZiwVM
ayN1JnsynDHKbFezUg8T5t86LK7mr7/uK3Bdm/2sSJAaXclvdW9sfqfkX5xEBJlTTNeLQloPAC3G
KkXhtQcXuwB6+GSae6iph8dfgzwJKhFTQCOVYqL8T2JrOLno8721O2y95ygqd5ta5CQxyl3xG2y/
jLXeAEPsJO+9OltvO9Dde8pS3bNkDT3hdy7WolP+1ajoT6LNbK9D4G2F5YbzZw0/aMm0feqMYZ/H
4M2Lh6dZ0AAkKKQr2lMO3CCrgPB3315UlMw5ortB1LL+yCktwmuYdqqvNdVtTsjCeYX7341M5Uhq
+6mo+aE7ygMVoDpyURiljWzwnqBErCphV9GhCWPDs0XExMOQr+CzLrDS6AN0gufy4/y+J4PBOPN7
PWEVTTgf+KSNUiqUzrJfAuL55Tx+iCn02Hh9lr+1jGTySY2nSxzHJIg4vw3rMgkfJ42np2Gf9xt2
ZXIoZZGxgZw1RLhlDwXNxtTa9VhsjhdygDbKk9MHjiXncGECq4kEjbO5Ugj5lQFx2MI2N3Q92vFE
IWa0EMgAGGXs7cuaz3+VlLxQIFeXZA9qRxKND81+N0NyBhf/duPbv5uJ3BlqBHuZWsPAl8SdfNUF
8j1a96Z6ebQx1y7U7ji7uv2yHCRbdro03NjoF9rsfvDuqLFNdfOUXI8E+oXB4mJH+9E4KmIqciea
Zc+1ZQORpcdRdXjUDMGqU3+SyttiipI2XUVWh+OlcIxDSm8cCa3rlvvkdwsBkpkscNdmtPF5pw2r
xqH3nVWlLOWLM00QQ04BWQZ0CnY9Ac4ErLwX/Y9k6bYvwPLiENTsvFe3IK2nQ2lbBY+472F6stF9
OlYs28bBwjm2hXWM7IEhEwivN/Yghgen88a0j7/wO2i0pMoa/Bzgeiq4NzPEB3CGsjBu66IpI74v
rvzVs2QMZ/zVosYQT19WVSfPNDJ5tIxWd0NBpt+5QJ3CGPHw3lSv3oUs5wWQnp3z40eB+Hv0TUhX
wxtH0VaF2loIPt5+Sx+ke6pGU3Q7U7xBH+DJTdAVJYj1wj+EYi++SMQHlscDA/7zqfvKggEg1YML
ZwfIpr4dYAm94qsqYdgtL1FeFQSmVHjmUJDDFanZ/YaumHbsu0XeoTP6yHOK/7FJqeEyzbEyJQR/
630EpqHan5LCTHB9DErVvD3E6vMXSumqA9LL1Gqm2Pm0Kka7zTUWqw6C/YNoFQC9iolur9NA31Ap
Xo6XaxLVY+hqE553I1iAZ9U+5pW3yoaeQJ1t+i2qProj4fLqwmh/ujh+9m4jSPZq93XigKYN2xEP
4q2pj6SXY9Xv9nciETH7EHmKaTyw1opz0rdGNXSwVB1Ko2DwJ1MgCIHli/OHaWqBr1ngHSirzRNq
TegiSzSUMYG+tHmxevJkdQtY7JKT2YVUiuAT1Mls7Ze9/aYKgUr7rd1X1uExrFmkZzbqtHfaBrZk
Tc4DxcCuYpkkdJyY4T+seP+g810QDSHaKWtEqRcXCVuEqQ8FgwJdx+JDOzAMO/UL/p9gO5kFsYIf
Ia9A3LFclyS/8KCZYuM0YCRwiiot7dNcHDd2sMbw6Bpp5ia41H7iRaZIT4sZ53FoKL7WW4/oHwPY
qkEPnVwcWJiMXit2XWjl9tezTRa+lcusrVbP9RuQlG8TLll16MvW6AqmhQ7kAAqCcnACj0MDx4JI
rd53Iu50bfXji9dsh8ODB+EpBWajf+l3pPVE0LVKlRkc1biBRCvDkJQLr3+/DX/Xcsi3kp/uSFbj
/7n8wL0Bjjuv3dz5usJyv09a4bD3vrQuA7UkP4n8NjsgyL51i5r/GsdeI9CiZSBU2Gxr2AagKFmZ
WUd7lnx+kU1uhoXVBGHco9D3gIuxMVMMdfgoVxPCU28eSIRcTUFnE4aPsLvIz8QJN9rnmMDFCQwo
frQuduLnDVoWSu8Gaj2JyISvg13/35QJ9ECn6rgQdYQuDF6CecwmY8lFXJQTIcBREXmBy2pxV8hI
UVKLI0WuYYBa9G7+s9fivDxv+BqXz0/ML4HR5p6Vw3Ha52vQyL1SeNF4wsgC+dF66rugDeGvvbVo
OlQVhCQLOtt3eDOdpsaB+q94IVBXl1frSgLAjMYF26Z3sxW6fGCRGQK1e63ro4sIVuMXVNWW6+B5
qppPKucmivjHzcBnsNexGeC1tbZgXzwqdA3KPp5467Ho7+PZjf4qjpWkWqlupyhn+xl2a8MMCjgU
fwTdLjcB0/ko3ekV8hkYU5JCtVjuUcBIy0ED/OvzV3a0foKEDZ3+CpJf89VCVljijejfBRTa7gk1
nd2aIL0XnMt1bLxTtHzvyXhtTBMHSMFpUWqBZCa5LVJps7NrVSZWHhiJXILelT3nuRnVyK6vSOL/
/HojrgyBTw7JeKFVfPNQtCq1Evt0esD0SJSf9q8sVRGq0AgM+8wHKvyh7yTP8jSzE1eZJdxdR9Yb
edGPErH5HZy28L9GQPxyRPuRV/Yy+pIji9sf+49iBZp0Xuz/Fq21Q164sCH6J1Wi/HS5fFTrwi27
T7mE/h/N1NEwC2g+FGXzv/3nevbFCCo/1jOYjLeCoAU60L+0824d5JVdBqj/UOq5qrrPGyWmU7HG
bIgwy1mOvnolZEZi+aFnsMXwgeUQl88otXUBSl9nK/Y943mRcILUU0Eyt0P2sJVh7I/afA+EuWRs
aNlHvQKkdxioP1kiqLbw3RHG+40vvdPfxJHUl+abVkmErj+a9swrFAEzIDXRnGLvNwU4RYUlED1J
SBa8ETCeygPcyZ8cV4sMr3Bd8eDGHBvYWMWA69VFLxhXz0dZwEhP4urKomnvCakxkSupgxMkqPcn
CcC2x0f8cHD2TW5RFlXpY4z9aeFASWVyZOtqnGULgWVj5r65nd+igfcbTaJjh/7LbX2ANrueyQmH
XYsKNqA7oHQcVwgI97BPvRBJB2oktwPGQqYD8KkggDDaIfa3ZuoC5jcJVBdS/2PZyXX4R7/iNdWu
oHF9e6ryhGsKSmh3OJk9L0iVNuXR0Q9fsZj4McDZB67XwELPwut4ZXb4xobx0BZFC9gq5qI9D/3s
Zar8YYSExepn2T8FqHtskiJUxvTFQ7yCU8dCPDwSwqeAAqpLSIqsjPx1XGI1fDX/GiwzmSwY623A
zsNpS8YgpFXb6pwA2BwrUu16lJkOw+/h+fjJysS+Ja6dyJ0gCChhK2y1/igrhPzIQbMH40Y5zwDo
GcgmZJwpIXpcdqg6xkxAj1cGOG2HQJNbb3PqUL46/hB/msEYuxH961YA70l3p0oaZghssO/sQfW6
FTQwssKcDpTvl0mM8pcysQo6uE8KoJHqPydo/MceRY5vVoe+k6e7SrD3F7J6iVC0ZaNAs4zG+WGV
aMR9IzH0XJyasPgRuk+89YtlalZ016hvuDijkWasB+LclTn0U5f6kwDGEBKy8XtWA0pqhom/78yt
S1oAsRnLyhGaFWWSz/u9vSvqJDgznuE31ZBs/vxnkSHyq/CJxqh4eibdB9/SR7VHGBBgjoRM+HyQ
bJxWyIhUXkZzf7HEC6jbSnRtro2W7DYDOs/aEaPYoo0lp6BDHe8S6ku0UZiSN95EiNw9cc0ycpsU
DFJr1iTWD9Ugi1gu2bMHhrKUB9iGV4Hy2sECIysoTfS43xZh3Iua+XLQPVcXumHnmoJPQuM/hrYn
z7nW8b6Wgz8tNMs7681XcVWVa3N451NA8wXMi6qCVn1E27TAgwaJrXG0n6zHfmW8pulWKbLB4HVk
GVBZuFERGc7NvOfIeWFvmcVlN7nRiqE+svAiqFZWOOodKN6klIyaXRkjV+yf6HBxetYfwtB4p+NF
vsqLN15DK1WhPagl1AmO9BIe4lcCLl+sW9ScubvzadrR1Cd7BEL+F5lwA4rImpreWN15bE8sSOq1
i/E1VCaKGr6Mpe1haWWNUL/JgCzKSgl3nVlEpyMfK2uMyMDNyuZlCSC3KD93sLQIODkk9UUHofDg
JgyHkLBJ16OCeh79B4h0EFbmw2CW0WwMjVH75LTPHLZtzKirp1Kue/9bhw2cWPs2pwyMk04jJzvW
n9SJ/oIgk+wj8S+KPsBDj6g7rPAQX7eibkRNIlHBflzKky1MQkKZYgi8SwgE2PRYGyk1vva8PcuL
kudJMXAi/JmXGJypIS+GbIrmfXqW8sd046uVZP2qWf/OsCPhuW/yEwjpSdvSnSgYSrl28b6oxMwF
2xFmsJAvS71NNn0pP1UwMDiXE3iKqDviekctmQbLUd7r11d6/OEK3RknPmYYlgLE4naCMMbk23lK
Z3L2di1itBhDGrNzIai3grJUCDPTPFT34prazCk2bKh68/RQSc4FTKNXoGFASNsLocR4+IOYOjiO
nFODKz4DRCvtOSaAvM+1o8M6hHSMtJ34DG0doEUgLwJFPeqiGy7mcXPPFbbAmTEigOLt6q/X5UXu
q1Ep8UwsMETd239DaMQHF2JrD2AGCZs000DwGpPCq3DidhPsy4HQb2IfIW0+3o4dHHn/Nz8QFJO+
FPhdBg9vIGITBzdvMljXjx/daYzFdNbegPKs37SYbKgeZu8SIWP7rybxHmKtnP/hGkdXhmw7+hwV
fpRwzlHdHSyN+qN7XAj9PEkW4nm0+g2jb9qbrXjrU3aNSq/DfWPkYAbnliq1xZVrjv+IrmaciT1e
AAdoOIjojCiCKqMBxZyitSmHhQlaPYzkuw7mdm/vC9qCLVew+Y12N1ije3tBSHpp5Ee1ktF7McDc
IAb6I1x2kxBEgyR1hipQt7/5cGoJfgPGDZUT+9jtQmpLm4u7pC81YGyg3Wamo3DgNBKTNkkvRTaK
XKiETLkDyEAcDFWNYVVOP1TaGWYtuP/pVavDPLFrcrrfw0p58h3ZZbZzAxnk7eGs4dolKSVHdLXq
QONcBry/moMS/vganyzVGfHizZ9BUo5LzgcpN3aA0jcyVQZyYGZUCyddAd4RRfAKurG6ZIphXNEA
D+dfLdsxg5FjILXxD4PrgX8yzeYMwXtpqkYgr3TCgi2RsodkzeyGBt1IUodpiSTUWuRCYafgK8+J
WfTvekSj6W9ywjScULp580TAkO22xLxpqltFwhp2ehvAJGA0L/zwyq4KCqwkY36NWg3ox1yGOCYN
0URELJ5koTfCrdL3/9N0EIi0AvXFwXxxDAvz4oPQIh+01N+iwx4p0RFLJpNFvOXUEf1lOFtt/O99
P0v05WsKoD/gAxuXQcVGJHtZa691WkKKU2gbf8IbyRgDI5YA7KbBr5Ikkd7JEp1Aorf4Wr1uBHrs
Hh+So+m+3X3iTy5/tzH3f1NvbJ3GOZoFSDxdJ/Opthg6Qx+3vfOAv7KoKrgRXHeZNmstTfPYyiTM
vS7ff0HlSLaRXSDpGd7mb1+nE+ECP83kgrQsOYBKNwf0QQM+9Ylj6DjBc6jjEu/5U3VppbvQVCkM
WnMrozJC5NIFU5cOcofNxnAtszt2lQeA9I/F0O7QJ3V6rdEWjakA587dhTEBujYeJqYn2/0i0Bn6
oOV1SUxC0KN9Oujw4lBQwdOvqUstYMC1bIMIJrSSEsR43fpQ59RpbPxMNuHiqUHK23+g0tMZYOmc
CqDor5+Fv+AscS/ST1AU4b/z2hJPQ6jpc/FxPEJaXINpo4AAA3elNr34x9TeQPLVRdAv/ZvTBPJG
9AAeCgqZa1uG/5qiNFN9wzm4gZGqWoKb88vHOxcB87ThnwU/OYtYI1fRQd+v923E7Iuft2VjUFPW
49iiEZoYrdeAuBjKP0Qo2fLIh7BvihkhQq/gir5Pl6P6ALlPOipmqydxxQ72FejseB5jZrJqBQOE
F09ecUF1QngmGinOTdrTtLSCKajS7QSWoeRPELfsOtM9tTRx2WDSJd+mzsKxM7pemKdA6u4EZIU1
9dIa/cAJU96cb7+LE9CIPCLi6Yy07PuYIEn0arKUZ0aNUVdHfDjn3MNPoUQlkKkypzSOI7cV7d4w
7i5LyKkMuUQdpac84ujgV+wtnF/1WiooMW70vtfKcR+m1KgO6fOrxVfTpsHLTAgqeItGF6N5yIOW
RNuFt+fBnnn12ZfEHOXAf+kR0a6CKuDKKvkxoW5ciMCvf4RsVYhkSmRsOTvP6XApXowfBYtG/HBN
aB1pD9k/NVHKeYebWnkcWF+TBDUGd7QOSi+nl2Ptbc0EYTl0PxvoQI+qJqiwJ6O0QgB2G9brEBaO
+6eSJ/e+ILdGrvbfQH/uHORQdUVCFmY8b6S1yLO5aDhALAEmLUg8chCmklhoH0rCIFluvhF4xU9z
SRzPYAtfrjNij6FcQ9BvVnyzH1ztd37L6bdLoruB2dcSERcTrcK/A0rLJpnS4wn+RFABQ2VzKye3
9OZMnCX5aUdQ4H3n7txAiw08RFx5zPy6eA7qANYcDfsXHxI+MGAL/go7RACO+/GQTZXjDm7rDfu8
hvU8itPseXg8W7w/6knlYUyBfJr07XYKVUF71N9m9X4mmqpo2WXN+zNEzDbiV7BcZVc+2ZYYcbDo
FuGTeJiiB2qJUzHcGobiPGZtWH7+qr6/4lx9VuaAkvkgJdp3f5MKUWA6n9YWcQGU0ILxttu80srD
uPtIQ2+qdT21jSGSTOSOyhV1uc9CsO0oVQHynyvRt2nx8dO1//yyxUb4OohP0yr65pi1UzVl1MwV
fgbA7iq66SaWgk1PgCCLnGAVxnvXM2c3mg+PJXCfWrx+ZdcXD0uX0YYL0Bi7kb7t4s75W22oJVHU
brbNSuA4jdQoFR6F0Dyy+V+cuptG5W5B46vLGtMy07F+pUDTKV9l/NS9Q3SpwI8OdI9NLfjoGjSU
zZZLhKt2M2OdmqxgQz0buCVf01+LSSBJ5QQDkRHnIjV6qRAIArN6ccc63ouk9JFIkkexn2JxvWD+
n5n07fY6wm5wJwf+VLqxAQofJ6pti3hbW2jiF4+AgUQdrZDrkFaR5wM3WzWbFjMAGXEonPWARf2W
izQcX+TKyL+SYvxm+Upkxreb02eA6p2QMxTlECdeqyVS8U0GLkzKm1sejlyDDk3eZR7ObPYCfdXw
o+aLMMhjjOWKZHOUylCPAe/IjkbMpenn/cL+5oqgzsH3rTarc33lHwrGNUHPdcXUZ79TLw3lS25w
MMORifNGSuYQ/1g1r71ENsUdONFZLUfu0zh2BRI2spUi3EYdSHgrDSAGMeT+qEBB3Zuk2FBzfPFa
ThNJHkol9kpKQVpWyOI4jqWxlJb3dbpiRyZV0HVgCzpQG36Y/7m3ruXIgDsYRTXw1M4VqrZDynTe
oCbe+FgEL7dauQHb6R12OX+/x/nXkaNt+b8uIQvbHvqwcVhzXnIqFOUcANZL7knr2qBAImikKf5n
DPcDPvJ8Yw6N0ZcPpJf41kzMC1x0LomOQzsNzB0tanO2YBreVPfGWDztMA64rHXoiAlRRH6b5EbT
sfvPJh3e0Emh713IWKeM041zT85k87ePVAZpkrlGCLxB/bYN8f4eFHz5sive8OSqaJ+dW4n0Zfea
sayIWCJ5GcHiRd/4kP5ouzaIkdZmbrRTmLt6lK1rJjosAM22Guyexi6Tju04OMlplgknK6WC0mOb
KY1l81NO42AsT10eH2AzfYNPTNh97ee+aWk2vUNkdCebbIpLKZ5qDmd+7esp8rrDRzDfEJBlCxqH
Q11/GkkPae/KMF26EhUlwyh4USBBn8zWMBvnWUfsx4Znq4TcZPapVjoF8aZATOUd8l1ncmXyZTWZ
AjhlxpNlxv1VM17UCsveDxl6hNa3RcjBJ/0uh5S7lptx6F4LWdhoxk54TY0yNQjkkfwVcxPDlmNh
0O73JI/QDRycdwPPVe3LaSJczEX9OPJLFc2LDIwihjp/3Mf9GEQLTYIxule4SFcCgpSvv6E0Qlmi
BTLsZHAlVcMLsU6xLAAewVsjPeUxJrwadqQE1MCL9dK9hI42AR5ZFixB9Onk9Z6bS4VqtCfNW3d+
rpGC2GG7Uw8ims0CiCXHQIXtwnPtI5Bsktx0Bp6cjdVyB4Cff8O2fKpr2uB6YsbZow8xv69x4dIZ
SoaK4lB+4xtLoe5PsjL/Th//wY7m515cKqZG1VLAhKvZRXELDLV/T1gaYU9Vy6hMZSwbJFXu7Ygs
rJQhLFLtyfBWwoYHXbP6dPj2mg4aFJAiVN5yUR7BW2mvKaY5T4oT/V3cXlsadvH47UQv82QSdui9
N7ATkg0/Q71Q98fUzeIpYCUFn3B/ARbYz7pLePfa19mUY8YlJDHhJ5F8H8RR6apM14npiH897fTf
Rm9F6RpzDvTlYD+F/iToO4TLKPKPj3U0/j4hhPuzNDx8LPUk3IhQLbfPs5DFTSMbs89J8itzLHpl
/WVUf9u6BVkB8SajIpd2rSUtv1yqnMwLll9C+h2giVUI6//MVyZBOFR1hRhJCrOiZk5+gN6w1TNw
qQRf+g+y600kJSgH1k2m2zShXfTXdTDH1tBFngJSZqsMGVo+DxolWQ2uKGozqKy7uv7UxLXpUZQE
ODy1ypjcneIv2tWQEQY6dTcP6tTZgSzrnEaPQcrJSotlmkQbTfxA/oaedkS4ScvWzky689tuLijL
vSS8kIndJtEmaDexPHjWJEtl03ZrMi3fxhuROfULQ2lbOGGaQ76NIqabMSzHHpPkBdLgEEM3ElGc
KJIBwII61Ka0F4W+tqKVwLwpFUyRd12tmNZENqO18Wz89YQHX0qNB+N7fZBFp5g3ke/qlBKzA+nz
+lmSJUnvLtBI/OoEFrT0ctIBX+cw5GScOxZwapb+yPeu2AZaoijYS74q9Bp6lYRNUlAfPN//qzzE
UDUgofUKcHTbTo7bx9khRvOenuHgSMaJVLL8G7iNedeRKdcPUBUUgNBaYfKJNR8RowKOCRd34svM
I7+RANWB4qqDxOLeQsP8g+Wk3Getsq3n2LpnHO0+m5AwtwghPD4Pr0yUm+x6rjaJvpAG081sI9eA
WlQdFysSpPlU7ZSHrV2Ryf+E2QHVS2OH7JXia602iW3TDHxyU4iRUSSUj62EzrCfM3RO6UbLpzCv
F8cvTUdbjlBIj6Z4dJ/Ol6NAxcGl6RhWfsjwM3zDTOg0tzhz2LGllWIrUQdDlOkrX8icCVE+ZkKl
gHjBSpCAGI9pimSYHteMYP6sLyb8YrKLh3ixSHAz2CVIiUwA0riTCz4gsSR7eKxNPLZo7kJe3ipD
EkJuJT9cwe+aNAbEH45hVr7fFheolYnDpLhApH6wdapPfkKIEZmeiUM0Iwqbjq7oujeze9CcpewQ
JhICV6bYP2i1hKMr2hy+zVBI88VsVLSvChj1sboc9gclLp1cT43tMvCPX3ITZYjm58/mkL9ee3Du
3Qc2W04W1fV8HqmRnXcsXy4oSNwPi9nnwmEaJPJcPw1VRKh6V1zd6C5qcI2z8rrP7YYBlMG0pPsb
b7hxTSdnswbyJtE130Q87K5zNkjTHdgfSMFzYjoWitNMo6cDU57xMOH1XlBB2qn7fKFYBVCT9e7w
5vAquZBLFSOM5MsJ4YIB90sxlxQe6IjFUwfDkIRN1L2+z5+btB23WXHlrjP4mVVpkZCy5z8mi5o1
/nMhM8I1mrmCkeB0NmXWHZN9Uy5ThB80MsdJ176m6dPfVAWK852HA+bRDGTkgB8kY3tAMNZlLl9V
begGP3RQnSRavA48OeHxBJBCOIV0q1jzNiloTQNe7PL4YX6WW3UJUHILr4ZDD70hMmwesL8jfOZc
2Olw/YzA/4qBeH+TOXapoGEfsc/QBfHRpXcCAVhN+1xHT4+H+i8/BqXv4XSgqY0g3qM4l0o6UKrF
quAtnJQMcGDAHVqj9q5MFWRwduu+ENgSr+ocCpMYAd4DORiScXpwjIMQSuLbwNLrNbKuJAzfrVA5
93Ao5/YRrPfhLbWdJTrCBneSCkazqpGv6l3bld2g/GxoQ4Wg3enLHqvL1qXr4kB/gwuywNtH+jGV
ypFwyKG4OyBV/PIsXx0cBJig/NpbWnFbPG4z1ehIRwRqSqf+wd9m5Zz84O4snFfZ9S0/xBM+JLax
moAdRgH6AN8jaaXZcJ3vCasIcEoX8l4wddgI0kVBs3asI7OhFIRPyZOG/i85MglH5h7N/plFjphb
8L6EyiP+rtVkWIK8DRq8DTltGF1H5jSpHmDidTs7smVj2n5D2z6CyWJxSv1qT024HP3Da9zXkYcz
xvytvlvLWkCGPrsjYZ0k+0vN6f9AxfwwjDaiGh2bZCZeX6SDRNge2pCPXHSJst+0tfs4rDgY8KKN
6N+/3Pm5q4qNxJErgrYyqOBb7oc1zJYe3hxpGwkFIS4+7mJAeoaMIsYifu7enP9+ajkoFLlGfCBB
pae149mJfbU6/+dECY2IWG2WkXKXLQoBsvOAjHfiUHIr4WDozeBuj5GGcbb8JOKPgd3GFIdKIC78
+NlmvmpeIrCRnFhz9DA+PYfgm/k65wzRpJp2rP8kVoRlgs7Pki1BiXhEDE8gU2cvONbrRgKxT8aD
t2UIKlF9IY68Xjp00am+ZsxOtfr5xHgYUHTN7uzufj/DR0V0Qd1dv2/sOh/SmIjsHd7wWctG3/Xb
cLZP19RyFMRXpO4CYwlDK6RPpf13jBxdh8HP0lCj7uXAS28UxOPvjD+FBUxkUicXMnfWDVtXMqBd
f1wijLNCgQHtNA18zd9uiejZGSZQhBKRZUv++Zc2Qi0L5o/6S08vA2HeYCN8WUbJt6BBNl+/MYWO
8VE7TAtUuHLDhb1RYaJyuV/FL2fYBGc0p6adlwqr5qwBfCwIPsgs+mHCYeOdXrZ3hDKhXxtnjXyV
dLk+HvSRWw7hnjnkGmiMhs7TWyOYT9V/YjV2oLNqSTv3OiDVkXq7OlmAa4pNNvEt1WjCOKRyAxjy
OIAc+o61gs5b/Kz7xFtCaVLpJINZ+qQA1r+76mBDfY2xCvekT6kFL3j1YXGGFQzHpmy31eUlNfqx
ovtleeBhFSAMefaOTzBR4Y01D+tfabb/QIrb04meDX4cGWlPp7ev0hwKLT52zt6yiGnYhEy4KRR4
uqcuG90jEh3pklpPJyGm5BWSXuBlGEjSnMfZzoQMommo6J7XLlkbMN8w0Dv3GanRNUg9SL6ZCkD1
d4jbr6J93GOiKQPmgc6sjTrGfhZNF69zncCcGvtn8eJT14K3CPZHOe6y+XecUHkR8gkCZiyrs1cp
mocxHk8LMnFfsInKlealjyQKmsyOIMQQgWiJe8ujTn52T8oZpA4d40Ut8m+5MnJvt8oHC3p+xyS4
iCz0XGtni+JvRJVFFJiL6Vd2bg0g6genb3OWIeByStEd2GONAGhB98Cq6x4gejShIU6Ub1Jc8S8n
QMr5iYtAmST+4jzaTHoqCrULySnwvPP/AwTX076BSMvC4vWjUxc/o4OoWdmCWvDKSVfPDe0wO3pj
/oH0Kni//JD27/KVomti0ikWdpQieNs82ePEuV8LcCaDQqZJhE3hPH9Ca9xVOdS1mrTXrwHnkTEj
gsHZifAqpgGU91u0PHE1pwBR0bHRiENFTodXt7FaqoPFRuPzNsyku9WfRQ+RiwSdnSrPMATD4xLR
GiiyNzAp2bVTfooOWgKc+RMmSLl61rZ9ZjBCoOQS/ujQo7p2gijdb+TAm6GBg0coC8int9XQo+Zi
r7p5GT3lDi8raGp14MZYXu/fR98VUFHfUd7dcVbafSpLENasgJjxmMYvCN1HX29tzzkzefWeg/Pl
Fmk/TQYkFnHPxb1yIIAUxmmzOC39RsS+xEOEgD7RcyGX3ucy/QS+cz7fcNtoa2ud8Nq+Fl5whiIm
+Vx1uMlipI2xQnkhC69rwZIbHzSAgpXrvU3ONchG2/pONw+GOxpA2M2HHVs+grE59s2eooIqdoBF
e5zhOGeGwQi4v7vMg6n/EFh8hRrSLqk9TcUrctFuJhFvbfWGQEjYyd12wKQTnhi2dyD/w9hCuTA/
gdjov3wfc/WbVwhWfntqUktp5ystzWYayDSi0/EBR6hrcyiwFKrx/hjh1CEuXuYIU9gVTNxDe8O+
KM8Dki9qFKOvRZhLbi8nOwNBGXFOCt+jAXBMqRwmJVQgYyB8OjeHJ5uoezC6WONt9e3qH1VsHim0
XPoohAcP3ZPXQjHIMioHy/uyNIC8VaaIzEbDadPgjrVergdSybHvSAQ5EPr0B5K4wgbefI4k7DjC
yjAYGA4yKuXgwRT6ruZexlKhB8SsMd3kR3Two7WoS2nkqs+xRzmxf3csrVlXVL+/djqwIoPTptNK
o8kgV1xyuZcGPoDkENVR/OUiLEnVcX1lrLK7BI4lEqbAFSxIklxBisegW+pxknX0riU2PCKpHnkE
NfgcaxcQFzfsGgArAV8BhHeha67tWvqGNcr1vByfH1MI9ql4BPwDLUpMmsN9Ymx//HXq7Q3equ1q
u8Of9Q27Xkq3nn3/A04fToIwEcyGmiLZzsZaGH/RpJUWPbkf3gcCPGqHZ4vgnT4HZyL38YoKr6Ew
Uuvy3aWmhy6fkcEKeAPygGP3ysjDx9isnSFyEfJExuq/0vjv9CveXQew5QfqSgA8CeyEXvWdKVWW
nyMX/GNYekA7nWSy/+gYPOlksNeubvAaJHf6DAuqHVfTYNpef+bahnXhancgQkHFoRlftbUHxW1e
nA9LzdH1+Q1LAFh9r+rrz+5iTXXDlflhlaN2EtcBoxToQl2yIyE/RFVqut8iBc6eVmLYTOQRz/el
FqQfoOrVXP+vYDEh02HSY54VeY0gj8q+45XoOs5JA1DI8YlBxO1RXw2cDZK/QBaTzNLFllZmwz/Y
DPfANc5ut3AyMy/focVF+BRTqgZNomg2eOc3amxglm540xFb4M5BLXr+uxszWlIkEhFfewDiA9t4
AA/+R1uu+OpxrDvWXXae8o7LNSbvV/w0pjiC8rG324cLcKCMvk+ZDPA3W8F2/ksU8L6qxVtf/Q6v
Cjsp4WAiohb9wW3azlmYeJSaSlNMB3jFJ2RR9IL7ggzzq5IkcGAFsOerHq8ScL09/sKoXSlG+iM/
956cxfUnjj5c2ean/eHwjiyItXvL5pS4FlU2sMpJR6fq9ajM2l2b5Zzzyfm0Rn0bQojgNm26HeLp
7qLv8e/jQWt9WMcFeCNnK2jEJa9GbqtsK5akheiqc3DJ5Qrl5IDfx5EMPxFMTaM5BVAnZLmABLiL
suKSbTCE8CS53OdMXxgg9O7ABxWUgBwsji97X+75TykcvS+//QzJ94oM6z7l1XNbN0sCYoRamWC1
RGMElCBV3yEPWAscfRw8KDyszAJdgw1I+8+JtHlb3E4MHJ/0S9AN9W3bk6msEtRT93gRrknt/WzA
fA8qTDAfoRGCCkvPUgvYWmHRRf/6mqx6B8ZPFwSp2iiG9nyZimMsp0ksDVfavpbYpNs2ijxJpUDt
K5FtJiKdDQX5tzFvTtEs/K/nqB3McCROCIJjMu5zBQTGIb1LtDJljmJ1DbPnrmszEfauucS+Ozkv
SXw70mNIrP6XweaNSyJIzXFscEgb8ZL+v1dF8dBUiXFCzGG4Ysq2Ng6macf7CGvT0VLrBJ9gjl6O
tXzAx/HTKTy/asZ0OP/rNL5Dzif7lNZor14v0Pud032vw6YqlWzbQlG4l/WV1tPZyomHHkBJEzOV
sRFxhWGRARZ3bdvUX5LzVWyoFnZvhVFXhusjuL1kDC16gi9+xVD6thAsYSTbIJ4NYu9HO1A7ekI6
DV64j4Xms9y5IkDFu903NbFQqXIHllgRDHtpiLRFgId8v4qWA4QhM92p8rKqnehfya/S6DsbJotQ
gTsSK3snnMw5ZPgwDegctQKvuoGba0EVJp7nhjmhKApwyQcINigaJDtuc5jnabKSyLHMQkZG+0DY
TamgjoaALCRgP2LWzX3Nttkk+kXmFl2N/d7Owp2X4eS5SJMf6sDK7I2PshgeQiXYnWnjGKaAkRqP
6gRqiJvkBxR/iL64swOT5bRUEfkaxPNqIZyh/JhDi2tq6Q2azeBCQ/eOlOkZ8xeFVAnGL3I59ygK
urbfpF9ANXs9J1/2O9xSc3gFi+omVBGs0ceoE8PKsEujPeDSxI3kiYCsiuFCv++d0oYdg9EjIx/4
oNVuJFcpEnmAP6tF0PiJpD1pW96zaVydLLsgGELnm3nGQH30t+bl9WpheuicWkwMQkdt4PvQmK9O
CDN3hDTLe6LTG7bPSg6a3VklQMVazRl8WDd6eHaW+A9liyiVcSwCl9u4pnuSrJvCrimOfzrM6/Rw
HFPMcHWugMRu7cHpnCK9+4Ng6qjoUQx7ff+o+UzWZFjB0K5H6m3H+8vd0oy4sDK+j3oSnXRC1Gmm
oK5dzYfjQfOM/61Hk1uZZ/FzRN/n4YoOlr8XSCzr3U5aHTxj/qQi5PUnz7ghaKfe5FfggGixkjqR
gxCX/Ux/5qVqUk+OcaVag/VrsLKrgfE0w2OUivi1NdSwW2sMFcBArCxUmWDrFLb45YOhbRPHKVtF
NbQq85xzo6+PQxkEMRzTdm8Uil93MsnrtOqpfUoxq0nr5/nJJq6P7lMu8BVpZB6KJoT6KamOiqQ/
RP14QKVZTfhLB0vGnGb9qSXCNFYGINQxkC7UikbJ6vChGxRI7lbJkbUL2Ax5bUOU571AzNMARBhN
9DAskN8uHUDd45vDnuSxvTKQVSk5gxZHYO5/4yVfXmq6fkj6L1a/net1F5NY673DCF/qy4HYxDPv
XsWdwzzccc8PQsLWbQVrI7agi6AndpY2YXpJ5Ic7xWNBbbUlJaIXIQUzhaZ1rZZ843t9aHgit/u5
Ix69I+b1bxW/dqPD27Uc78zSDxN5n4LwjsgKQTuqRPbOQ0ptrM7RwhWDAhqz2abTCDgPQmy1BB/Q
QF1Z9WSxJ/7avBXbe02s8Txd1W5/19iaO1Qbu+yJklaOW4Zf4HyFl7yE2YqEV9AtlMtSYFfeViy7
wssfVXTjnc9W7ssNKu1cvkM46uocvWPbZ7c0381Amy89/HTv1JfNxcDzrFze65tdUgoqB1HQFg7T
jN3QsYAAtEMvQX+q9c84abHW3rOFIZtpTgL3n0nVVjEN5u4h8MIPUEYW7GExutaVSWA8EUIx5AKe
Hzfxcvqt+MKS+5wkR5662VqcLiy5/GjjXKBqnS8HS+tEqi4UmgLlWLdqllNIFA1hmTZp+el2BNA4
KddR6yCFyCnE+GhUM4MZJD7Ozm32LAl1m9qc3w1/iUkKu3tSPMphpwfZFB5m4yi5gEpwcb4tSwRO
7Ttpd5KmbwMDUNYWru2DQK3Y9T9esjbEqkXDqJWxj12RGehk1M2Hkq3IjZl8Meq74Hca3Q7485l+
Hsdxcqo6lcklS6jPhZR318GWBXBBCcZiNZyy6FaQmXIzsbxiC8Y01u1bUurG18VySR4TZ4CVI+XX
OB9+L/MiVp3SAA327i1IYSjRPYbZhR5oIrqOM335RAH3Ond3Tb6mu8p4e7Z6i5VrYPNgW3bfO7K4
Fbj5v49Ko0IdVl5cYl3bbt/nWSI9z6rNcqdHlOY5XHJHczLIhh1Pa6vhZpKG4EsZ7DfkXL83Pc3P
cbFksJ3IFn3xuSTthhw9CB0ztYDkoBDpqte4KWTY3uMfh8sAOok8NXa1QhfcteNDMoJuwX1nZGba
gVNZYvbF1Q2jmAPdrXK8OuzOJHd1B/cufocW8yRGIq9qA8MyScNg1THN4Z44aUYorOHo9B9gyEmn
jtl8D1CA83ARhhSIWozSm48WfwCf1Q1BzAVzCGy8H6qOlud9VMT2aJnfT8vF8GeXxRO5zWxJfXUp
nRQB73yCWXoC3u0uMLOi4Psk3JTe+1tH1CQ5Pfzbz3IXY5seYjqGMapg/jNXTgXhvteiuKcllU/t
J0PVQ4fD2Us7Y9SRPmEfK6eUV1Pt19JJGVdCHKuB5dCkJGTrgAxoEdYahzc7iog+cnUoFvGKmHx/
aGbr32cHGZyA63xp4IfkaiaTDHom5tkIzjwQKx67lfGn0mXD6DRxlJAmj6dEUxa4lgW0BKLQvNn8
V76o1C3jf8NrYN6l3T1l0CpQf/brLyjXsUsNauVt90Z+CX7S4HqAQwxJkbBqGfQ6JaczgwEcyzFA
2GUjUgw8MiNzp4zHSMwuVx09PKf3EEgl497nFLzWW2mdUpqCASIaC0xh3xZ9WgWR1IoB3JAVxRnO
CQMBb7upJy56xME497ruIKtaVqZXmr1kwn11KafbixLLYA0dQYAMm6xGCeqdBxi26VWT6BUUzAij
mGvb26/XCPjXnYsTy+WgJ0FrqqERKoSFtA00U91bKwb/cNik+CQ+G4dCJFWgr/JVQbStw9/cs/za
ofRnksuUat/ewFJVPvaiaxfoKFWURCYWIiaeZC76TeHMkxRAtFLwtA69KiNXL+NFMatGQ6wvyrVM
h4BAFU8PKnQ1Yl6gYFTCs8G4fSu6gaPYhdG4aNtddmPAwT80KuZ9kmvs/uXa1scwt7YQMVRFyYfb
hbWm844Ln3tlNgV/PP5eLxsijhr4aBbdGaeDMPH+ICRLbrjqbWpIdime6j2O6fIg8M4kZiM7tO8c
NW9VGHB1IWbyco3McJFuIjJPpfz7NdhubUfZLKeK0y4c3cSnY9FIwobAd0U1HxUeYYDW0IEKfYUB
B1YfrE7DlGFwWqI1SvxneWZC3sTBB0nGVJHSNIp9hCZS8x6q67vSZWKcwLOjpSY1XnjFPVNGpBB/
wXGYNJ0Hj4K2xKey6Jx74xn0RdPK4VgLGfl4JZ5eDFcCoxwBmHpKkpAJXOtB7UbhHpmMGbOXzcqd
GDpOOwj9IFxFhkaSFZVz++4WDUCJNJj2a6vYjiSWkauxagF7+VggYwaNO8aoYo5uyd9sC/Bvw3gf
tDqbyW5I6D8uqLgnqVaxO4s5iRs2hDFWt3LlLNK8RuEE+dozwAgl/gthzPNjjeA3qkyaCh2FN9Lq
gxYEFAco5iV549wX+af1whTbUahg+doNYH/Pw5BEvVf07tUAspNhGtBJ50jrPbfL1oEMFWMOetC3
lLqT/VXjWZCeK+Ko5z1KCEMgK8m0G4qCTgDd6touuYbCwnR9Zz2q04vx/HX8bXO8W9540qdIr4ZN
b8V9yvGUZXhuQj+pvKWOkc/o7+8nSQUiMpcE0mVhivkfTVWFY/C2PHoxt2D0SLvTTjcYwDBcPHqC
Q79Tq+w/Z9EnytQpUf38MxZFULd2F3xWBVYeCBdaQ5AkbhEPNzKgZ5Da8wveB8Y3vztitoaZpidn
GQ7dUEp1MCck5uyYTqtSY9cXeRmhg/3gVF8hwSfKbvDJn8hDD2W4aOqtvqgRpnZxtqgJ/MZaGUcX
uB/nl7YkWH2tkEOh/m497xOjqaFq0Z3HnuVWmpTwuV249b316cZni5cwBYikGYfk9GWwY9nZsjBN
PRBDcJgY6irC9K0qA2Q/Wi08HrMgiZrSpeluC9NcXAZZ/zss/IuqocYOAWQfa0GX6TpNhpibKpzd
BHK1R1SmjoQ3PO/AskgFLhNMFurmUbizfxe5iptxI/pLWe2OY4QoYQMxgilfHT+kvpVGM6iY7pjT
YqVBmYo312vyE730jO/ZdjSdCZWImTCD0u59NuxqAdZdnjgO3wRkxZGYylmmXo3Mph30Mqf2N8WT
UHTKDeExLOu7cl20Ovb/KNaHTH4hPA4esXvu4fka8z/g4dlsC+NPm7ppLru1KyBjGBwYSv3R39Dn
x6zQI9je+gptu9X81PpHGBgmAz/lE3enrynS78ZlhNzFOXGvjOkzpWltSSp3UEEG/nC67IlgvvJy
lIioQXLT8Puah8H5ci5kZt60luKj+RvcrAmqh54LBhe9KYpPP2kszOq/vEz+RUsEUCxmGYFo2VW6
zjoRbhph+zbIP+Szu1dtaLY5UI0UVCDfSniXpXnSUns2j5DQXL5KtcFFy1lqPQy+xGVAib8LNGOu
rE/LDTcfkLCTWcS+GszQrY/gr7D3ndKXSnMfbWGrmef+wmEe+GIs3CTEpMejPywpxYdZZWFTLmz0
DPNXg4e71lkYK3Zzo8kkanI48S43qVFhXAjmVvm4eWRKkujaFCG/xbMsBpJFmhnu/Ud0/CdjebnZ
XDMqkvAr9+vMKm3MVT3JBVtGAN445M+mILM18BN+IagACLvoAmisNyEUueRTl/QWkbw3+CzNYNj6
nmCAhLtfMZyvroBJww3I2f4X6KSRd2cMT4OkprEOqNEjUjM9ntAK6E48XTmq6A3eAj1GOoPryv4n
Qsb/NuXITRYcBhEIHkDsCbSO8nQmPVkr8wI8hkPWOEk45RaJ8VH6RQtcJ+OGWepIpsta1YBokDa3
uhztjBpWrUH1z2DqFiVKXffDMN28xSO6lSp5sEBWad82jaOjqUsw8ySIHQrAnWJa+BSRR9LUE8vA
VmVGHrnrznjOp066UOQZP1RNjcQTH31+Bv1pCfVi+E7PaRiemqltmX1hFDD1LGFApR9ppbiElVWs
6XvQqKn6F/S4qHITIxOLZRUTLl3KHdcc65c2iaCnKgW59wLujQitmkRsvrd+YgXQlO0SPmoegC3u
9vhTvbIJPsxVsP+Cu8NPFJRiS4DaVhllOG4NdDUvOiYcOt1ABlVNXBc46wyRuqtcZrTut7Kt/iH2
VThz8YZHOjAUG0qpklnpsW2En+p4Eua1E7xTJvtcQZotQNFiEZZajoV+hzw1M67/UHxgtbzgSTN6
D5IMME/1fvt/RMggoOgSK+Bl+A7zjWIMXNqYctEYV0pR6tKSTGGCOU+VnvorPvmhL3/AAal5h5sz
1srjbjaNhctivP6q42JGwYvwkMUQwKKsSW93mrsU+tfnUCA2GknJfnSLwluyJBXrALev8Hmos7rE
GR6MHhlHNvO+ZClOO1cOV1tYTIX38DyL0M8wY/ICB0ok/TTH3IjzSV4+Wqxz9cHim8OjISaT8FZ5
1pMNqpSrHbXM2M238ajo8N78fYIphxVHq2kVSCtwVEwhU0jHN6a1Bao+FswbtVjjm3+w2YK1xEtQ
ExM2o3oTKPOlbuPjFhIbpcSlDcH6pdZqyQ2mM7aL8nM8iPpCskwL2EZV88dlQCtT6MNi3tmsZKtb
EiDaBLPlDfSzToYBXNXGi823JUeNOlYf25TbpIq/m31lATYSfc2sAgW/lCWaybOm4kkqw8SMovfd
96fKPPdGUDJx84VwXw1VshT1CH2nli5BOdBnV9Injw+zQPxwUyCppml3MiKTLQjc/d6KbPeQysbW
Aq0QACQN6fQ1GUO+p/TJJ1hs+qrjea8U01EeTlgGDLeXd49X71cNeRSdN24giv9Z1k0nHVqY0LSm
DXCbyanjyNRlaKxYIguDsKpK6NIoKhdu8Q5QAwCIVT858J/M0lJqsHkIFJgaVJPM4LCabLJub+/2
nVXFdLH6GPGu4bFh8m0rhnl5txFwUrlL9Ieheqf9kfxKxJyydgkINVMq04jdrv2cKyMYzeelpEu6
lRkVfTCq/cxDmPEQMpfmMIg0A20iR6/64pH3l8Rrfy2UGa3rQkQU2wVmzdsr16S5CH8grzeMR9WY
sY7N8LQSgchab3mXeN+zHuXHLzBzV0FXJlX96zQKygY9KdWY+7EBUKWNumjVPF90uytbK+7SJmfq
hXLDKpP7Saaiot807/l5X6DGSJ2AflUkSKMqefS9BTO1jG4pG8tnhfJ1YWLkdWk1eqz5t/ofRvEC
MF9Cw2Kvm1Y3Eavg9M0/TEfIAxhh0mozMGtcH9q/Htdgqeyfp/VZdhxqrBV03sMscZ1T3sY8qNut
dBlHV0KwVtIJVS/z/tmy4telzWy4t6gAvva1Gdq1kLd9aBw0gU3W9oQeb6wEB3dReD1vvtQwsqsN
6/SH2uxKt5akcbXnVzp+9JJ29p0ZC77lwjBL3Bv8+/mQV5lVc/fFTSh0TSZPsKQlkXtCMqzjinaj
V6RQ0UCi8uY/QtGCvAiGPJUV+KzQZEYX7aH2FS0aTV8VZdsbnx9ZZr4faPOMQzAnF+b4Xh0YfrWu
TerDieD5dnTjsj8iBIr6hFf2FmvYAgdKUJP3xuby2j+9njM6QFx9Js7AlEEyypqguAQ84oaysRAG
+LvKAbWMLJkYy13NVRnIlTtrYepYSlMIkUsoF/mt1X2u2AoPPkh7SdPfAkN2TqMY0OIYrWC+bFCG
7oSxxK/poQCSl1l8BVOivvLKB1jZAEChfMWG71jdDaRanMRrioxHYzW43Pwod3AhzwXAgBYJ2WDt
ttAvhGCcdW+qxYl0dUScA0l7kIx2b+YTZHbbWzitPKRu8bfQxcIh/mkoJaCIaFt+DBpDpBcNDK5r
HuyVgd70YfEWvcLSq5V40A2e3kY6YGqqzGn5FdJohZTl1VfsF+DhpFOCjUYSHQakzjKc1lvssN01
vRxjaVYA0mzHdVfCzYM28lsbLcKb6VYgEDOybCRtwUdwuOg8j0PDqP4bduzTXl3gweKruCcP8H9E
TRmpgDllGtBlubwBx49z2wISR3eA6bFvq7s3tc/qXGhpT0uw0eKiWfbukv9WxWmuas+nhbtXh/M6
Uhk/Ych6UM2Jdy5gEdGTEafbVLG8NiFyUDkGQLoiqFH2+danYjGNN4bAb+1UvxCuk6iBrKGMayVq
iWOr5PqfneSs0YvshzJTCixgkmHCehGhDGT4lI+FRQuJotF8uzn2G9z8K3gCOzOI4vY6u8485vSm
S70JrwqTwn9r6/fM1xWHu4BBowTHBP6fwIzZ1Kcfd6LxoRZ7FYLRdvO367FELcrG+VidHmPd3gC2
ar9hN9fhA7YgyY3yRRNyt5fQWqRGm3yPuLtDTrElqP35Va0JOJokSmpmNGWmEq5Hj/Yiq64L+F+C
ePqiH9moOBW2HUpQg5KzvKZJsEaj3XWe+2kC0vuV0zwYb1NiliK2EmxSj8+k3up+9FNV3+TNUZc/
DdS5RfrPlg7No/HBudyr07yZo5cjU297f3o1YVzkZ72fQuCr7+C9tp8y7LZxvx8wFRtKxbPTLIoR
ofbKNYZu4cSbCnxRRh1Q7Bqp/v94SHQEKraO6fcilAn1c1r9u/38TjOWdgdf9Z0AmIOURtFBH1Yu
JlQJMPn0TAqnAMHs8sWr+W2Aq138TbWyGxB/5czWgXS9VJ16pYHUVZf/id/FUvlFrP3LzVtaO4yO
77jUog2OYtHJm8tU2CT8nOqLS8XeeGVY+AnKhWQiulRYshCamMSusnPpmsZx48ApY4Qch42TGIMj
D2QUfqEyGpPo7XbAc9DPv8WS4pU49PBF4c8kA98Fmjphid67Dteo4DYCX5o7NiVjSKQDsWx7ykhW
q6pHe1X9xstQ0RunxfdoRrdABHw4T6wh/Ha8X50SmwDUc44+kvfTVDyRIVezd87w6tHa7N9aAt5E
kHLvw3pNOtxpinTAjhfyoHlbVDF1FThu7go1SaRk27tHHAH6TicOp6Jlo4COsu50DMrF4SRY9V1V
I46I8hjGMpYC0dedFGPGlkt5dsl8oTCAPvKPyLnLq9eGqbANXQrDnuQ+a1s8Icrgxm9cud4ILMcE
vyCrVumQ2YePWMh0bHBLkYeMm3myv4hEYBdDZVLMlglbXQFIc4n/0+GJk+B4ImIuyE0nqyDlS3LS
iTAEwJxuvYvbTcSrJm3ayNPb7sS+Qh/SBgQV6ua3hvEjbPJm+fbHYwz1sWMrBLjAUYKET9a8MrxI
Rbz7s44jFIT1RmclbYZgShn1S1bkBLWX5u55ygTL1K/emsyWAf1ib9fA9yKqUcCAGLqm/FFbWst9
YJ/QFlBHFtWgfQFkEzMMRvP+j174gmrufj+fXI7tf+6G4foxzDLMVri3TjURpHYxDU2fZ4V+eGj4
BwuXgFWnghZQ834QljCTX7X2Po/41OLJbxySl6OE+3WWAarJdq7bVUV5mZ+BLlId2gXxxtd/b9VL
kU/tEppXd49jl2k6tT5XAgPDV1rrqFYpDvd7rj8t+J1Nj8u77/F60IG/AaNfjVq6S4u9vjh4UYgo
6vmFZ2xOVOzwFQQkE1bOg1dlu6nCMBDnOKzhJStzXP7nqZ16WKxyrVU9X1GPZoLPhNAVK37/x/kN
8K3GkliIBsaMJW7aW+QC71RHRkw8YkalfAg/RkoebJMazN0mPRvhGxD3NjlLT+6rGmxcTLlXkO+a
gWCN4w6xCtZ2P8gTklq5Imu61FTVy8pmRCgl8cLZ4BCh3gn+3stk5naC6xN0gHs1dEf8PHrOw5/s
oM+VjXaJlqEtg4VC4t0JNAtl8iMdN1+sD0VDSWjXaug6lxRu5cF4JTQBHeWp86udAgZRy7XZ4rEY
64V417POJypMW4+pgzNPaQqQanQIaZE0kP4qiCjnF2CVCc5glKPI9YfOfIX1s4GhmUcxFaXNwtev
PDH8EdN4Q1Q/eY1JtS2exIe5Pts5ddfThtQUnmBStzZCcurlZfkFVn7f6APH1qdaawnhL3l8BWgR
18w/hIixxsFSdcYECWnj8yc6fJ1HlAh1RoemD6AZALFMo2to8o8Yab814sJ6VaennGhLGHg38CqC
eLyv2R6EHKJCJu4X0c3VMiXHLaMrVkazrG4VjoTv5mIiP/PRWWE5EMT6/lsXWyIzZ/7IN+lBFv6E
21PAmznxwsIJw6WsNtcANHvJfRLmF4wkvDLTQxAYNhGl88PHvCdDav/IGjgfZN2u81mA1zCBYFTt
vuxkun0Srwj+bByKbdJy7805USCoXEC2vvw9u434Q7okm1eq36wMv12lYXTOMkPYBVPtoeM88/tP
zak6XQqunHlGcGmy32UCSsglveHAiE9BCCmrsndlqdJMmIlhAO2++vI5QNXCA7xQ93V6n9xXuCCm
1CYwtnY8ekzfeTRUYxs5gXOYCDISZLCAIHq4bNUIhe8/DWXqR67IqxjI7A2nc2mVIbE3xj/8Eqlz
eRbBxe7TyGPLRqSOEBD3wbcynFu2KXDA7iyvYv1iX4WMcgG35caPKPByQ+Xh1PyF2vK2NXpDN/4Q
LOPWuhso2hMTUwM0ZlJGmG8qnZJEHcBI93qnFnDp5asTaR4nuPkCezIPu6FfQWEng0TLRCgQb6ty
Aho3DqsUP7MZX/Z/gDASpWuha5OyqnWyi3mru5c4ELck7Pco5eVJuq9NcZr5+/BAIgA6UYNxQ7VY
gc5u5G9M6GWSvyIxDMQf9g1L7mRqUXmrYItl4WI/kVgxTaFH4hktYhNJCEExoCcV8CKj3EfgO8bi
qUxawdd3mue9x8Tim9jc37XYXnQLFQ6vjoDLISUhuyxC84P1s2G8LILWcoxtVJtC8d8DMBB1PVox
oPRwU9Iai5rXNm+wF4jglzlC2C9qzqy2eaYqTdgMMCyzkU/wfzfvoifGZ3nKKKFDgpxS2SzqfsQU
IfwYWLRdeXeofFdq2ejGbH3AQaXNg2X1lZSwkA6buZi8aI4roJBd2B9JTym3HTIoO7KHgA1vdZIQ
wmOarwGpv7voXtb/aGj1MQv1TROsoG1i4b97eIGtN1en94fq0EgRGcQ5/QDFB0kyoSFPq0RgMIE8
itOhFRP442jAMbgPhHvXE3tuOdtbaU/cWq0mX2cfV32uQW1qrNOzfj6yO/1MpF5Rcu4MFh9oViQc
Ga/KLb53xRR5IPlEDxMZ33ZZjlMsphgSGJqnfwd0o3Ch/vNasoEh6pu9sOPhnHPxm19RmiBgaJZ9
IrnNUersWIL0PTrwZrrzMO5frN4gfTutq9Q2UYcT57B1hj4NHKlNpFtSTyKmwgADUhdFjSPeuPPT
0u0Qrt2f2WP4zHGQlRjM+i2tBtKWo4sUDIslNob6m5TS/o+/QsyIVoZD73qH0fbHS0UqhdSgjYTq
XYl4oqvFRnHLhUQvYcJf/wlij3PerxQNandXKOsVkBhW9KlJhOniYX2eTx+vaUUAZCs6IgIU1YEQ
1lt4MNqovT6DoBpWm7oNeLRwsVyPd+dh5+NHgg3nTUOpLxI7D8mlUTXLIqFuR00WBgVhJvUEjiB8
JSi3deN0SYXY6hdzKjFBajViJNVzJrRQQCAFIA3/duzcc6g7ake5q2SCAkldNtq5QiB3C5EqmHHZ
ORVt54a3upiAplV/z2S1Yqs0K0jzBKZACu299HqyQCllig1PbyIW/ED0godOweDY1Efqxxe/a1+G
AaaESSkNpuI9+lz8J90S/2vh87tMFiBGY/CxQ1JejTxn2G45/LkPQA467a7TanvtjDKGb33+BGT/
vC7Qr0RTfcZPjaZYhp3InwHenPJlOBSAzUCpqBroB61xY+HGPAdYzeVDIjr8eB85qc+h9rwlDiUi
wx7BzdP1g62dV10WQaM2NQPpWxL2WQC4izF7rvGiKU86qn6gFtgpidCypOt6v1846i78T+kpjEoS
tjuNahkJkZHn8R3gBerNYgZR0qatbmG/NyRBTPvRQapL0eHG5lhk6H8thAhgBi/rQgp3NS+5O4cU
Cdk6CkcmlAkN9FRlBq14/rG2izvlcdi+uFkrLoEPfiEiEfywt5mH0uB07NFYvVndCkx/ZLCyYxvu
0j1F1Ss5KnMT44KNUgQbpIOqpGK+PxevrzzBow2rFeP2NGdv4vNpi985ynQxlC93G3eZpJiVVw0W
uLcv5v7ZY95t6UBFRY4yN8UPQhJAQ8M6T0TxxQ48lrt1/UhquXeJKdQPxPYKiZVjS3EOKDVmOMaq
HzeZ/i6/tYELZFiiOORbTFE5zwYTGzp4p5zCoSvadIjdSWj4+FLchtQPHYBVPbBpcGxfw2W1QYWP
dPYpahwn7W5CM5Ta3nmohItky93f70zKmvXDObaFvfg6ChEiD2GZsZgxY8eqcsL3j6UILNV/USCe
Broff6TwDP6Kisnj7g/vqYiMzb6hpTRiD7gPSQHsY5e3q6Jz0kFwZcpL7KuthhAtpabSrHw8TZ7n
ll/pJ3Rj3jpjwnVymBL4wiMiTwOsQ7RMmvnzS10T3s3tXtZoFGQRzn2ezqff0oHJxVyvnotjm+3C
2pYFIGZfM73h4SQOhTAfR9CBHZWpFj/HNhZ4KF44Db3mCJau2X2E/+yLVk5xS+lChfZ/GCF+r59u
RQlU5egFMAtj5yBY4Qg/2x8nCpFq0m6O5Q1ee9zFWaIDZu5XL/530r0kns6Wa6XuvJHnv1ecIDAB
RW1oGDpKJ1PznUnJ2iJKsVgwBCXcyY53/6WIUEFyLxOpEcqqzXokTTCfCK+yLYyMQMpYIXM8zzdr
AB0YEgE7yNoEngkG5GOHJ+2bUtYdy1gPcW0s/EUCKYc3QGW+/i+61P4hxqaOxYD7TFgOm9lnnynD
ngY5brhteVjejCiT7O3WnOciIvWvdP2DqSm/EhWYooshoYoxVnhMGDriht+TEC4cLdw0OC4fESYI
FXtAzm0ZMdABe1Iq9XMagpO3pn+SbkS3aVxQlReE7EqICuX5zfJXndygpSZS30Iltubb+nsXkJy5
v74bIT5YV2bUqMyM/2JNlxnUDkujjYuaRcOWlzEGq4XtcknRFfy2uEo3PvGRih4dhD/NwvvxdHhT
BHoV/kYthnYLsnREkDwjOdrTttcORv30/RM4gWGsp8Pj3VFGT1V4cATE7qsOe8JMJ5wNBIHs8bz9
yqye1D04k4HpK1PITrrayb4/wj6FyHOg51deKG4oFR2JUv7P8mc30kvCkI0naUrRH23mzjGkqW/c
lpjGNZpHPWes/M/cqDXkkLvtyDvs+cI1FsIUTBpqyArt3D8/D54pJXcvab1wry8989PePpjbVcFm
nPXX30N3m3CRTzcYrsomO1cnOjAEO2SRYmxgGXk4WaDqVPycO5DXfTZ6AvLZhqOGGzJ8qh0fnJfD
jHXwnq1ZU6ZSPa/6s3E0HMNF95S3JsZ8BzFBBXd+esOPQYflgyo0gGKlczkB4wetPorZTrPXnry6
S1Dj2mJUo2luYtCXIuH3TqyqZf2LpPhcmRVbXaS9B171uKG/A+750pFLepJveGG1NNr2alhfvJbt
0vzhFLvrPHkytWgZRwa5r7Tcm/haMOvx7K3NfnNWrhX6gQlPW1ILPMvPH+3XzCDY83LuJzg+Ur7m
/xqcw5ru3VjO3w2T51oKHubDY7/gK0I9fm95DXhnWCWco0ugt8du+qE60Vsy3ZWzIP9PWMm+CMAX
WC9tzUqN3fz0LQoJ2eZLRQXSCX3JYgN6D6eBmbPTohrl/j63P4Ut9LqijGRJ2aEs25WLxgMYS4xa
ANrnYQ//ZEcLa++zzrMwOeG0FDxByTXuEgQaPAhPSVCHkj7JxWzkYJ5SZxJRhPz+sCoPp50VeFPo
Gxr5ZErFhLUGkNBKfToAA+H5swRXVHPB4lOHCBaSYWKBmuR7mFDRMWdHrf4xMq4kHNmRuCbbcow6
fGjuRnTCaL/PrP32/TtvDTrgvDy/OM5q6nb0A0pxT812QalPdy8jCGQjShrTv8y2T5FYXwmWQXx8
5mcTdmzC+MYeXYPiN/ZoVNR1BPhq2OsYFGRE7s8RFPYGW7Mq3y37Y1o1rfG/+cRiH+79NCeZKTID
edKLaDnY21pQsxplTPP0voFFX8uboHQpPtYeBQqMTGZpkFJomWt7sanZGYuOM++tt3uxH7ZzTxdt
9td6N72hAHRcXT4IjWRlbbCiHRn91UgSbOwOK1900PJpBeZVq8LSFlUbdoRoMn9+mrhT6C1/0qCl
wPFrpH0iZvgCflBUFQSphxP35InbEahkY1QPpHSqkBkmvk1fFXSgrmKwEbkK7eUP3E4SaxIaihz+
k1HwrN0KpusDxTNePfBiUQAKKXO2hO9/OxTvWxfa4ReCkcuuWovdkdOd4Fu42zvJu+hWdExKAJhd
PPk5ePK6Jxly1vWhDP1GK8mSdFlp5DaQwvikBG+d0p+ns0VlTthxAc7nRMTewzuF5htHVG7glYpH
H00lDSf6c+kBNuJwmgzyL9Mpv7SVDAkOeXHaCX7vciGaL+UGYhxoe74nRDkqAWgCr41HAD6TI2XR
CtDzUJRFbUb1aFFoOkijbji+pggKuRZ6EiWh6C9YjjbMupMN41zhJZXttb7W/oHOgAIRn5u2ij0A
0P+/keWK/pyCjZbnqUe3q5Ncm9Yka27hqnxiX4Xoiu17gZR6tIymFb/SbL5SeGN/nB1b5Gnt0Q9e
aoBlaMTqGrth2EKTKyONmWPTjMDXtvnI2vVTarJdI3s2IxaaqH88ft/ni167qeVHUxels9IAe1ML
tPeg5aH+WreWPs+mqVNHYkXi+NU9TuzCzYDyOBOA9VDcLXanbcbhZUJsyxmQxI6fcdzIcb2exN9C
I0kCRHkMh9e6GTgFUo91dV/J4nSS2jH/rGU0CGKBLmNQT6VNnICMSg0z8zEPjgkMWnplNQfxHdIh
nucISRA0MbE4fTwEIDn8J3n1SWiETG7oWgWpwPHarbAhKmdgHhJJ3iENv23/mts3IemwftY7Tq9g
JhHw4h+dA1C0g9onlViBSSLk0ruz9jz+VSjOgS4y/IDMvAJkTYzZaFeBnlqK3Mo6tSgE+399khkr
CIIEPUnw//t7jwHmtlYAU8/yStUy1zU36RzxH1hh3vap3NzghqFuI8ZDzLGJV7PyejBSn4eQYJpw
5puG3xs7ri1Pp78DWX0ghxjITtjoWzsOYYMc0olX7PlC3r6BqQ42BVflornWrGUOK6VSFNKg+k/5
3VErG33kWRGjpf71qIpi3rVFPTfzwHYDk617sSAjTV34q9qlWBPz+mCbujDV9qWfSo+jpvFqASKL
DgPyncJDIASbU25Xb7OFEneoT8D7KCyuNMHovQOyFyLqnEsblkaYYbexAJ23+ZmvK3AIFqtlQXgc
3aM1nGTfoMgwPArzJqTq8QIVBBkfiMPP0bSgq7OOzvezwtKYoztKr1PwRCDJpddJ/eZ8EESHY+Xi
3DDprW99LBxra6X2GcwhI/sZIdBHTCn3lpglXEqVYgq7khyisN743zckCRCb14DUrxnPVcQzOjVP
38MAQv+MoimSkWlImMYsLg/PV5mpjIuHk2wmvghDp4r5uwYAX7R4WTrAKbmaSyNKuh6IS2p1E4LB
cBMWdmQT3R7sFC8/G4UBkP4BkfE5YMPAvlvYZSH/3NDCnS92KSVHuBkHz82AJz3JwYkmxOPr371+
aZp0CWMVFWhCHT3w5gQQ3a7ZR+SXkdnzFoqnNrDxjve4R+nIKLzLXMGRAnarNP0rGComn8bte59/
nCBxivIeRDTq5XtZRNJXfgIqt3xuN/emY/NLinTmsY1le9VdKfu1zkdYFPNxLsiLBhHXzct+8fTn
mPTvW3Y8S0UwWCKmYoW+lrKDcxH1YeLyauj7jnsByzXCuLHqVISnodA3Zd7lV3qFkfvC0Okn7NZC
kOwTOsCXj94RIvisjEdzRqjiNhuk34q4/97ZGzZHJMyltoNFq4QmUFVMJJjxFYutSnuwP0iC1g3F
oithVJzevzQp2RQ6HaY0C9zq/7MbFAzjDge6/WMqUib5W0JdBj+VBCsXwZlHhkSDM68aw0gFLRKN
od38nEaXyy4ghuUSfGdy46/AafhJUyoQHnPXbnRx84OiJf3goXowZyVXbf5yZKvyeO9Flv0oK/6M
buFbGmwIYlHxMSgjQYphkFZYs4/2a/X00abViH0DRoQL3lhNYr2AhYSyxlMT8LY+t6gpN/Umz844
cvsyVW4ZyuZTUXBKuTS5+xxDCC0Vnb9GecmlwmaSDs7D0Ssb9PtRb/f9xkXHZEGXCrEsXh+bmuqw
mQWVffY/pLbtp7b3ak1IuRG7ByRlr6kPR8kxreiVfTJBXdMEZjfOEGrdev7a+jQLA53Am63tbPVu
HRHfuSLKPoUN/jn9zy3R6dWyi7RaLxAw3uSf9+GjLrIFQhDHwtv4kL7DKvEEcr2NkKMgCgQazXDs
AEZ4MEcsE3CbrMJytd60mBmUwe95DoGZhQOEbi4xoY2Famg2Ot//IfITdTs/j0omSYB3tN3dYnKO
/4FOWKqk+QJiLzGjjQkrsFq9jXpfr8SncGJbQ8vkA+0x22L/FnBOZRGl/vJprxU2+Wve+0H67rWn
3usX2I7KcfGtM/UcL95saEzLbvtwo7TdSTshQu2YUZipaeivUlE/ff0og4oE2Ol1kxXqrHhmICen
xGRb8NwM/SgGCt22h2fn5tTheTXdg6KsN+r0DUou73uT9F0v9B3+HpPJKCaQ+7mAQw7G9ganh0R+
v2zEOzXLb/MbZ5NU6oevGsYW99x2XiyYpqI5ggeiiSRQ4+g/GRFyEiOtFxbGl9ELM6YzG/uwclyH
hOYDsLAL3Rk6CLv2JulADfZxdBUxL2mibr5Y76DlWoH5HySfa8JfJZgqqZ8YCa3He6Rjx7AzCwJb
fNHx3RJAyZ+q1/fXSJiYt5f7gZrmGSf4hbHpDwDdGdv6lVXElw2TP71H8qt+ZxbiCJ0fac1j4feg
YqlqhcHsRNFoNqCHF3mYNrdsxkfR4xUQj/LeHw1ExG7vtYxB6EV845GPCdYKTqbo4ashvS/H3Ga+
+N0S6VXzfgYPq5pg8uy5mdLMO6GCb08ljKfFYxnS6xRMb4s7HPsilzI0dOcK8ALPmWwCGxalhFUo
o8bxWqbVXTxonR5LMFmrvM08XTdrLgfQ88Wj8R1kp625L63W/h1ibhyueAwTzren7xrgsio1b8FI
zc16ZSiYCKEjTSU+AvQGgcSrBfN7SIeNxumMm58IPgHG5BtKOy+Dwfsjqi8d2reqxgUIu+9IUp9E
uLFlwWPC+jQGxv4QlvEBgeoqcpOucsdOF2KBQaq/GFcZeuu5nw3JwDWsx1xgaM0iO/yzT6b383dc
ykYOSpvGcFlWwxRIcSQ/SUonfSFie56m72Qu2TUJ98BR5nE5G+Azt6Jnw6GWQSXlKXTyDgDnchTn
yLAhiid7qbEEXi01Q9jqHB+IbYTA8m//4GK60oods6dGhKG06QEz4Mnijy6xDF55KrZ2J80UYXOW
M0XDglMm2kSafgFVTL2Vq2b3bQa6bObe7UtCsP9l+B1n+qTkSF8E7SvxwCInyoxBn+nhPm+Ltkuy
fuhbP1BHGu4C62jraoV0FqKdNm/6Wujm+P889ZOS0ZdTbSGcu2jVRS6INJ5rf3iZ2WpEE/HlPIB6
TiTqOpBiIxYVmDYxRHzVBMuuZsqwXUHCf9gsJuhPoXCwXEAuGXT3laE9Se9VNoxmRr+xLYd7cIsi
CqBX7wXtZlrf/Cq6BvKXf+ThdwEiA+tDxnwZEocuUfG6OymSQxQkD6aqA833y6z/IOjUe3meyViB
xpf1KPytVffJ2alvHlEn2DAkTMZvzXC0mMTe17jEL94cJ9NWwL5ZG4z6ITb5N9npcAtykG7IvzpI
NOBPk04ItplcdMyERs1PHyde0fvUeR2O9SOkuxL/uURFIkBFudsefbCdrLSxgUm1cMnTFsm5ngiT
+aXpE7ojNb3sav/8A5heK0LvYxVOJv3gUwSrmhnolPxUlzXzVSWKfeohZVZTypLIZAOhn7KfJKNn
UodNTVOwLgMjb7DvQWCaX1uP/+2xEPMUWZcq3L/o77Gze8Lv5eb7G1YMCTa0dkoKtp+2CHqYyiHc
+7CfNp/fH2Ot3TwakzbyqF/5Alyx4NREv/ckhbrE9y6hjuZ2QsIP0gj6O8bwtv+tPIz9z9hhpTsx
21znehNYFBd65hWwTB5EGWD+ejVek1gIKtfm2fLIc0skG8nXlUlMOf2o6a5mQ0vgI1KoaqIXy0U7
epbQm5vxzv7+c40fFB2WWYXeqD9X2k2HlEdooswTs1nQt084nBaFcxstODNLfVwLsn4GjUEA65lh
thFzRg4i27iCJcQIPnf9kWnOuF5ANiUqPcZiS3qYLdhZV8JXO+iGz6oDLnSIwinxFA/+F0/tNKm4
bCLTYEE/flTfN/aFWAq4swqdVWFTOKN5OezguwbkrarHHTQgPajh5TXMVKsLbEljXZ1ot8sfETi8
ys4JsQ5QjFDkalYAcnOLATduT0gZxoh2Ltz8jL57ACWD2wqQ0LmPO7Z2+7VyJ9UcNLvf4cryoou5
6JejN5jE2+pFW/1TnYJ6l1dsBmX1EU+6fe5jha3tVs3L3DxkBODFwy4mR0RqXo2AXw6ECexanu9R
jNi0GvWpA1OjgVLCWP1Wsgbwj+THsSySRqWbpVqDoDP9hW6SsJhwVn0IdAKvV1lRzd0OLDxXhoRZ
DdYJ/x+yDc3ZgIXFOl7EmUvoHj73DP4xmZzQqbjF5aI3M+eMpa7NwvseDg8CG/5CWLjwE57VwWfG
IuLzTXoBJGIuJcnObYmdoW7pSDR2003H9Z2pDQ4yTM0xhupBqbtbch+4ub6HRhHEtK6EMqS+NUG5
tgtVqAOzoacbyU1sYvP80z1qCLMWwLPSKBDfFlxhhW1cI92vg0IaP1KrXg5DapqF+wpIH8ks66WG
9DXVM8hkHUa7ufLLkJOMjqfsJ0vmDUzZ+p7qJlQFAEOcSkfCiT3yDV7xY3TuDyCorCYgHHkdpcXf
JSrKW2vMGCvCh9f7NOfVE8wB4gBqRzt80PMYjpTZIqCaMBD6YQ51v4oPoPTHTLSPvT0YNifQrDKV
fPQbjcChNHMTyn6P+FuMjJLUlIkusJg/lhUcSW6BIjn0mqvDNzTAP5A23QOMvcteqMVlonsMFhR0
2HfWg6EoOBSnz5nEXysNH8caID+l6DMwySp6V/Q6NQm+dUuNhZ+KDahVfrZ24FXXrx8CXbRv10Ny
CbhwfhkGZWRUXiiRHsCMn5sbMM2rbh7SqToGDoV0IW5lHVKOc7DDvQ/uFfJ7DNxlUPPw8zgCOc8T
P1UZN7UiEunT+y79cNzQxbD27I9oNJfCU4yl5JOLjXUSOmn8mUr1zIT11MbuSFW6MVHW7paorvPZ
CyD8mQoXHRRj3WczlRLPYOHwIZ9+5gDID/BpjyIzLO938HQsZzbrZ2qlksomdLWYtOrOZIf7kgSM
6tlUXOJS7fdD2aTlsz97eraFjUHyifUhAmDpTMEXp9c3+DALjYJDKFNitbGbUqinQnApzIbq/IHl
frDq2rzjug9V0HXdMU7WxssexIkuvhDJ78g1jVbdd0JVck5xptyP5UFRz+lL2jmaoZVCDpW7IkDd
NpWetxX5GRGL98WYVA1AY0yvyyjx/GzfSScmc5BiwuzkTHBBy3N+9WOnUA14S4xHcintHIqa0D1j
fAFr4b5ps2JeI24AEgKNIqjCZ1TJlSTgc9695UztGMas/DJOOKGkz4MhzVv3hCoiEJYTyFYZwPCI
wzmvQ+z6K3AmyhCEqFCZF+luPAhPgvpLQM9K3Z82rN/SE8CmX1dvXSYhNVxBVhbk0L+TdizV26K2
tklxLvfTMWYqGRl3v0Wwp1aac6shnIlHeprReTGnTgURny6R0KYHa/2yyeW7naWx9GY1e4L7WbQ6
h1shAk1r9wfhtDjYOzDTgyTTR6ZYotuqLBoGEPVEi1/bVgl4VdfbBhPxy/tBikIIpNdkNB2Pyxrq
ZeBwVGNBG0ULx0ZpWuV661w8fMiE0+2Pzmvppp7zymMecuX1+tso2xDFSV3/Arl1iqoSvsMXYvnr
YWY7znSq8TnMAFpbeC9egW4z5RPMZ3BiQyZpxcFph/2d6QSX0LxA2E9pTxX6xTVO5Jz2/GludT4w
e465WJa3tKn44AcQQjlSCnnOgxVat1NGcsizgmEfFZGpIBck/bSxbXi2Z2a26zisdwQY1ETN+Ke7
y6g3Dy9J29SDFl3BBkOU0vjJBn9F2Z2yQI0gf26yNfpjtQuusN9wQYH72q2ZwB5xlTsi5OHWH8pR
LpWQsATH0qamWzAAogKbsmQdyjY8hKMzrJKeSR3Z9qHXVlcWX++9tAw8v17GPMdXG62fazi2jSk7
Kt4AB6sEqnN/d/3mpqROC8aFTP8lE94c24Vl6zl9BGwdr2PXxcOWhsqSIkoRhMTABcZDU7hjZtx2
kDAb23Ri3FxBCpUN2jfOBL9/uS0mDvwkcPvKjI7+UbX/DqafQsnVLVtrxgGYGCvJhKwaXMqY6PlT
btu8AtQQDS7MQDyGnFas8JIM666iTh0M5lMs64SM/14EapKM6Y05q3hod0NZupcywlS9lHuTLr0P
+T/66KzK5DEMwv4cen+bu1CtV5X5dKfyfXwIj8VSdaas87wGDpgA1OcD5Lomt1kqrmUTVuok3LOM
891DnEAHzSjMejF4sXqyaoTEe9bJorszsRmA2/MI0pHuTp61AmYgu88CErNsuVoGFzLn+FHPab//
szzAjCr56magAqIhwAAlhYaG07xUREzhrEru4gW2qXeVvbtoVsoAN3Befqve8DoZ0hmycPfE2oJT
jhHrt4KJ3YIlEmjyfXqPjpZh2Jj1KMFHpwhmU1Pz0WdMV15q6cbmBU4w8ziKnzhHrfohqvL+l8M0
1huQRTuPjbgGKGXiG1gxK+ZeowT2NSckssY3aBoD1JyyvULKHtIy0odmDw8Un6RTDasi59S2P2dt
yqYS2sWkDZEymYXErJXGSeu9VSS+niWlP+7xpdMFF00ZM0nk4nN4y42YgK0HjO0KKZa0bE6c0rTq
DOpEeQGYZ33DNDHOSLBsfIzN7sN0gnGGnN7v3qEgGVYwK2idXlwj+sM1bbaNLz5Hr2q6ezjDljVR
Lj+sQs2pKocQDGcNDkMJQDX5xipS56XkvVSQrpYCE/iAbTRhwYEJHHCOXyOcTM1eM1sbbTW8FdR/
WC8orhIZJwmtx8z8dYJE2nxdVV2GbkzijumdFU3ADpk9pVZFpoK6Qx7SZfa67P467uXwxWumQDml
npT/03VKbwtEA0wd2/Lo3+42rL1T0vK3+rM/KfE/jGFLoPvM2M3Bj/Y1wqAa4CWTS6t/zAVK0mlI
SFp6Gc6wzkXGXTi+W6l1USiDIZTfkMi6msyuPaxeAq1rpOCiRSEVwQ4RfCj36LUWwzWy+S7Q9ocH
jZpOasuj5tHwB+DJbatLKLXYVONA3Cwbi0A9mT8wM552l5YYSez1w7ntbWcYy2hV6dqbdN7xVS6z
9GwSFEGODibwSLK59ZEuZVBdVpHA5ZOFdeQQX4x55pSl5D1BewBY/vTQZJzeygrtOYFS8L8RgT7F
JTSDCgyS47ro2lcxGQHTlAnJUSrCSB8fCdTrfOSwUgeoqwgvmFMy75jqhiHctkGsnWLfhBqEi1qh
WkPRNrhht4lm7KKDFlkTrZndZthZ82v2lCTHbc4uyTKUFJzaab3SI16CbGVMkS3/349kHoRAXt6R
tMJXgYCBKg45lXPEyGHww9jzJ6mFiXwaoLYuG4doERT2a9y2V8OWjMTVcOaOTmwH/s955k/49E1j
G8Nu/oUnTEmMgKioFah0akbEiI2IiXaTJsXjbYU+ON2wD/UyF77SynCIE5RaQ5dttQTIt0anBBMF
PIELHtBfmbt/Ppk+uvdSJzN9ORQc4Yw9HDJv2sqvNaoTi3vBmA7z/yx1hu/c4EhmT5Nk1XhPfw73
NKH2wcxxy0o3W5Vub7Opj9P/64Lz24gZMX++rRyfTHyGU1+rWHzcVDM8XWXZyMsQp9MnxbaCNJQm
1fvgC0BpiFn3M0JL4ptpP9YpuHFZELGScS7P8omJF8TXM7HwgcyxfUH3wB0yOGY1B8L70DhBqSTF
FKuUxJW5TTVEMRlDnwfF9OWTuS6uGc4FHtZN8PgTO7f1/4AxS4TTnVqCPCzNGZyZz39QOtZRSla5
fTLjgMThdy+DTXX2BP2oFrFq4PgVSqtKycxQym2f2AD5J+35yzLA4hlifcbvptkdNEBu5Kbqp0uM
Ri0dDNjgX94e6fNUGzcSEZp9NhrRyBCemal3oD2paTbECEG78UCW965Yr9MWfh+ofVc6uRDuFZ2f
kUZY2DnXclCZyTYPI5xoGbQjKguLppkiGV6kfqeF4X70MrDN10reTtD67NJO+PRx06QhUDGQdWak
Nwn5b0qDPRMrxsTKqSzVilhhKv/1dJ7b+oPVLhfmhdr/Yp+msZO9S1hOuc1u9pyRRXIuE8nvjb0e
4MfTO6aJlpfDkqF6xTAEb8edIXXgvdc2YCPYPuO+o/d3gZVojvf8f1NhwT/EZeZHuFUHhpacRDc9
qZUlc7+CL66RBinlGFa1JYdH+AdZ5LG2zzGolB/WxfI5zsb413I6E0jXGQq27T8w+MbVujqi4mUK
B8X56EE2PpLw55/CrBuLg3YYLicPnMT5mkX/PMYNcXWwDiTy7Rq4w2jZRSWDc+nszyhtcQOgE7WD
5aY1jmUAyE6ZwxkuRgeNcL8G8B27/uwfl7wxC4sWE1MCqw7ORwEq1AlTvjzS8AAb6jPD4+uw7gS5
NUY8roCzNcZg8SgOfhmsUT9fX8+a8YX46BpbYuasxzzKk9rCLXWKa+NCUJbMYxCrwd6Gr5Ay2hNh
Lqj/BgZUiGAJz6AUM6+Fkk38L1kfgFHdWoYZbHLkm5FUAt6N2O3Sx5qR7zi4iLgLdILzIXoEMjwk
YfQ3FTb2zCGSh83ZcYEuBOA9+CbWgFzvbVGuyBeFpeaBMljTKh8JFw9xoAttpN04r0ZYvXt0IdgF
FSOmV3jUOH3UYUbL20kEl6EiqeOHRcNF2BSP7SUIy/RA9tdrUcCDZCWaftRAt1tJVyHfH31/3eip
zTUwG1GnAsbWPjkx7W/FTadZfokHTjCDb1QpwKt64NIgKP5tphQYGEp/lObt6cpUrQ0iqOYuXkKo
HoAcRw1eibddNMhRzuTvJZBo6t/KKdV/r9lTzqteGrJIeSl5osdnHNwURjzOLwmMhnFVMHM5l79p
O8tQUUvme/hLI4GwLubz68oWjwzZKA0aLpVJEFnEd7ZsAelCiZHW49auGHUw7tSE/BBcE5JwA56M
79V1338OBANVYSBhPRXwtYdhs7KuUm7ybQ+2viaYlJbgWHgmPMLisCNfAMdyiw4nD3cEnTK924Ng
dlW7xK92ERiiwM3BFwppJgnqjBmuhNoSFDZ0BTYVSJdVbSZ1Uy3imHkBiJEIA0JzkRXV7daQ87cj
ebV80Y/Qcw0OmvNiYS60g+ZVuod+PDy6hOUjONe/Q7hUF5nZsf3Qv3I5JzmKn3oMwSmapHG5aIa9
UvY6kRsJudCCC2sN4P+5v0CuHPKPQ/hGT1J5u8Ey/3wgHYlCJ7c9pW5U1c7q31wLo2H6svsIFnJG
UMUmqs0eBQINk00CSNOh1Xkf7Kht/ibbZspVXQGzbjS8tEACkwJ7N3Bryf+HVakmrcXy3VdPEa4P
WnVku2zque7BvnJyyOTZJ9/Ywan1lbhafsGuMbVY/lcLyGYTl32kgeF6tmfGZeizBJkyvE+2grj6
9gSjoorY1ItQspmr3LgN2LDFqtPnMKUPJVCd1EtFROloqP/TFau+Dq1ycqzQCOcqokyRAlVEnUpT
E/hJleKMT68aBE03g0KWuyq6saMr6ZN48MiYD4xjAGOsVSYNjwFkYcAPefeWBAedRDBPVR7KsUeW
SZGNSyWCYsmhtOAwFb1+g63hFbDHJJvaFba1Zz1mpQJuRM15/XqsubViyiJZn2/tXQYRhOl2kYj5
uepB30UrIjBDmzrPiyGfL3tiI/2a3lSoYb8mQJxpyBGBnvdCWVCxouVVqUIH2Tc7gzZ8LeYJ3xxN
jpBGi5mveiZG0xyparNRc6Qr0h3BhuyTAgWloAYTGGxpFzlZMNIEyI275Ry6VAf5HEIgcCvVrK9I
bi3f4qSCooAJOUflRnvKPiGWChzwUBxXMgPPhVx4azGD04i3D/X+YzbUry9QeaufZJkFXPnVDihk
bk9RjII2Syn/A6blFFeStwcoyJTsMwvRMRkQharBNNekd/jmLGvLOwVujoPOrOXMmvIxu6rlH3KV
MVxBlHV5f4K0E//3/3oozeSPIoq3oEiBzeOZN9GeMEVGis7Tzm+cRG6SjEol9lCEFDbY/RZopbNd
p1NYljJAIVljbm6dyBUv7CIUs2ieisIXwfWffr6RhaC915I5E/qwVgWiJoYPbpProqjtQX2I+Fvf
rHY4Nx54rMlZBsc+MqcHW9UQlIKEGLYJaRukJ3zFiLqQ+eW7IqHmDNBpiM/xZdpwbbxQOpf7vusP
nY8KD5oIp3vXEJ/1ZHD6pyGwnuFWaHhpSobVW+VWnFKsZ74SnP9dLeIEeh/YKABFlR2fhb58EIrH
DocHaipgfzNlvPpDtSar5aiD8sZ+p/7TH55NRDtZgyYyctMrUzGvWcJx1s95MX0GmHwXI0l+oCOe
ul+yDK+zXy9aBvkg70ynLRBnS71eIzPPAmSR/4EDWQh0W65BEUfBhgVKgOBmTLmXFONMNaIbMzk9
HrIni+JR1HsP7w0t1ImX+QOJhhPWKsxCSDQr24f8J8SOR5U6k2JYLftUr5TAUwCwDThIZ/9yB4t7
AjEYX252J4ZKQftoqc1mpg7qfDtkOqb/9/Gg4PCthybD7XBXSmDWtiJgUWZDgPjOrnx1vL1fH3mT
YGuQfpRiq6FGSU5r4vzPj6zDhmNvHt2RfVDgDKOpzJTIw2C4Ue4klCGTgVDit8iA+3fsX5TvEL6F
4w7SCYub3zBFq4qqwkH7xqjO4WHgYnRlk4dHzCOhQtVJDD8maTvnHAQT40KUF/dfGF91q045uZ0z
DcojggGDAZSYX4ydYIqhzep2NJE1e1JoNvN1GjO6GRbeFSu28TLxXcbDDIGWjxDemrHre2cbBgHc
GDjViABTlC3f4E1NmFpTU3ZLHGTd+f6vm5olFOLNBVTe1Wxzn7yBwhM8vUD9gXOTND1hNtyD/rAC
JOgpJCDOgQH1dPfWq46mXJl8XotJy+7/nOxbvkzdJMnG/k9h6tqMiUDy/yBb+wI3nJ7Y6DvfVsMI
j20gDplRdR6mUe5h4/TxRaSe/FuB2PkW6fzwlXBBRudlu9YvbP5BlgaXGDseyytgnC4OICXCRJ4U
N//YXELgq3sZARbiOQ3JxMrsN+lNeCFTJ3cMrgh/hazN0sJA/bvyFYDsoFGd8He+emivDy2jQBd/
Cy97khbPTUTHOQjCOQ8ofQjsw59R4zRQRCcIQkwuch7TeM+cduuWOCUU71Qj53lSvutSUR+Ry+rt
u7cED4/HIVbJHG4sepDNe4sdz2f5mehFtJsdIAxUBLlGZdSxxSQjrjWi30IQeS090YuLMObQRMnm
8TIMnJg7om6ymPUtcPXx5VvF4EW8icDs+7YjKryXOFOUPSXnahXPgREiILzgFUcjNzo2mK1ZnIm6
laHibmsU89whb8/PyUS5K+g3/4q1uCUr9RvYFHOwYjxy8vItkAsTEIBK0ffgjtB2eaFbMvdPyX+y
U1/R7R9O77+oMGWzt1c1zLAjKcRmBZR680Q7FkBIcvfYgjs3b2Fjxpw15RBaep3P6IIk3zbf/h3m
attJjWoXv79L3u0RCjuqJ2IVkOJCqvWGmysbY3JP1POryBxJRRFneAk9CVYAKnitJAB90g5BbA3t
lMW5VzFpAw8qo/TimYdryLjIdzpABSYdT5Lak8O+ATXerPsVy0vOc5tQtOH5kxUFdrJWYrhnthcd
LCrfMmWrFE0YNaARV1tewYuHPx2cjg1rI5vcopUeNEAZbzWwZkpQzkyiz6csFfnYKBoFmYZ+c1Yj
goD5aURuLxxE++u0QGZ5SMflMIxz69SE7L4JE78faDVn8m/hY3qAasZnHutujfAjZN/2BHuz3rEd
nLfY2Dhxmmv2wfayTG6lkKENeMMj/AzD2Ezew2gNYXRcvBE8GmrNpux//ffxa5kSN3rhJ80EhVqL
ZSH8kSO2jUhk6WStbht2BWHlmX4/uUHJir/L063nI/SLA1E/19fR9uPmvNn5wqxstOFyCRiqPuPl
BveUBzgB8t5N7VJqliLdBbv7EiltGWMOgsfGc/qro7Gh7FwsVyIA8dpdGX0KWgFwRfhcsGYfiJUL
r6IB0vi4lIafgLF3N/+wjsYGi7Kv1Iwvk1F4yBKMwba1OOzBh2j6tOx4EXs6zzlRMDG3ENse5uhe
0NCXZCe/OCeDsVDEn/NUYICS3QeqL4a5Xi6JIkoETM2/6qNvL6Fh8ICXryMAgJb8ke9u157Yez2v
BmXDiep+/sH44PxlYOvcKj7ZkaBK4cVrAgGPXBWpNA15/KgQdH7swzqqtOyYyJPFXWjbhk8x7JJ/
3waCZnamqntb3ZmAjcUErZJ9NCxMdQ81rBpbbZAUIM/bXoGfm2ZyXZ6WNB6YsgSMD6BetPY90Ktg
iAq/sd6HkhwbFBYDKI5UM5R+agrg+GwG9Q5hDFYEcpUdQQ3Sd4B3CIrxBMneOdOH0km3rDf+KGB0
zduS6BzCifMWQfOLf+Y7X+xz1kw9gxnjSNpdIA1N8K6mNRCyRb2t/q5NW2jazmhrcm58vPn1dDff
H6pLMv3PIUiWprSDtGLaKF4u2xuhJ0wEEAiAvWXEox/mXcB9wplifUT5CuuZVGXcCyKeUXOwfe4i
b7NJmY5saSYNrXpc4e9SgT8JWGn2CMG/TbhOQPPLqpF2rwIv64y0c/x9gFECoxSg8kwZIKakuWKP
lslkYVBjdhmT16Mo2sYDGOcQkzAhmJ+vlqwpW4PjtpK0nOWhoQbsq96tztRhpeDJ0KTrkjXJSjf2
km9AxxsjN4sgqGto9V+PIjpPGdkVvTuPFBxL+WWE/hj+KdWqDeMdTzIOn3OXWieNjXesWhfbLukD
zKz+eH7XL31BkG/UkhcL3UMScI1685lXgbH+UttUsjB6wVRV4QvTSMTny3g01q+LHO7bcIVdxf37
ZaOpyovajvOwQvifuOS+H3Da716eZl7d7NXMOYtQDsNVVS2NLt9QEw4OoH3foKPx47ljYyHTE1yG
L/Arj2w9jRu9PfmawFRU2MH8gR3pkg7mHE5m7xPLcTLsEUEQ2Xz0Ogcxe+Dycnl0nXvPaPlButBw
eMxfgN3CHN37Xz3jN7Or3Mpr9eE3yMxm1Z+buOxLvRK0SA5Aj2IqXh03wqlX6LGhb4IlwJsJNNPj
0qzxc7B35eCzgaoI3cPVeA5+8Jhsl/5fKH19GMCFM/SCS1qrJd4kH+AcmBTh0HmRn6WKRK81OeBH
pX7q5cr2/iLPv3OraFXbG7ctaJh+tXp20A2NuFSAbtTYhUYadLgF4Uv3CKGaPXI8R4q+6OsEIbNe
OJ7hcA9heMuX1z4GuIDyfG9MMC0Tnqem2272u+z2VfqH/cqJNC9/T+6/ZynqgWQ2kudRG7wEcmAY
YvTf3TtiJVHzJHmRLHYpc0kIOV1AABPJ3n5awPS34PSHU3azhW93xSOOVvCByf7vMg55/ZiY8/pn
M6V1s2p9akRetNKR5SPEUZOkG+A1gCY8s8XS2w8EyGoUco1nPMbkCZ4T3rk8IT6sDYnEKDxOfHLb
0JNN/gqaEbzwSdCW6Xkn80PpPD6Oi10fObxjAGWed5zNVIMYYTTigTGGubq9tBEFaNmSp8WkGV+C
hyqM7ILvO1FtlbA/yNfiS+se35SfHBselANAi/TET0Nm8AShnrnD1FBMf924mmh/Rsy9UFiVmjeQ
9T46GaTb4S/9+MWmlsccOLeaikPISoBOXjokDLR5BJ0Atzde/eFowlekU8TT/ubfpspRHvmw760o
XC8nXSzaVemBJPIavI+EGKBz+FsXoQ05jYUp0dYLbBViDaaxF6Hxlii1J24mrTl2vS66cb9Ekz2w
QoyAC/do6WDIbxVm9LN2k8Eyrxg/7tTqcFs0mIDso0FQXr2k0oCgm5gl8l+doWAHN5DbF9jeM/jZ
xSPzOHRcl4GAmDEnxK2fsvw54Aj+MEV1a97K/BMggFNsumNoTSXl0tK1Fl0GGWOxV/sSF1zyB6a2
faoOnxyh1sDZAzCM3WCczZIF2hI5g6VAKi5PczejMY0aGVKY/NLIrNKXedD0Oi13TK84OWZz1i61
/SiCw1GMVlCQnzQP7V4LG+rb7E+ffKujt1X8fL3k464J4OStsOICh/9J536bcW9T/eSIChnA7VuR
NylrHmeZcZ0x8MmOnklG6WHOntYnzLbXVE4lUcCa7arVwe94nHq9lgiwVYK98daD9WqKW7KdDx0K
A1dtFHLtcgaPsD9jP2xNa6LNUDGYkENOKuWK27uQEtL0yvgxH3Fz4oevRjWfV9BlK/1Q4Kxk61u9
yRuRii+SReR0Mw8B4rnu93W0u77day2ZdAro2Vz8Dj08gScmuN/400IDn3JA1vxnyqqUB0nm1G6S
ML6ShM+bZRkwfwaev/XOv3LNrNgwAgU77xG8YYqWbOk6707TZdUpROy2SxRqLmF4VE/u8OlOMB8U
yTO0LjkaSkKn/whBQZbWkzC2d1rssFeHlDqQzUPw2LagZ9t32OY7ArFdAV/p3auHfNP/v52z3Z8d
vjp+ETEF8a/CMvEKCv+r5VtmVXjdllCIjvCsF+ugoZHdO92qi/8ENeabSw8yEaInVy+bIcBJJ3cj
J4vtsyXgp6i7fNl87mu/tIMjGlGyiDCFrQFPG95MXokJos4jX4I9Rv8WLWhdGUlk4H2MjPC0toUx
TDuMiCnDSbDF1Wscve44/FlkisP4nYVTY417DE8E8lXa3QezhAUjSLVAsTgSF2pcYEygC5jePEMy
JBIxGh3kKGD/NRVY45l5KQxYoETG0rh26s6rkVa79PgPKx6ozfVdxPi4cft4e1P0Tw9prx3QLISl
BwzGD7+crCyy39eeX9AvMyCTufCsW/lHXcwfI5hUFgwG5LbQJecEwmrdupYeVRJflKsgX2uSMrMl
crwnvCL7r/9uT+K/4TFpX+kxfu75V5ipnA2/U0TNv8TB4YQ3i70IPlme6+7OI4xrSqPkKOyGqaOx
1g72umDqS3B4dURltobJex4XTYwoJfniHEorlj3693hgIvMJYi+/pegEme0cEdHwbO4i8NClKJTj
C1rKuBvII0WU71B8HvMxw5j61sSw2Y9XzF2jJfPeC+pdr+E6frIQIBkVq+l0+9HtAYswDYAiDskb
XM8OzmpR+uhghM37/9fvYq83NLKkMsS9xJBaZjhcYDguyec1xyLy6sf+EXx7TzHepbGLqkV4Io1a
h+lz223fecz5lfATUefbFY3UiVVMhYWGzntCrAhGCr4YvzI/D2DSBEFGrQ2YTQubzM/Of6iJjDKo
6k4V94yQgKNAgiPpyCY24O9MBYSyCvMApjFFTJgM+nMb0u+TSUy563zuWK5/DJPIbAzxnHU9gpa1
3oukQgWNXweL/vp8A3pRRYw8fBhyiHXV9Artm2sGLQ3c9mwaxjtiIz62mLY00D0y2NIbxxofGDjL
jKNP4+3ViLuMC8hD6avyMXZLVI0HvuPxY0TkgbUK+jPGDZQKCFGqRyxQUV3nC6mHuEAY1IhHljMc
4zs12+goGN1XgZ7jLWkJJ/D/8zvOGkuGoEoTTW5V2nNVJwx9IMHX0Ep+0lF3nU8S3kTbmC/Qtj2C
cFKk9qIcMlSFsyxFZ926Dw10gUEyOiXcigaZYdm1tjXyDp7wmuvr/HaPYJLVqXWu3InnaXn/GxdY
y9yXTMnwMLfH1y3j/Ffathl8Q5H6Yg+LUybeVbiyByUHZvNDybuj2A2Em3M3+K8m49lX2J99KJmj
vm8GMPtw3EZaHC4lm/tz0Pv2O/Jlw4RsY5D9m9OqiXYygmfWptwNXiHDIqqoDKyPay3L5SJRIEx+
Btj+9Zlk1+HDtWNBJvDFOGzlBQTHG7TH5cxCVFEK56W76b3xJ9QBA5xVOEzsl95+Q+aaAeCplXAl
K/1jAuNyZnP9ESjb12JMsSEoAz8s5WpQrA8Mp9GyR++pU+eP2YVTiC4g9xw/oBwdub4wN4oLfvBT
aPaRIcKzrfaFTM8eXQPspPZldLbdu7Ny1SD/weGWStne/VD9HInkIfdX2LZuUoJFrxQIxNgwoqfv
Y80HZhwAMEOhScyWDsBJ8heOh/JkB8Puqu+qKwx4EXeUxDHNuwhsjYXNYZXDfSwtbZaSptAlzsx5
z4f+GshBkvJ7qxsX0poZOLXEoob43I4yV1nXCiCqU3p7mcOAQTlZoEHDoL+u6U6sELstomHrqcs4
MKgFygXiY3xqogLhTg0P/bVNWtPWPs4loeGOEA0bjJZKKL/0mM71/RwOHZOhDffaV2A7NfTM7ic1
Gvpa9ftXGtKGWRNTNlf7z6pPrzAdH2kuvZfJXFWUPvES0v/QS0RL4Pv+CAucuRBxPZhqtHSZRxsF
2v2c8BLP1/QJTszDHP7TiY7louqFCuRyV+UG0qzi3cNzz8BWhVZEgBbqLj1mbkJa6rzEFBVoctK3
44kOekc83GrIRhSPRkw4Vn6cjcZeeVi8DwXW9GFcYUrL8p08NQu29QJHYxh7rkizuFf87IsZh0A+
I5tTCoBkfDnMvC1/BZeZgot9P9DU3lf1kGsTbjbNwYmgDJMXySL+KSzXE28/iErIraxBLlk+iH0X
mOXQTkT8IRsM7Z9XiCwT9o1JxKiiP3zCI1cgy6KH2dKAJ8g1G3QLUmKYbhupOF8dWgcTE12nT8F5
iUsDeWXctZIuj7aQrSQH/muQINCKInqfdkWOB8A3ufHm2MW/RGLJYpSaAr1cXzGnmBC8weY9VfJL
J0pa+NeioOBggUA7q2L8PtPT98u0MzjHbm0LeJjNflsI/CpLPRAJDjfOxcupXZ51NwZpdljGp8Xa
me04S8oC+oP9jpVrGW/LwmLn/kvtO6U3VoKDIElz7iZxHqIp1zUAtL/QrKQ/tnKT2nwGuWDOgcC8
lnWMidqiuZspvJn5Dn0MbGONyeGS/G4ayf1OhKXSvUfI5mfqJXcoEacIr4E/VXYkUGgwL3gRRLp9
X6t4pwlS66ZQhOSrEMp572vA8wuKyZ9pbQ6WD1aw6j8cJB16z0yZ54gRWuOCUfZxcrSem8eYRoqi
bCAhbaz0tsu/vvwMNJ9YYnPQF4aaLSjlu32iuaxuVIYxKb5LNl4jwGqmmTa0vNR6QGcEPmrlyS/5
XPycxK8HvBkpNDfpfJKw3K2qphs7zp9vVFsxi05ekDu96YteIWZuscStksLAq2d7wFrfCFpPubCR
suP6ePAbE8GoJZ6EEAD4LknPH8ca/IVJlp1tRIPB3HDqnd4frp7/Cy0Y45JFwBa/3p2kOIR62Z9Q
TXYKabExhvH3SbB4rIwWKJLnmSD2JsbzX3fRAMt9QyIKQu3+qDTgBNsM91pSDW6PIdz8FqLg/BDE
NmFJE6jyEOnmsJ7zs54snsGWmelkoD98YT5QClQMYd6g/vfjdv0NEwQC+527ONFUCOf3YhuNKLXL
i2tZAjnX7PgsaQoIurjiVmkuVF1plZXzzXmEVM6ZhS9bPLFAywQaKWr1ajFKZheDONz2zFAsxgD9
pH54CMtq4WYmOQHXoGEvOl+VAi4pS71thc66eAxm2tk9Fk1MZnpgjvxb15dRlX4H88W+oVV0ZG3Z
5ZiAeP4Uh4hL7+ikhRvncR6mlhgNSGUDDrKPEBNM3/JEPxxhE3Li/X3VJEympOgghBEmyGN9BEoU
D0FDSLyMO0bVIW6lpLgAimUmFnxDVNYMxmqx6XmmfMnmq/t8LhQBvyiYXLjtphSFBIY1Au9KF9j0
9gEQdXsYvjgkiSeAwHk8yq/Kq06+hnsAEH4yOT4uwuaQ4MUCDWfvX93NptlCCBCafh79gh/TvTUc
akhtz9wIxK/u5ZffoWXX/+yk2/e2vQ+mlIs0XomiyOumtoqybftAucLE4BjUK/VdkZl45mYuou6T
W7Nk3YTWVRU16mDmFTcg6F9zgY6Qa8XUrT0ODjvAxuPOzvTQeT9AesIpqBuV1f7UjrAgTkCjqz/y
8VXHSZ7txoSGH8pr7CC0AK9NnGT31G7NCLD17JkeaP+9cgbksACFSVSbAUGUTfYFkMe+/ZwilgHE
12WZIxq+fGt4ZwVMM3M2rXLZIL2PaZywrGMu2FsYOMwLbl68k3ug6j0WRmOVmY4+hJO+uihAyGQ+
3y0lK4+qJuYWAwO1rUchRPOO4MY4E/FnIotdOcSl+EUEOm4d1lusOwva1NhUUQZpZF8U5AIOa881
ZjoCdPDnWsx+hpEclHAD7Vu1T0csBRmd20hjBl5DCn9MDVzfCBo/0ms7Qi/RMYeERMktMJPdBWky
Il07bj7s0vmY9QstBwRJu+CvFElaXlxr4AId/toSTgq8uemlsG2esbu6QvWl45wXJbaKQw5lCRFa
Wdx394rpeX6aMw3MOELisjX7H6i3LyS3/NFkZrb0inZIYRDsA/74etYp4Lw3K3kXkJTPrDcw0/IT
glyLaMrPpk9eEJtJZs+ZB6qpEe6EuOH/d9/ACYUyHZUiMEt0ja7payKqoROjtk+qI2YEBOjaH8tB
cqu3rDsFP7u0NA+nkiU3MQhiP04p/iSIXHDoQorb1k3AOkiWRYliQz41lClw8Jfl9DfsuUJ3CFUY
t7Ia1Jv3GXd4L7HKjOoK1PQwZO8DsrYF1Uab0n9RqWHRnFKCUkBJ5aCXsUDK6y1Z0fOGx3GbHoD5
3FnYe5D7vemXCizuQbdcPB+nxIkXrFxTedyH8t2OX2gp1vGdBuDADiUR3ReFvyu++VrK/z2U1ZZA
lZ4M58rCmY4PSuEz+RgE16ML+6nK6nT1WKg8iOq+e9RAlRytKRUJO5U+bbtPkYMuhCEI3LaNN0Fz
kk6Y2ztGO/ctgJ9LlPiAQlLXbi0zIP3ldzwXgOLwZro1KUprTzYDxQDN04zIkaxb2raTlAUTKULd
wBcMxTaHxjUVASFWZ24O9ENec30viHbTOf43WcrJVfX5I5N9RnnYxdkfgu8npCU/tmHShi+2xheF
L3u7yD9iYyF1raw3nzipoopxm2YD7djelNGMLbWqsQKeac+nOiB6SKimNRlxJi3bqoltI1+AiN7A
8gvoTdBuv/4g3wsSWKOArs9WT/tyFC55EDQWqxuqXDtHoOInCFQL2Ksy6MsZiXuUUAGGMr9WBAje
sI2+1/IOdokdYcDl6AllCyE6r+Gb98L2ZXr9z6XHM0+bSCfs8hrUtBnmpntIVp3xXaNVJPVF+nKw
VNVS3ZzLh7wYNHOjN4adegyVYXXQjAUPNQbpjhsddy6W/vSThY4qQxzE6aDjBCHX4WezvD0fIqsJ
iUbWWY/b6OMKk29zIJ/mKHoxdBXSLB903m9nzPtib5wC0zaRrVl2YnpAWZUamo+HD90gUsbHxnPT
E11FlRLp7rgsmXy2MpMR/uEyJVlNlKlT8Caiec3PVQcsfH/b8DAw8F7ciZk5nMfLA10em/ofun1N
PqcSI64lt7OnzXhYYo62bB/VhJk/lHOtBO6tIIcY4sBq7bMDcPGEKqSWguLPRShg04hFFYAWbXGr
8MzQXgoeFPDeFzYgOzmqhdWFIU27/66zOTu8kYffnO9/4VEUkACuxBMSrP3MZdzBtB8bpkTXRXz6
nQE/uGyQ9fRTfoYjPuyXVkAogTJLTtJCu9sMaPp/bf1FqYPVpK0GIvQNzByNDlVks0hl37EMMoG7
PO5lcyKJxrtFyv3ESp/YSUh/HXTXn/h4ttAz3vb4hzORAbkjKjGZ6sv4g+rnJB9i8z1oJ+suI00L
399or+c2SUYd/Wo51ZjkG6/Xg/D3tfHRk8lvRrnPA+bBSjbKZKEAi6yUyYaghN/BOKkFGXNjlWxv
YNWQkb6utsgtFJrtRKtEyLzTVQchU2OxwzuOywP2/hflQ35KuhDOqzOkSv/PZ2D6mFNISawd0Xch
Ov7w2LcA4GwWVjWrb/2fiMlwZc+pjVcj5HMIUXgeHtxiw+ZGxMzORn3MS9rwDWgTWyXznyaCZ50O
BcfCzRqLQSFHEi4gkl7pASnFWFykaueCNGe9AkdU1dFzK4TKPY4aCyJDs6/KRGyravFUv598F4KT
Yp5KUHe1+jNGgtl+SzsgFWNPXCw49OGeIZepbkEKuGTHT/jj151lgc7whAjqH2DV/KECX4XlKDHs
rVoYVDC1i0WWAz8DwuXz+a/1qvGnWO8541JUwxmrDtmZzF3YSWOqDPfEd/ezZUNdOmkFct6jlTq8
cPWMMHjfKYSGwgYvkZsXwz8KLrQ5TI8GjSW/09VDj4i2Jh4HWzOlGmmcfuq2TROVkIUB4W4FcqiB
VscT0pEeepr18x1y8Hsnx+lUvRXygMAvfrV8tWhxyPNNEiCRE6AhgHIqHclAFhMOn91OVmmYrv1O
cYRHTHv5fSbUIQ92XVqBwn92/M0cwlxIxWRbiPmwfLRCZhKP5on/ugu4PfUITtjAxtQcXqBG8UfX
6SeXYi2w+keBaKqrpSXVxhlJYqh7Gh6rEeFBDJqO25t+K21ZIjRZde1nkLdQMGn8wZPzcV/2ceHz
KEXf8kZAKQjDD3cIU5bg4H9vJqW5q4Cgd6WxYUKPXVJ15NtD/Ze4/0vbxERcQfanJxQEk72mDgDp
q47os5lQbnbwsQ8g5sN5MnevW+svRBuTFxi+zUG/3sRPKLGZTDAYR6dwmr48PsCLh4Gkq+XJeQUK
83QiYDA4iNjFdrB1C65zIX9nDU7Fmh+nC55XJpAN90EYXRLWrlyDlxPHOQSkq1Li6ObMlmquNIOC
u1BRmgbc8uQaYg0eyezi6odvW6uUvbNkQZbxSnUwVbFofl9eleil7L2S6CPFkodSwEkHZFXhjITF
72jwQkC/9AbocpK9ihbnZpC/1N4qaXuQT1r7XM21z9V2y5APKqM6l0HmmOLpA6KzTtJ5Si92Su/Q
jPKdvpV/7FkxpCGL6rmky18jLGiXoc3GTVj/4yLLA/gN9tRXju0Y0Pe4rFwDBs8pBD3f0oyuDXcr
1bdneGti6S1pDffmmHx6lCzbQEXpukFFjODZrBwMvX7cXeKYY9L7/qUB65qRpYt6OxnT8IMbPKI8
w5dGFgsTXGWn3KTTu5W3c2wVCRdxheGin+OOEoln+R4/tHGBI7qtJklZk18b0CqZGjp+y6dhudY7
X07J3uCmUcIS4a8CHrPXNYg1kBEJvT6wyx3RvHulPEFcs3sB4UyOTjQKwM+MZ48eIDT985SVYcp8
mUQIB8t1KfJM7UF8RmV3WJI5Xc8W+FxvXUvd2Uoaruxdr34OMeNLJPJNHzC/799SkGCtcuLudqBL
G7kdWPg0uwyB33LtVzvtJanm9ACAi95qnnu3cgiqScllKE+mqT9H+Nli7XfbG2na+2Qn0kccgHtI
21ZfNLm58bOz1XxjB4P12cb2L18B7c505gKH0dT0CuvfjvTBC78Z3awOebOVY1yGh6jRBZMc1A5o
r4HpQp6O7Su70MoBmVLfevYhK9XdGoq/WnzJzgUhOGpLAYoKe5s+vvnrwgX0Q8akhlWkFyGr5+53
nS9wtLGNjM5HfYzZQnWACli0l9HVGStnk6P3ehSZhI3Wg+xw+fAjEhFJvqiVy4mnvh4Pt3F9Q36U
+mMVDX8kv/zCTEFE23JbBIJrv3q1+bgy9FtyaN1LKMNWcsRyY2INFlRULIsQHl4xtvQJdGHvXG+r
Xri+PBaQF6KgMAhaz1AcN4EhG4qnvLpHEU88ybDakUBvkaComY3h0cLT4TbrF2OkuAYci8W/2pTp
N1pOFbgYlkdCIfM8Fov7sAx6dnfb00NICcBBgxTS/9dH0LQOKPQmrUWAm+iZFiVU7tVVK1GsciXc
nPc+nto1ndFi9qF3tkXvG/cFGnMpf2Hhft7oA3k09CS1EkpWmhKLj90kZLQ7fcxlxndrmMcs8ONt
gRI+rUnK3jMjAs4SYu3H8o1nU+WV4ujLntyF9ljXGDpmhAj/zq7fMkQgKSzfx1328uhABcn0cEyV
mY6tsxn05gF43lJoZ05ehl/aGrMgPZaengpaU078JLTNrRe/pl0LnOE+XbSoiUCwC1GvmCUsscWv
/JuFj3JGRofjEhwAZ1ZRzJttFnXbZ+XrL649CfNWDj4kQnVrcvDx04+vk6rCiEBI1Z9ZENrecfnX
C0+rQJwy52bw1QBB5sVsCZ9u631i8NEBzdfrhv3W90oOGhbs/E9//paFPH2CiyON9lITuFMw6l+M
lfRgPv/ISW3ROrVF8oTk/1f348N4Ev6QxYc+hyCexBQJQXjgPAXqPH0nF9O/j7f5a8GQ3mT059Y8
CWAoDUIuFdezPbtApLTWuObN4f/oAWrZcU60IztZR0beHt2999kXZ/ET12VsIC5nXvU/KkREc3LD
I03B1xUVHXkP5DXgmgByJT6nDdU3ih4FohtyxDLOEaMTJ99AYVA7qhWgMBBjT6ZdBeFtJ5McUoiI
WE3nQecFhSdVVVr4cMzYYAfPdr239DkcoQw3Dn3DiXjXvo/OsUkMp6nOGi8g4ap8VXwrp38k3m8t
7rfkpPrj1zu8F6U2PlyMNvc2cOtThBu+k58/UE5vxhtNzmmTFM9T0Eq1fNq4Xsxtp/j0QaNkWhwi
5X1uHbTp9CuGOJ+w18pgrZ7JvQZA4G2lWaQDeUgIUBinip8SkjOEkOg5snON5r9dsYjRJF7iIgXb
rKj9Q8EmUlWPvfnnU+QZ2lcS8v9nOaQjqFMheUbs0TYvy/vAogC+g8p6G3IuUqRNh8GRRUIdQj7w
ul+vgm5J7wS/LIUPRmT3ybKz1ombvILWaMGdxqbQajuwiiiJEyjLzj1nJRX7D0Y97gkBa6t3OV/U
dq9PMx3LywjdI6qqowKzWBrELRdQiviYL3NgCjISs9dqGqIeE1bTA5GgEcaZcGOJnl8/z0NQjbdN
21JCRPEqyf60T9aPch1gF61fd4THqRRf0vJGu15BRVg2SfJ99HgprWigUJjMwjO9CxhZle00Pmwn
xVK/OLwVCxDLcQRP8KabnxQ4yyFeYHEbd4HUcWSKQPLmAZMMwehboH1Kx7MqRbzLnZplpCZXuHrv
K+Hq17LXYX0pVBTqSF4mJd8mF1pdIhPiLqXYfP0YKbxt+DUtdZSx3tYUIS+Gpco3PcLGtuPSa+Jw
sJV27eDYsNlSJQ5CceBW0Bp/qkVb+v/XnVVlElq706CJUE9xmCi0tId6E1BG0iBMKUGVMBKcVKCn
VhnPkDLJ1Axn9yzHgfqWBu1fGrZB0qLvr17HCUYzM1Maou9mNqYXFmmRLfvHUmxWpOV/UAR/bnHN
YP8P+orpWJd5PIoIxWq11qgm3qXNJy67Ahv5BaN4eGFMeQu3AMguuPHsTJqTbpYqpPkXkmLG/O4f
erclvrLbsRNJa+kccIUCKJlIkQlo3UY0PZbsCXdy/0jyeL7fxVEoM8+vFPx0BLWs0fuDw8WGJuQN
o5rChynK3CuX+DQ97lK6CEzCuLGibksbfnXL5CrXtxGrXUbe/LoIS5tWvz10GUoMvI/BFP4sXivT
3o1gukiSbMGHv06nfabcaq4REQ2IaiqG8H401V9EAOCJaeccfXAvl/RylZLvO2Mgy9AtH4zgY8/p
rMUZstBWgUUsi6QAM9/u04MM6CtbMzOffo3EPJFUCFP0WrVcvXAAdDWm6nduqHO7bxqZjM0ZVxCq
34RRHPsbGe+k/diO+RFLhj2Zpv3cLAJB5imohez5Wt512j6Rghp9QR1fWPkbhnP/2wAqmlZdK3hF
K4YW+mEOO/BoO8las9KTDTYfKIyS/PuGkBnuu85NJu+PRT+pRXs+2Zfa8vnpvoD6ruPJno68jWQZ
OGoLqLMWPTf5+nQu4kNrLwi4CZJ/zlplmxBGX+ptF7NzcE7evspKNPTVPBoxlgPKCy2EdLzxGABN
mIP2dZ0F+Wa2HasQeXfLn7AIOx+FFPxZxrCGXHHyKUMd7gNjxSUnO4SaCehsWJKvm96PHRxbu2Qt
zMLLNDd1VvlGnFUqBRPIepenb0NygKqPvLFAY+Z0mN3CXlJ8SQEyxyyFBVFwIFNS/npcsPPjh8/d
Ep/ePmCEPJ3vTZ5hUCUDBU/O7Wc5zmPKzvqV49UgoA+SyaWB+nYui1ING4HoIX1AYmUOQklKPrqj
tiavM91LwY0laIvSDbXaaLg/RmBoGc988n6VgH/w5WSEymDC1YPmqX5jCsi0myCEwPcyGi8Aph/6
L9Tm1+tcC3Z9qI10FyYSHzVeL3Yo7WjqGooqsNz6xMZaMkuAXa9VOkM3cZShFOzB56vO/1VPVZrt
n6USIcaBf1p1fB1z4a/ZoC2jtqTkq6+8ShSqi1spF/5bMQ1Np3GQgGF74BtG8deBA7+WlZbx/qIw
83TdPUy/MrtrRg2+RCpF5HJG17nlABjoy4HObBQyeP7yFh4geH5aLGl/SUuK7Yo0WhNjhSk1aJlR
y18pRHYBc6R/MYBnceOEwyEEQTVbk4+8X8jMQUbcX/6BWySH05a21HEPWZuPEm/oPk9fxynPWiPF
gNum9fu52HzAip++WD5KF68TZGp1GcfT0gKFoElKDkjg++iCXyIwhSXtrhUmhe0pdRchfTMkaMsK
0Q8pNwvLX3BiFvBmvdyizvJw8YuEh90O1WzqbUEo8OGChSBhD8wwAWAdZjd7yphyfq4HFA+zCL/K
dUXvmhKWfS4vHqCt7P1tJS8cZrRDXwtlPEpigdq92QoAo8NnRr1RXcpucnQ8TpxvFlRQvt60x2Ic
Zu6BL32WWoWPA17ToiibvRiiTo1ga5Iblbx10B3ZXhnNAz2zRzajT8LHht+2EIusMAzCy3T6PIi0
uCjvCCXV70Y1k/66DHW7ymi52knH0PUidC4UFAKd0YIucfm2VdBfAgjt+XY+zFJedI1VS8WkWkTM
cDlEYlcsP3QcQzP6Ylx8dFLiNmiZEV4gSyU+wVYDNHVSWFBf86bEvnNntVQ7dILinPZSI6DbT/4C
pfOhqjcKw4SK0zohR4fQ+rYRqYu2IXwgcRJ0eONjz6bT710eUvREyAvelMQisi353FIWZsQ/9Vqm
R44JdBeAVYECKHcAHPnfSM1OqHi7zQmUvhthPOZbT61HOOuUYNuGcA3V57wYVAcDdmdrnTfP5KA7
9lVJ2qX9Wj50mzFtxUk1GGsGnvNimwog06a1o3d2OoeVc1UYeYo7Ce+qt2Hkfapvrkl4GkwkRgGq
EBa8Gn+2ZEMfJEO4S2NTMdAJJyct9b+Fd5DY3QEYO/iuo4NLcrClQzqLP2BcbnPj295Ou9T1eCkQ
Atq9g8mrLiRzkeUkxelt1a99KAy5k14fejZnVN0lTcR3Vrh/BUanITCips5vBT2hm+umhxfliaQ3
Q68IU9CBPuHOdfYe18wap5G5WPXczB0N9narJNoSK5pff02IjbAxCMU7u4bsX3nids7ztKXEG1f0
djsZjNY63tNia4BvlDfzL8Xj1Ecv4Ai66QcB6iV3PY/NuTHer3wQdLxT3BDNdEOzXb0akPFWLX1Q
i8xRyQb2q1ldhs9iwFFH8gr0V7iAAMWNmU8VKEItRcRsSltCu1LF2YJFrZZQMt0vBsswnSh6Rbtg
tAmyPKt3uFu36cW+lzyXUQKLGoUTWjmiRXzg/qp6RmUX+qIayWy+RfRjJ3kchWX3yRut9SqVrr1p
0k2pESwFQCs2pEz6QUPs3I8ZnPZskf2A1SqpDYDSLuhwY+OPW/nzFFvFOBGKwBBfRO5n18FbQoMN
AGPCmomKPqAi6IHEBsVjj6TGF/uAHCqzAHzYEYsJyfXhzTqNqBCSdsZDJy0Regu9ONeg6+DZcIgz
AlI6IltvzB8MfeQFLOSGexpwME/5DxJk+Fl0kOP8QZdiyFkNqPLzOMKvOf3KEp5gl3380K0U9HJC
C1gJ4qf68cVXXWDWuQkcxb1Kxwn8rIA0HC3I7pfeiXQSaOO71yF41Lrf2Ucx9C9Uv4uunD3wFAL5
EsF9b5eEXVaSFMDlbMFQNfUbNeO7H+USlYy3o2dymPVfzLyM47Hj9nMlFrwpw/XN35fS1P50Ce4d
hX/TUrjnE8WrYY+mRlYzfI64KSiHYAykSNwM/i5MzxSnhixJ7BljUXcBnyCV3eaKu4dzdJWCMNJM
hdYVHNF3s21VQrWmqLDqPo8EujPqcz5zSzh1EvvxM8Evrk9KOQcwf/18vycJGalZTbaooel14Exe
0zvXQ0YTL7JpGpSMVuBKaO8epe8h27wcTYv4fy5NR/TOIpiRoIgXQekqL+mrQKyX4T8rPhkBbHC+
KvRQ0clkpE/z9vf1qvtVnlwLvQEpyIzDuLMO5XNDfUdthhNim6cnEZu61440n5VytvBhstK/CxmD
PJXe6pkSbg8QPAIGgSuUsu/z/ZEpidtFNTbqelqIw9FFWzKKQmqbS9LhiXmaCx9y/Hvuzy5gTtnt
VoY26W7ot2pRpY5Ula7Z6ytgDTwbG6lZZXeMEvp1EihsJyw3qWTSDFyakycgQa1122r/rOiartIv
gKHnT6NwARj/Z3p/53jdSn2mnChbixK3WC5vL0dKm3umpuVIqcpFWS10SPtF/sF8i/QiA7/Qnhoa
yeo4mayI5EEW7+wA0TIoI6I0AfUbJP4e9jomo9vCNORloXhQCI9D2n2e2sjNWUdQBOknuQ5hBPLP
FYDS1S9uiC4WyfvSxi7D4JW10I7hdOLFl955nBgyNUjht5YgYQTXRYurOzlJlMDBO/6zrCknAls6
0nVvcVxYT7KF93Op8uaM+HnsgdCC9jdko2TqTBGuA5zZt+JnmUI43Y790EIkR8reLyN1fsd9lRTK
//1riWEAwF3ajHZ0t4A47/+f6MbuXbZa5Bke7NLxulwY8YdUen2pGxQezrbykpOFDydUJb7azA3q
BGO4lH/64aN7faoB5twhHHKHEHuxSRqTfd+6NnxSt14MTxSMFpPN2xRq1esL+GPq4WMUSdqqjwV+
CtoJ4jQJmJu9oXt/L6P0uS/+NrgtM/H2xQGouJvCXvL6szJRgXBRGA7vg/+t0ecuRL/+Yucc9UvR
E8+mBFc7TIZmn83LuqlU5/XL+5/1EJeJGLV2opco6s9ngAm4aHHy0dXqAjcuvwk49ADnkI0lezso
RjHq9XMo+pFzIBrSLlGE+tWwE5HLomlx/jtx9hV0L2cSLpxYCAZ3erxzQCF1kcLluTpsxUvHbzid
eWB4UTNnMBfDsiCv+ocZoFb4Trpo/oDEfzsfOm6GabgA23zg8g82LrbcEIQ6xIK0vRa2q7+/8WNB
ew+AAXyF1UsxN2jOCQOF25aHhwwmkpUt23zSMgZSLO9S2P/K4g6suy5e9KTiF2gnX52k0SWWk7aC
FBFpfSrqSwcf/wGWk0d5NGw++gXJtKrOUzjafzi3A/VVsgrSTnAgpi8GvuidpqSBgo0n0hy7tpP/
I7vNInaPpuXaj6tSOjlpbLRnCyBzsaAXDc5qNuqWTfBKvG5mrtm1PVeam5MZiRJBzoUt3XRskA7S
p/7l2ZRT9PM8C7yD+gx1UgnKowPZlGTDMexzxCaWGugf4Nh8Yi1AVro1E13rgjXcwZbL7BKmuN/V
WBHUjEo7uatbZ12pCYMXGdQtKOMHWYOyspJuRdsVQlCt+Py8OZs6H5YkEE5tXCHXaKsXadQF2JB7
w4TyThF7BeP/9NbZTwXTkvmgd5P+ODmUqpReDnwr/dWFO9Z8pV9i20wqUNZXLN+57zJIUlw0892z
5F4eJ7nAfPzdpfyMbI22OMNAyb5YoTTT12eQB8xCMvcSMmXjrSJUSt+MtpUt5S+02LzosuQID3lH
kcr/BSiRqpbl4KNLK127CFbA0yvyAhQGT3TqIU0SQqzeZ6l5WRcjI8/eZ0Qer4j53442HC4lFCM0
uDJMPGYEVpT+WJOS1v53bTZcopSq9t/9S2w5CtX+YVJq8eaGmNoFFdwCKKZFJiyuXAtlcxEgX9x+
f8wM4swLwtCx6/xcMajqUU6qYbwo/r9DAyIKcfF8E2mYe6qQmBbvcOAz+1rXQD6g8lwWi/Vqv32V
o+VSndIXcKVtwwmYqxVk6tUjMWPjHS7jnk65mDkBnDDgk6nznov8Bijl0tUeT4oeJo0ARis5tv4W
hqpDvg7HN3EmoJkaMJ+Teat+jE/bo6ZvVcryeVORquR+0PvEkf6svzZKLpbLma1zM7jeI5092RAb
hWQoTo3y5bMMbTUnoHGGfa/EQRBbB4eruUf1ddmZP7gAPlCSHTbQlXIiW1b+Wns+dxYbZoQze22p
20KD3t/8i8oea0ZIFCRSPe5+KJbrcoFTD9kRjEqd29Zo4qdRXDElFU0rfsC+O0DaUTI+VmLDHx4O
cfeHbcN9i8o0QAIWiCYmR2sRkTT9XmHIEAHuSNPC45lZoTXqpdyD+bxhRsxxjokaFg4KJGTCceDl
G8G5TDw3oJDGGcYv3gH5ogzEScR/gglTaqnkvZIJ5m1GjIEw85EHitPjD7AbhhvcliKjW1WpAIym
l2sm0yEPFETYnXjLu9Img+X8wyo7ccuA2ftMyxsYt6LBTsfjxdDgqGmpzePsidsM5Q2iJdRi9m99
eEvGNuPkv0cq2ierEhX0hQKD/smVFzlIs8JgZc0KC/odVSTd0NZas7tTMW5ymch9/K4F60DAqiPP
Pit4cUfDoXqlOq8vCneuZEvyA24B4TH+mVgT26KVA8bkV6OkcCr0sWXSMzhYXyD44HY3068KmjQj
ubd7lelz5ZUlhCUUbAApknaVWWqGZHiiAL+TKK1AUeNVjZKm8A06aRiAx+JpQADBa4mKe5mh14Vh
UP1bD+vL0wcXcKav9I9VqK7aUts3REvo1NOIAnotjWkxwhMUqx9izrhHMXqe+ku6FpZcUHXPs8Y3
6Q9jtWgzVNTcsNcAvO1mrKr9TjNw9x0IZqHE0H0bs/zx73lxwQ/Ff4mYgeQ6OYbIWcI8YgQ8VpHD
BFaq0S+qNrTGdkq9AV5n/GN56pzHPw5mXd53WGXAwBaq/5cUG7p3SfnzquTpVgysTu6xZQCbgYPE
XDxWpvWl8lC032Nuxw0BAWZ8vNGXIcHOCz1iavo67caKpg9UTyCT0RWS+Vz+OtAXgvZcI4PHKTyU
teD5Cl/XpO/GUnyZbTR4/NWNkHQRsuVL2qEvbaab0OQgddtAPWuj07LFHyd9BLvFobqC7r6bFV7t
ngmFd/0Zf8cD5uAiGgYE6rvnPhS53nQt+pGqDy37yZyw9bEW7kgyhP23dwBiWPa9ykReLbrdw0JW
mKxhvbsCfL+ByKiX1xR6+2TkIWivxNgv8iGis6blp/O5hwl/PxrYHGQfTBKO05be2IT49Rqeo4UT
hx0L+4kjQx1AJkDMeDeZP7NdLcCLQYKiL1q2K3NybrEQvD6Wzd7tF35uYHl5iWEpPqakhoijf93A
qO1mbkAwYe35q7+VKuTqaGaWTZqGiiODidrPQzXHUQEySN78eEyGHWGhO0KbC7z1F3la7Odw8ozv
Lb4CxsgSKDpJlBpETP+ske6FaJ1rGP6pRP4myaYPRMRxgPXYLmG+vKRyM8YT7GntmH6TqoduIVlG
vK40jYL+Ug5mvzjk5PNBSIfD0KnFOijfg8R4VcnHJlxPxlp52CJma28hC+ctFDN/ja1ilQc8c5mS
zITP7Wlsz4xhnSFrAnTjwWtpHSI8vJNxRD+GAeGrSEmiBSEbyMZG4cfV7b0qxK6CC6NSfuqRvS0G
BDHqcls6bRzJBE0Z32BqDDawXnxuOjWR/EQaGGXclsoBjL4hBYvd6blpAGfjwK2L/rtvlt0jVRsK
TCofzCb+Js8YA/hsKmPkLzK/rhnrVt4Q4hwHvg3vvpfSN9LCLBI7um3Aw+g6UcT2arY7CLhYpPz7
HuPdMcRFpbbCEhVjR30GupJECLe/GQheDRgLuq9AdHXvX7W1/R5PbrCl7RomcGK1o/vAprfvbw7m
byfLSKdKThbeZbP8x73PpPhib1p8IaS8vURNrV/8d+1fFqo6iWM2cLB4iw2DPHTirDuhv94CoaSx
1nQ5Bc1ItJkaingRWUEpgMn99pJuDWDaqaaMVOfiWfOMHIJeuJP0lCLIyKNH8XX0VbONrnXc9KvK
ae25XgxQwZzSiTQEcPffJLs9VE/ZpApfgUfIOJEp/SFdIMn2jDuzTK/oYHXcwfyQUL/5KwfEuHVp
jMDwahFnIDX85BB+IZ0qq06jxrfZDPFWERd/a2RSMpFLwegzvLRKQ5mi3LQk0cyQVWln+4tHznvI
zQDqLVnWesN3XkgiEfyb2qQEdmJx2Lfxe1+fMZUlZ3cDMQFdxfPZMPjfKz2fo84Jqxrw+zpKKIUE
E1c6njmt4LzhQpjBSJw285l0qnGV4O7ABEuJeBdgu6hws7TjQNMtX7Pd1jFWeCsxH5tnfjp1ciwE
A9dv+PsrTJCJVCvzX9M7VH2EHVFdXk/Z/qSizo9oCthQ2eHPwFVs0NmitzxNLtfB9mpky9GPlxFD
2TPgLzGXWhhhFLecS+NB3t/+8t87FgAvIcrU9sTJNSMmmsBYKGo9CYn0zLAq26HybZc/YLDTH+lI
+2syayQW+yY4oHwZ7kYnSfE0IUvyk81Yv0zZLyl4x3eDtqoLr4RAwAd9E8uwG+L4b3G0doxRk2lo
2/CDHBBlyjxJv+wI1bFg1bhoaQAyY8DhNLU1Bc0OFYW9z8JLIJ4LEgiBsixJIrvPUDhlg7Cjusb0
3WfcNBGEe0LCqjRPNKEnoraTjXKJU9ndk2d9OSUcD0XMNMPHUPIWSuQG11X02M/pZOIB2njfT6x0
9U2kdfNni3OGsfX0Lefgew8A3MRbVZTkyOFpyW+J8TULzQHzVi4rCfDBhs69gy3JlZIOkxiOoj55
BIJw7oQwLCnmSRpeCkhYx0cpCSOD6a2QD28KZNdAO6f15zUMgS3Iq99Wpr1zXZyfUdDHCOwGTqTH
GnNskHbNX0aeBC/DVLieJ1Oq8ZzKNF7pGkp2FtvS2mqbLkSvhieGWaEVyIeEwAsywRzpJro3+PVt
qoYLneKSgfIe/c1pbNWPEqj9OJx3ICjwLmNcvSEsw9XECSjQDrtE1OGkjiPmPFx62ezkW691De6k
xPLBVpIh+kUjuLVL9wlPdmwB/BkeZgO6b7it47iu/NUSapeQSB2XrFWmTgxK2+NqI06ow+ZDKnMJ
ZNvySTjr21Oyh2Ptchg1JuQbVdjAzRA3N9eDxBOQFJeC5H84WfY6KYxFrRu4uNUDmoyu9yY6Qtkh
mZq0il0eD6FxkKFtv8WUUhUsaGkmN67J8jatWRJBxH58Si2M6MvKj8fUH7rsGOJ0/dP9hkzIeXRr
8BEVlZEywSe6LarTOpuG9CbRtggRkwNu+xzlb6hUIsRdfXB3t+stYcwwXJaklPAkQtQ4yH8X2ums
PyQpNMxKoFBSTzyVzI5+vZ5df0lwd9g3fgtHzolhkJ2zkjS4NqtvTqfKbIhYjR8clKorRzvKnPC/
YPdMlIr8GdfewV8sIBEcg9HFZKxUWkG0KB/pR87EFeqgeZgYQp0W11099JgwZKlnTtdGqEbtVWrW
RHgvWIIySe4KL2TlPZVDUA9W5mKH683iOj+y2uzycdMoDq4J/IOt2GKPN1Fli3JmH07xO8GtxlAI
qHWBDkvDCOjPukZW9RBUlbHJ1r55aQuqYJMqTWE7bF0unydyzi1NLyOgkGubN3BjOF5cVwLX4Eu8
XRRHtmyedtSJyl9NU/K98crarcuE5mHyE2QDQGU7IcxRd1HV/IkgDxQ8dqmSWl5EKMP4PA3s4mKI
MWZvR4tl0J7doNXKoTIqFgJwqWnNx07pcD1Itm+1Rj02nOH3BAdR6LBHndrOG3QajMc7OWWCMCxc
OyIEuCz5U3qFSX/kNqL4+PI3etiCPP6wAFuetrF+ONy+6udkvIReZ7BWYtWF+omjfFxUEmFM297l
6mEgbRBzCVuyGvSo7dQ2wvBiCC6GwMdHnKrIDTiBv2Kmh+lJ0VpzUGgXQF/uP3zwgpN9j1Y9X++T
i47HUijaAz0hOk6wpIPOi4nQJOg0YphlFd4t5fko9hcaT+U0SBMwVXi9AlP9NKQRoAMaEIl5wehJ
BN8dl7sumcxZbrGd0pFT5R4h0tC1rIU2b4Eb3S1M8PxkcTMEZ8xHleObiv4Xeb6e6MjTnIwuspYs
kirLKdotdjQqLxVAWri2pSO8OXm5atWUoCQZWPRoZ+3TnkExkUcqLtcfII161t8j/w/ayB2L0bYB
nkW/ZYmbUg4PoOSfoWP45QJ9H4Rxp3kky4DVQkrLZ3s0swmNY+LW+ugalEsDG8p3kQIzUD8e2OJ/
JmJONxD7K8qdyhOFCwH1iM7HDdPnH9L5h32pGGVMaxj3GY/JLXqm0dpLUC5nIkt/IAfmNl7nFY8t
tMmtqzV1VIu2eO5M+lvC/N5Pon0ey9ADnVOsQ3GGY/1c+MR8tKg0tvE24SXjXoNQVKMDYUADvERo
C9OtSZHFcGqBBbWqKQ09359PEG+b+9JTn53H3RlkcJqYetL6Nv/YkOMmXj3BKro1vXiT8iIa0oY0
eGU4ye1q5JkcWPA9pOg/NA2gvPSm+UgxsTW2/D93h8SfA8yffn8ZglCoAZHHQa84L/Z6wd0FkmYZ
MlLR7yxDuBBVEqbPHM5s3gzbptXDsl4o2NY12P1+fOVUL62WtgwT2XC1+tPDIV3UBQzSA/vYNSDU
EYfUarGHxsUjRzlAE6BggCuOh7R/DE01LRT+iejuwt0KelgR4+4Luvfb5Gow359a8tMQmu26IokK
ukuXPEiYfOsriSKco7iAwBPnrgBSkKG+Gfuf942fJwrIAqg5W6bx1Cjo6yxeY3yBLbZANZD+Uo/y
GXNig/jL+pW0Hmx7H0HDVNXLPk/E9Kp85P1FN7cCA+I60Ue9T2UiWxg6iAJIOhooBytBPgRWmrl3
wrBGPWQLdbDE4fo+JK79mFP8ZdPyru7EB6eNNl6URUr0JmqSozj0c3BJGE2Cu2e4t48Z94C84+ae
ogKS/yyj2IuSPxNGGXBKoB6187AKBfeJAcsXO/bldViDMukvivrS4iyFILMfb8Hh5wtR/IF1wXmL
/rxjGbm5zaWO4mPl1PsFvhT5aaK0F+mFMQkRYm6z44e6ejmfi0QBpI4+SG9GHVoPt2Y52mMuUbAg
NVbZ8M4Uow5AV/L9bONbL9rmSrEUbQwEnsipW7bOWaZGI9I1CwJwuw3Ji9WnZRzZyzd+jdMGOKKi
0w2zGktY0og9RxzA3JdQ3hKoC7AK6IIQSNni2rJl61I9PDppVfLYxOCuEef+xQKPmSIeVn9ob7jD
dgTcqSVt8oXwCr9epWNTwqQAWnnOpt+ETZfavsbaKsipu7br3doB5EP6gD3wHY8aHdQKomE16yTO
QUegnGogTDLBzDqoolX7Nreu/gMDUf52ZYVnL1W7ykTKHsOR0lJfLdrzysGcaA7sGLxlB4LE42js
V74rWQgM3AdLzdFgts9jurRwuPPS//fKnV4rvFIpzJhn3/MvO66V1cK3xVjjZFXLs5u68pFD1kix
XdJTR2HVQlgEvfHdB6TItivsTU/Jvf5w2Hfgmb9VnB7iT/9DUbowTMZgZ3Vjm+/IPkdfUalBF6XW
BiPG8YmYx9EwPztmbXzJek7F8Fe4Pf9i6QBNlcEkDvGyIAy3ZCU5K74G7sMUNlyxq4KoJkwkESOG
JLReHlsPTeKWCNq9kIiZdOL6bHelGNMvk6GV0HTJ4GKEhID7MCkoEQ1CacKuTdQ4zXHW6J2D2j1j
/L56zWCcb5p2XHdHES+D0K4FOIs2ZdHQTlcJRzE1wcQbACVqOUz/3wjR046crYRq4wgBJt8Di35X
sO1qJ2Izai0SsvUuNEILERivHEe4yaHHFUSpKwQlqjP3J3Nkx96NBXh+7YAl9/1Na9wY0GK0GHjP
TmJSj6JknlOMzpnNPmAPij1YWFKPWMV/Lgaj2vmhlbYAWRKbyzXTyJthHES3bcjXz5Q4r65eF/Vo
/miiWwuEld7wQoBEF3FeGWZDqLGWrInumBAxicN0cvf3n2C3fi7NlSWam2ZVTJCFDpzZeorZMesc
qu10Cb2Ky0HRZdAtWUTT5f+dK6pm4yM9o1opbc79ynZn4H8rebIl1PnhrLoJOr10RIxIWvfQEpOr
OeJlitp0mddJfgn4U72r4jNnu+7BKrrgxuo/y55ePFhq/8t6g6ziJCANiZwgfFUHs0JhQBzvidJ4
baOnuwINmpZ/syTay9teCjbZXVdLxlksFP0GIszQOblgflGPj3V3qoFuHW1/l4pdoRKQ7IYir+zf
7ahjaUEs/salhSnFgB7e9253IXlAaJzARDr9YgZl0DGcIBkB3sOMjx6PU8KbAodoY7B3l0Dw0+mD
L5snxkrdFY8G1I/+R3f8is/CuvzK6POFVm5yX06Kctl8zIr/bEvCcwwzvawH9JaeGjGW3tvKvnDh
2HiJPfp4qz+1g5Xztj5POsyMhEbxfbIehMJ76EuEuBeW5xP/xf/qOo49RrBLrsm3ekAfcLNfZedx
uComwz8N3o3QQmf3i+vLAp/LhdXLxmkQTGPbaDr4+OclEw1yWz5Oz5LEcKavkIVQJ2LEIsfJWeZb
ts0F6hPyj1gql5TRoGxKqM/E4SHy3FqDyMn+AMtqJjkzm+zqrB1Y66yLO3t9SHYrPtcbaI6uGDiU
ccWlLcsMboYdItoE/qh+wT2s9hT7PQy21QpPfhRoXmeFJekOuYxt9sxYBk9hj1HvS+8br6mRu7Lq
L6JhE2FPc1qx+8qPu8dcr6HNNkP5vBIW7JxbCJ6T6tJFXwjf2bJyWafewhOxBwyQ6UhIUca2OKHo
DALnmTr4qOEHcKvvQVgsXCKpirRW7GYMuKYn43yfZAQLL81u/numS0Fg7dFVjg27STOTipVy4FXV
8A9dzqymtVdmjL9W9OxPnI3lX4pv8/+EI5E7YK0D2u3IRpL4Z+tmREq2gEkCMq/SucUZAcDAU82w
tTynI8rznojFL1OZJ9REOlG9RLg/TBVwiYfz7kEkmU80lVMEifuZC6kiVgTf6umx/Eo7kzHJlN1w
sAMmWmCRgvrf5mRGToNMYWD2HTSYw6NZVIREZBJ7tUAXblAEIwBq+KvJFH6QFa+h30e4lxjUg5pn
LuN8D0IjXvdXdTMwJTaqvSRratvC4mLJ7G6V47JX2GI1k2URFVo37PhRqXqFopYIZyeubpbncGBL
SmB6zfacn7pJUguXTix3cvBDynq3s/0UtsfaAsq4mxA+/KMfo3wMJjydrnbs9rx5810KKV/f5Dbv
2wUjxyYIhzftnuWhyp3ut05wL6GlHgNsHRMTJ6vCR+YtyFat0NoNUL/Pf+k3EUu8v09HZE9+BYsh
eqYastpJbtCw5dx8mHUQwapjWifTe712gNa0QGyy0zz2L33YjBVrGw8dNlwge6buQ/VdooKBoihX
G7ij3JbC1Qomqg93UOn8uTMl1bFZ1i1q/5DiuXxG1mDar7IDVEzQn2FyVYO3mpwgqgP9wwQl2/zi
NRMyHvsfv+IiF7hkB4Fy2oUAa73gMtAiXCZeZXbrOj+cHJHOMwEdGa5Ch0g8oxJbm0+icjSSED5u
2VpFuBWOhxZ+T8S6KDvnp4CI/+wNkmy+pQkoaEbLT9JzME+LwowilwpZoOhXx4i0DiqNABR6e3Qc
d6nbzgha45vIY6lo8UpkILWtNWqC4ftubE8rW042MPZOJk9MOvokqRsqMbEOsHBBMbF7azDMCxON
YueG3Xtrko5XJCG3EudEURv2EjArjJlFJhp/amDYeE8FfpIruPzcRh8Et9hV6aWytpIN0qBglrlE
vDl4pnP0zWXqbL2ZFTia2AhqNX7aJsSfiwpqavbDSkp4ZQ0/rtog7q8WckkN7u/HzvoQiH0luFZ1
q8swyhfs7AwQo7Ku0xmLoLemt4+3UfeB8r2nHyTVlAyXTcyA4xxpHbNjsH1xxsDzp3vnA7jpmhv7
fHat7b40MxD5phmbv2wzADH9cMvOXGT+1VDP6/2X70VgYFgY1UN+obSAwXvEmgKiHA6g8NfiP4Zx
EIKSROTjkliy2Pin+LEvRlp3O9gJZ50hVmTheajmrypRysHt2oIQdQbS/Qo4eQ60cw14O1Iw2Kd7
nT6Mhg9D56N/A2awPnKOt3Y/8BI/JEZqKCdotAqkLomzHtbf/8aIMcNlwlFShLCTE4jWbWYm6ulR
THfwL0qEeGfBXa5g/AAx5CQOPQ/jzE2ZOk+66JycoxQ3UI1shvfTBOQdZ8Lr8K6Jg+y/Fiw6cGN5
co0djk126zzu4Tzu7mzmk6zwEPkyx8hoymEEWTDDpTW7AzBChTc3ZcTZXHZcbdMQyvkBfBhyWJ5n
Y4RILCXXB4xiFF9RQGljB2db7IO0A5u+fPbTnPsN6JaAFmA6SIQnmG2XvO0YyImyZYKXl5JEzLkk
Qy3aJKQN/noMX42dSe6FkqTeT6IC0uxEWOTJBKhPm2uFoAasVXDKQGJu+awvPA5aEPD740Sj9Hok
0s4fAprfH+gM4EQWl7blmeivtttlROeUAgSEYTR5FGKwZtYY1P/+WVD8Fv0qqIUuj1bsNYZGD06O
b8DnhEoN/d9k4B5hktXU4Z2FDJuN1dLWjBEHuYcBK+vsQyH5RBqDNbS7h4FYBawuZvGZdtpZXj7B
/CnNc3WeqBgh1RPxnIgp3bQgMSmmtEVUUWT2W3+LJ3GK8kj6cWzFOoQHMC6TtPPczbHPvcj8Rrgu
VLI/sQdJGv/YoiTLN1tleUFRp7EpVAKXMW5LwhBdxPZFaAwytzcUMqDRnO4SdGBqutTJu4yVHgGu
9twGNxHJYFO0ZKbxdAskfFBFvgvpecove453PS8NwpZw3kMG/WBLuX3DDxVd3QFjB6LjYAydRpUs
t5WncmouYwmqK9nLdIg1LF86SN7pu64Gn5BAm3kH9VtGL3a1SdoSs82GO3a0LHpgiQkSoAJodHjE
MrnPrVPYJIEoxosRBvDwSG1jMN/fD8kQ4r0S3y+EEwbxAsA2EJi74BHvxNb8qeF+gzdtzSelCNsB
cOsudHc65ezr1/m1wDMSzj4do5tDHDgSMoqTMc+rKzviiUmFIJZGq2xoqe07TJWygjvgwgPXu4wX
dpjrWXG0LrQq9cOr4bmMwLpo7fR/WsjWtd3Glmz2mvUUgxQBjMC82JlzLVLUV6R17LMfCBm6pHRh
6qym8hisu6GFB4pDLwHejJIqTc1bGbMLKnlxsFk1MxhirphR4ywCCZkbA0z7eqa5rsPe6zXM0vEo
c+trSpjnk9K7DZWrvWS73wwjYD41AIxKPMzVG7JRfhxv/qBxjCxJ5vQmK9MHNdPUCl63GYmX7A/f
rWWn/0MeTMnDUgMuhJIHXEqG7E9+XMhLyQkqdkn8i5o1/pVJA8uLQI+n0XzlZGffiWadHlGZYLEy
VBSACkw7LPF6Drt/fKddIxUfalFpl0G2hLb5fRB4TUsyIaNch4FWolTqaprEzCBmudyibCovQjbk
z7hnofER6ErYYdXIP45SRKGib2bU4KeK/O3KsGm9K563h211tap7V9TSH5tjW6OFTFN1t+Sh4VY7
++xx/4Sf5TfoudPMgY/L4QkHos1Q7sHknYuEzH+RR6qao2PuGmB2nOYMeRbJ5HBneK/+/OOz1GfB
kUtCLedwbLC/hSM+ms9qFFKaC556glF2dmLtDP6myjNeKoex16ehWTkuWdiRol0+ORSvpu9/isPM
Dkr3VXZMBghyfHaPiMEKaIGI+3O130jRR/o27cb4O2Gv/FHoIVMrHBz9e14BoEQcje8QAl4zvPNR
PxHguBziib4rX0D+01TBegUl1/QUMTUcyIpWkcixw9gWIosMGLxbYbJXcTLtZKovRxmfpzsqVPrH
eNxESVw/SNd7c/hNmBpCzKxCJmiiG67axzTUnVJEo2MI0Qi0rBnAdGUYeZjLJ9XbAr8/jqi6t3r+
KKV6Jm+G/O+bedX2ik+JuEWDQ3MEKFsE1dPyRnM+HwilZqErLcjC7VlPKPwrs8sp3klbE3vhO9o1
dCraxitEhfJBcPan+trXAi+i3Ey4U/zpdBeWrKh2ZKXlSsqfG/P5snYYqCNucmY8AemuNB6K70eP
KLAyZU9Lx11byc7CGBtE+SnJzEMvK0MmO+GZ89mSLALVOBNlLgHG+y27D6OxrrirQ3zs4jfYQUJV
ZX7Xscrl+2i4s/IJikC/lVEHVT0KUUu7wJXJPkOpql1LG+LFIBypW0jDVx7d0ZghL1J59jwxBv23
6Bdx2Rbm5IIJI4yp4i/WHHgvkpRrVj/V3Oc0fA9AZ7VR3mBYeBuBQt544yaXuooYg0X/f8DI9ofi
49Ra+9mo1GDFmHP3NvEttG20j6vqnYeuTnYKBLZKa2p/IRm8zSE6b63G8CeyZap+Grzv4fRbH4ZL
TmV9P0U1HyqGIZcR9FqoeSk7vXg11xQVRRbAlYwZwO1ascKc/qyH2Bb16WzizUOTyal53Dfvsl83
q8veAxi486BpccwotZ3+1csh3khMmTqmF3bWs145amKpSkmybvjJJPmQPGabhTFuGniTO9+nLFkq
WgWS3bWL3mnzSnVIXDbqgDuwbKoSSUOgonvOVwM+4jo/bICxcS/aIwuq67JyCU6mifmfcu12hu7e
CJmiI5Rn7tc6oCQ4syXdHPeiiuaJocN0annzJBuhuKQdDv4ImzbejoIUTaew9Ki/AJfdytyhMAX/
fJQDAYMONN3RnNzL9f2jS4seU3ZFl2fbQTtdJIZ9tyazcmcBdpuncgagNo0OqqYcovz76JNtDY3t
3bAIZJIkDvWVdJlFE9GURRlC9cJJ99TF+QAAR4ux/QODO2eIxHEZf6+uo3W4wboxEtoQzlquG8ot
yg05+R/fxzETNJuSZyszpza8O+EsBIGoLDg+igSZCElZMCrfT7ZiT4iOK2NmZ1WhCYUf2rZW2k0e
abAl9t4SNKVli/WpwFk2BM/gPriiVK+8aSj/wz6Yx+tM9zTuzPPXunwdBd6iFGKHO07r5JRuPSIs
kZr5theJskzOh3XftlQgLkKXdbAQ0PrqdxbLlm9bj9HaPBLpP0I6yyEEYgOx2QxvFL2ZRIcVDAeI
5eIR+rj2q7bABPbu8DUDIkG4+1UX5riVPeJoLG3NC+mOWvV3ItwI3BSFg8S7iB74m0J1zBGgW25T
mWsI9Y0mWW7CAViSmRGJtCxYFHpKlkJmePpTmlZUZyXryN46LbbSCNzUw1BYkbXGXfurf9WldQQH
6h6CW4tgI2QaBQXbIJg+62/fYjKxJpWVRK44nN7MtDhErLET/ivcoINen8yqqPfwApxYdlnyiYPw
pvYLw1MX8BdX/yiwEJyNl/CNcUBhz/xdarTpxbu2StUEmjPFaieLO0kRtq9DHZmHJ3dTDEet+VFS
IE28uQdecL3okvf18N5wiJntwp0GFLIb3PHOcCzv0vBelOGFMwux+X3Dd5LSTjvCP9L8WGqN4pjv
3h6QmAUZj/wAjDSg4stCXRYle6PWHZqGjjlDaTYrXHB4XZcgok6tJz9YHqBXyEu/+YMr+k2CpAl+
akt0vo7O0YGfFqKvIfFGMEOOoi49IgTTY6Fq540sFFZfOatGj6i4ysN2OXI+9yrKkZ8Axa6jQMCo
R6KyjNfD2LWCTglWgLQFwjeKL2eIVYHB9Sbg41c2iPP4X1tnodbf1uDcUd4pxs2wQO8wnjXay2pr
6orLYwkren332eAcOGiKnlHcxNsDRMfHNd917lN0j59v8HTTB+KFjrJe2646WO/dBRFykyP1gCK+
nv5h4wcJWAqD1z9E/FYt9P10eU4YdFSfwZ/pGZJy8rmJvwbBTdHRgVxtTChudjlaXXwev8Tse6Y8
dev48EnOraWRWvNnQF8uVvOZcQ8Ir9Cxdw40jCDK9rQ6aAJ1CviVhArzE/mZGMwXmFBlQJOXFB43
Vyrkpc1FhzvpKnLT9xvtvnapuRxV3m6EbS7on45IyunaC8H6xPZSMO845KFpc5zz1XOKzKgtLOwN
LK42zdsDQbT6uo9qNMf2nF95Ur5lkEcobQ1xTs4MzMVrfHY34ButRKbHbahg01wefz5uAvvoiKOf
0qgi3YsDbJsH/XCSrd7i6HF/eBc0dehL7TSsXM0cETrIH7eVWR/XcZSCLbHNDKjBBpcNimjou5BW
qAJB47dkkW6l1M5C+wbSmM6H41HCcyiAroa//M7kY5At+MI0zxRi2tGSJuN6VBdoWySJGj6f8GPp
NGLouOBugjmQi29E/U+p9FbC4KHelkqEZ/3KaIWo2UOwZlOXmt5D2LIj9Ff8FcW8ZSXzN5KgSDRL
4NF7k7casYq6uLoZez3w79wS1Xpj66vfNvl2Gv8oNoIg09Qa1+Zjrimkqn/w80I66yqoycpGVDed
GPRYeSDlxGupE6i6ka38KQbsh+rc37tSsyHkom9DfdhuoQTb61cdPJjAAnFmQDVSLyfDCNyGQ5M1
ILgVIMXE60rP3Pf8zKtnYV4jaWeUu4OIh46bikeI+dR2b4Gptkbgh19JLnChKQpB/QovbzMPDdtl
osg5cL/RbFCu89oBmTFbIn0hnQs3TzLulUmIKyXScoN0xuLcdIdAWf6i6QFR6RGDHSZU9+xTv96o
uosexeBlfelVzAMy7395W/HQsRRngT3bCWLwCIWYkvcLjqSZkwyVLmH1hUHQaAQtPGvA8CEz+GUh
AWwdfCiHugjNOVnWVvjzNJusVjnpr2lPrDH2GSvdpc25hm32lUNSUp24W4KuU8yX983RkysB7zcu
m3T1QLZO2kqraQFTw9RQly9WnR676i91HeXT6SELPUySf36OWJpxY2Baz5WR7tpjoe6lySOCsde5
4fwfUAGrp+9sIoT3vujaNzWeF6vJ3NtWJG0L/eSCqBWZSjUTP/1EYVYC0S0GTlxa7aXJ7KKv8Kb9
/RbeV+8ZDEQQa5ZvRJVYdP8/Gy5phdYuc0nDxIObzNl9ExD9NoA5WycjLgLJrX6gPHbHzDIKdrXM
NM7NPkQ4FH2tM45Gh+pRT64fGZxJdKT2bA1d4jmeuh3eiYD5CZG+hY3eIqM1JLBZ7wN5CGKPHFUI
vGiTy//pCYumedRJYEzRlZr26T4f0jCAX0mrf+pQfGppHdWHgnQgOugknF1YF/Q5gmKAbJKRvFsD
bUTa7jmFYg+wVl8OhX5za9EyxMop1yltwWiTW4Jnq+fZSi6wYyG4syxGTzLDJs20OhMQ2DbKMwMC
JDPHarOM7K5eYH2lpvqpzAZVm90TTQKNFSxvd4ovj6LctcadIP62Zd0oRymKsaIgtWlVxNy+VMmt
VswVx3nWQ+QZqLLZiA6wr1BUjOAMk8944EV2a+rPPPN0a9n90DL+g+cC6tvXvV+IvvK+NCifqOmL
m9KUZ97iNTPqRLqnTiL+fxW7Vh9FeOQSFDJlxCjtSacXu3a+iYhWNgWEXBcfT8xR4OYcpXd3Qf2d
g81dfEAe3WRFLaP/fVcneXqhliMtfJcgencH2ZGoC8l8xvxj2uSDal+bQGmJy7GZoQr7q9hvrr/9
8Y4YV3Z+9GAKE7fxnlURu/Sof5PZ2Lfxik+EJRVjd/JPPwhQBDJpNwuIOf9nQbdvzXaqOqF9o/9y
4a+ctEJvTQk2LYJRCFYN+OSqqeuLFJWR0+hV1/ozv4P2ANJHmFn45KKhTEKGLZn8LP2CRNGUKh2o
D8gPhL/9DrtEq8LY80etIIWtbGSjexME5c9ZYCNxGnYCSANmnex7d1Bsd6O1Y9Kg8ySC0zzadnDq
ZkWANLsdk+wnZW5DfC93pHEEFHSN3/A5YpkuozV9D99NynKK/riNot5K6CXeTDV6NthYV/ZK5GOf
Az/+pRPYX2/l3E/0z4Fbi4tWx5V+5NpSTg56p1+DHnafBMEqt9noZx4zCNFGWvR1CmhXzR8FuvPc
UwikO579J457nFrr+YL6xLr1rhUa/bNwBhezhMvgIbFiQZ2JOK4L2YEJIU4pvC8JWar+9uTYQdkW
CaEhEv380rhliNbX39cn38HbRPsOichCpwl8fInywT/Wi7b1M3Mz6tudRVC+HkwVy4KAQxa3mWEn
M2+TFYj6wHw7+9q5GaC8zzYuewVX703fAZjmCoyIPfOt369OBpwq+ks/q5vZ1UmrZLvyLHhl2eBS
+fw0WhhTfFGqhn8TFgIDjisQod4mPFWBWBy/UVG7aK4hozf26x8yQ+qGf3M0zEVUIMw0HwwHiqSB
Nnst8VDYHQgHwShZH34Tj6w1KprIVilKsI1ej2vCM/7/8+cLSND2cMCi+ilvo7MsxDZuhjNAIp1v
jrl701SIfDqGoReS7jn4rTKejPeXES2EYu/EPIhNtQ85Rhzrmg2CiIJEkirznQ+mn8z3O8WgOl/7
/BLxb0eNiLs4KegpuLq5+tJo/fjBhepBuYYWr5ABcjytU0/fhsO+GEu/MQcGoe2vzMLhFJNZXKN+
pcqSUXex3O8T31GGpFCRIDjWxMEQyu6WwmcS+Wv9GPnv2lbqKg/4kw7ljwTZcDhaoUe1xbbTEbfe
rMIfWLZ3lqcpqg7nO/SJZDF5L5GQv6yA6QpVazRFhc0saem4hSL0TiAZo9fpxXIgLKpuruBXBEn3
4PUj7CPRUU6tDJVV+G0Hw6dUEKrWQwFWCzePgCtAdsmaahIT8ZGC2bRTJ79j31mNb3CAUodS2Noi
PoFeKyaob0sZaeLLihILwCw5Anx1bxYSwAKstk1pEen+nVSXeQTQHKV9YTRBN1kRoTOBqEG0Rtwg
xBzFCY/1eqYhSnugOFAHp/9dRWb0xSbDYWALtp3whf64o8KfnypwAWw5OzJp3jytlrtRBWBphiXy
LOi5ZYCRNPIHbZ6pzz1pRc4FjKbJ/uaq0kkPU1mvsYh9fk8Be7LoCGUCKkQHWxAznJh1wtPAwSf+
clx7e2upTTtCFKzw43IhHutWl6GtAlsT/e6S3XMYlSN/K5JVKoVVP2LIocLiABtiFLvRAMv8P05/
jEgVOjBI3+rBpjh/Uavn+kuqxlu4TJlDRqNPZuyAFiQuWafSJ+NQXGHXXv6p4tm0CXPVwo/z3nmW
zPKGKMzHuQQK0g+nkZw4nmogSsAy+m5T1Xv9jssVWJ1s90r9KnmXTzeC7JInqETVTbQKTzW1cQ8B
kXo+u8uoVNww/rUFVmdfkWFFqfHBrr7713/oNBf/29xo+OEuB69LqhkRQxei9njEHdqkoTJkKpzG
eOql/KSMpK65ejaSr4pECbKgUmg/HBfsw8QCJy12cwWvMV8y9TdaliwdhkTapExKNad27lbGGpIb
k8k4Vjb9RHsZGtEBI5JiiLzahbPgixC4S0AVCTnqL/VRPe0Bd0qcaRfNKPyK9SjCCsL+Tkj5RQiU
jGAdSWfR582FiE/eQudUl+wRvFyGb1qR/NQl1ktEgheix0uIp/Lpy0BbRPsRQgcuRLzfp1SUqdmw
IF4A6Dhrc61mmGqTFQrUG1ISX/qQimtJwNUGBSun595BqV1Zv5eBCh8+eZfgMTZrPNSO6EZSOWT8
eygFJSGFPtNsy3mXgUQWJMPvbvzTaOGVfkjXp28xmE51apH57Cm6HwTKOfPNcx2CcQ7eCxT2r3NN
sAWPk4xKFxPsT2r+P9dzvHXCJtmjRH5AxQJgyAtS83xr1ldbGtPzFyXFswIAc18Bm98cnNKlL/Ar
51EOEBS8tx6RJKujOBhCnIhAaKM9zul61cgBV9fUcVwF40rsOvtrBFwUPPwmVEi/vBNYxCQZVsAo
/oTdjsBbPzIY7GBEU7o4B09POBPlCaIJFXMq/Y56KegOIIF6tZzjBBapLUEbuIBLE1yYq3PfvNYw
MfzPC5vLD7jcy5jTuK0+1ltMd5E26OFGYL98iIg5If2XhH5N/iD4gNTlzT85hvMhWlPwCnWz003K
A3MvyBWfCjzGtI7hF13AIE0qfOWi1QznZgyeO8ZKEE218XLMArpamFJTQAHyMA6pgra17FSkImto
WM8zcRlYF9cEqL2ohCJobmpf+ZxIDXUrsXgoMXgsBaOWnWPlmNudc/MUX/u+wyVroDFnkNTxXqCh
h1lG/bpL6htaNCVVE8DhTVwvtzQ0YALrgnYmom8u04Rotf+mtLV4ExBPZ1I15TSQRGOSROJy5C1E
ckXi7B3gV0yj+8iziebO+JeMRvnltFaql3AzlM5mOXEqaEtTBMq6orY6nulquh/htPiaV+4z3V/P
o+3Of8yYG/Mm3YUjDTmEhEouVqgDey83UsBaBqdznWEPqDFrwa/jtWsNzvxKgNx7xWlqVwGOrfE/
IWow+Mt5X3AS4oT5ZFu9EI1buWUS2QvQaksCadqGXI4d+rK9ZylvJWJ+yByPBqNWSSRIXRG/fSdf
kR8btCC5zMsHs+hlJAzyhHIl/FzUSJmfB4WVEGwWyVx8CcWz8Dr5zWfHvTrtZwc5+UFLuf9MQzOs
BNwWnltFEe9a3iBLz9fKXS7J0mliZboXcWM0HzIMC9PtksjC/Vn87WP4Qs9hxOq2rYi84TAyD5ws
iERB8xKvWyFgsQRmdJIuQfg87Qk+8iSWMqGtTF2fTaTNrbxJ3Li3lEGOVNl/TwMH19qOnFQsc2F8
WZDhKyAr4QohBxGEQybr8WBvlSRW4tjqG4BZKpdrKVqg5KfxU7HRzummR/iia7jupHw0mwF9wjpM
wrKWHIw5hcHvw7anz0UZ0wj+RhW8zlmG7BJIkPvqazgXbz80DDZpSlyE4wCuKjnmUONGWRqoOy2K
B1qSfUY7f8eoLE3LjfRDF5Hox2B824bICvC0eKMoqt6FKGy/dIvsUSqubFLzLo4w9/UZ8hOjKpK2
synRd9CgiXXzuWTNrud+JUWz5oh9laB3PAvF/NBKm0OZ9aTMG/xi459n3DZai0RuXRdNsy2qKzM4
SYrLL+avVm/IvJFj2A+SzI5F2Zk89M4iqI+t1Q4QZs5uP5QgYwfpSGQv30Fjqes9OZyN+vs+s4ks
go4a9VQoSqXnXDBnvAr3xe3S9lHu24MYTvmUhju67Kl5iHST/YC7wfTRJHy6emkpp7njD9B3qDJv
AbmApqhEtYOVFcQD7AIwAOLFeEpfd3TVc9OXHjUgvMAe2Al8Zzyxo1xHaFW40BHoGyIkSUgaUHiQ
jKnPSIKOxLNpXCl0I96ocEE4nYaBJFT254vuLoRuxN489MYxZMdC2Xpy+Or3ZWd8JGhLQoSZavWh
ToU+tSjMuy6ffTZ9v2p04CnKIB7CvhFTsKyPTqPmYZ9LuKbkwo9Xje7RwyZGcKD59m08cFqWoUIC
RGv0UQdm6xBgc6UlGYtRb56mxcreF4/801togfkYKHmBRtLk2gviQ8f1yNgLc9KWj4hJtzdA10IB
UERVBGf4cOEwapW+v0G82gy9K5YYjsMTGyTqdPd9Yop/p/poCXF628RVYinDp7+XenoWHALkSGSg
XUc6fqg6ZW/vsGPeFEryd2AmeeUZ29w+LKvJ1SsDb0aPbNewXRNx42r7i9XrcKzZ1GtCFTVHDEyr
/Nx61FvG2tmRejDdcw4CprRjjHIOafNTq12FoplociFeLLNvYS15dynSi4028zntLLX+t6wIkP5r
bkjsheuRBglpEH1AoQgFQWQdXOseDw2c6BpRD0DnWICDmz/DuaHAyoKqmXVedH7ekWyW9EndZcwH
ReeS+e892NTQKaMeT/ftJfTxWXdlXGZtavobogDcGhPX+f8DpR6JBp5y1fEpyhaWRpg9kOHtMihU
EiwulT0CANQVqv9r4yvUOXLNqvoJWP7g6qefJ11AMFdJy6O9r23/IydjUHnWG/6omMSXz4FeVw0x
BxRV6bobjJN3JgmNPdKPAM9XWH/XbtBnqIWVgAlwfCpIWZ/l2FY2acqPTebk3U0ssJ68dNcHaKFk
YHIvzLDUE4vzQfixRF3MwyMbC0odbrBMKM51curArUbULTfTceuq0PCjgX0j9ULZijmFcueU78CO
IOBjiZ8SWOTz3subcPQMexh1/EbM/+KiiesSc2a1Qu1F8g8aLubJWAWge/mSK1z/Tvuj7yz6yLrd
opNB51ymaWWiTNjYRsoarpohzIjIXY8Q6mfeuUQA6XwbE6cdHE2N9KSelnpwVGlSsybxBbIt5Ld0
GWQJGw8hhHz/If+CI6y37Vm0EHQ9DyAgXcyk/LQO4u3gxerPHxvS13NueXfwYTyu7z38r9E9Ym3T
4H3AtjVjFbXzL3yU2KxrQRc7umqiUpK82lk3+m6A0IJ3vTegKb76s7+zpOoOnEli3ZK7f2S2W7Ij
Q1Q9X1Tn/XhJl14y0qAPblnMxzvoXEcK5e6lA2Pj6Vdur4CC/OEMukZqxjT/xPSLSZp7AXJYW1Fd
N6USOIRdW8xNbFwfm453KTkzepE6WWij8O4xSKNbXBSc+viE2BCmNDTbi4hZgA+MRBRYZOk5CgrU
966G9Ec4/JqIVLkNMkqqxeFkhu1MzDRLD1zGK0PyWNuDVFSph8lhtPjmVJoU8Ep0nR2JAv+NB25d
UmoeAVuTyUQ6Ff7kOWDMm7TagjKdbVgNUiN81soQK6cHjgpoYriIR259zx/5OIOMK+ZtCzvLmQ+F
Rwpm+0uIT7kprPIZE8UNltyqsKUbGwrbsLN1RRFsVNZlQes6DMKthr+rdpjEkotMU14CWptOFNo4
YXFFTtea0t8ciBOmsunxTZuqCmvbRagTUJQbAPKNQVDf/3nHlpqYgzYY0sekmdrCInlJa0r9IAT/
8GtljyoY7NcwnzhgNnVXi6zKmx4gWNHh3JWbSxUNrY+Ss+NIwFRMYOnuh6MiqZajQtnBRUHCfgZv
geE6GgmpouuJrW9iCVTmqWE/9NX5Odk4DvZXmntz23Yio8wAz8II02BXZbBF4s2MA37+/o9aEwDF
+lVy8zLfxwkd18x8goozu1a5H/dr4Wn5awIFx9HwodwILp9QBCT42qltr44ooRVfsBMR+oqTxKFF
+DYMMQ2XEpFBRCuOrdVdMMyHkZ8pcUF8xTKveIGr1hNtlmvsfzLcXr5xd+Sfwgud3MVdxnHNV7Qb
4EoBBT2JGm/Zj3/0/qc2o6EWOmjeZuJfQcz7q5RTl5S6Fp29kgfvqpX8+7wjUH1JCoEUJj4AVnY/
CR6CCNHjQXHZgZlBt9VsUTaxrvfLXeUwugYhwyng93FjnhYcBq6dxXwCsVQUPKhOrtlHGJUWHZJj
jAFFETSMz2Ogv6a0pBzF3BX+/TbHWCTKD8Z48ngh4c/SyU6DysOOm0Vn8OmyJdDS7EU7vwnzeL2v
Qz/GiMmyP6HEdkiO3lNXb4TCkhWaxiP4/jPRXBygmZLJ17khkkq40mMh4yj3czHJv6I5opmZiWO+
DDFGtBLPUB1ijy0wfFzyKgZqX8K3xk1tuKeTtRuPIoRRcxs2d9UWFjLHUEJWvxO9eVQ+fJtNLyEH
Bi6MPNPWSL1q3N2thot4qEQL0gaxfUcUvam3+qApsdLK5vpZgKb/nxbONM2h1mvYHNj/yL+bd+qL
hgVY1c+3yY4cLCH/DCJn6/QHvTbF//UWwvTvWnbV1pykkkuJLcV6WcCW9g0WGzPk+0SZpbuJF1+X
VQkWY07ELg7dAQS8QgdFLrIOorVgLs7Q5rLcNusuDllbHl/pA9NUgID6ekQIr78mKOeyCIlTc5zJ
f1jeNdlF3MD8FNshDciet/xe4ofJHAfbHGe8pFtwdTpp8WSsfMiPRp6w7LaMy4ucIr0cugi0KIhm
59s0NyyObA0wYf3iq0IykIkwH1vgNxkkLgk6k0HtB2h/9MqWTiOLiZpfg76NSkGZsq1/d9T+4geH
Eo5URgRv1CKMBFgDEsBHY5i9DUB7vZ/IKy+bb+tL7L7+Bttj4iWgeVwqzx/kHpH1e+wmigA6vM1j
hy6cjSueE7o+y+mSpIb35EMdHaNmRPQ6iVz0sQjGmRO3+G34y+f2+BkPuVtiV5AUl/25PnVIT3wk
u/5GczF2dpLUneE25DN+o69shjXTLVRhb/yekEBd5qLkGr0k6oYIjjWkyBnuslcCis4gj22waEhc
BC0IRS4pVyKsQP4fRU7sq50SyEMZuxmLqF1DO99ywsJjb2H0FqNWcvA9fKwRL7t3Lp7NgTRmY2kE
+foj+GT+fn7VtfI74o9Gi6Wj4GDFAN0sqpe3vxlP9GnFL3jVVXymUkr5U8SLZ+7qtv6VJvKcDbMN
CO7Md1ZEgfe4tm/9joI12LWuCJhQOyO1Xih4aXH4E1C4eXMcjYHhzABLUe+QoKPoPMS87MRyDhXT
3aEreq+COvNJTiCTyBwN7Fxyyylla5X8gpxiWqPizhCCAA3c2cvCMRydLrZaZNTtwUbbEEEb4NjB
QXXITwtf/+h43KzU9/9nhk3CIK5B3CHptUyrs9fqpQzwl02cP+rasPdqgG4+uEh95OPfyXFMqCHE
LpAs0gVLA9blNA3sDd43znovaRQAkDSDfZoq3yIgvWYzqoe81109RngH83B/ddCA7Ga6R+i+WSOG
T7SdKiqQpveiSb0PcXqt/2vgjZzzBfB+roLLAXZBobsLecAQzwa+qQpNRnSkAxH+/bu3UHR2lvzX
rea50lpzzG6cIT3oYDzM483XisZufnw31ksUSOpUPyyErC84K4xwpsSJ6XUfeO5VVcM6+kEJx1pA
wL0L/QU6NQolvW0C3NYjtBijKha80WByxqujyC7AxbpE/tgscj/OnT+5+h14nb13pSPiZ0hSnCnQ
NDXSxcAEwuxN0P6K7Blyl/ztBMrcrDeUlE7vHwf5mkYW5/Rmousunm5D0LPB+j1G8rEkZdSXQquF
QexJOwO1B1x9HzYiFG8DqfLAIkqlLRqBIWCNIfVUBiPfQ7l4qM5W4yEaCx4Lh5+V6//ouuyL28I+
LbszQGhn/NiJHCeReoiAct7ELDjswbZWnYFRXx/Q/OwVCU5/DVIEMD2F/EX7d3QFKsX0pA+0eiX0
NXBwGF0dhgUYCr2Azu+SFWfFDYVB/aE2TC46EMqMN0izpv3bQ9kVSD+DYyp/Tm25HY6vtKo8YWv0
dZpG69ZqxnUKh8WxrSy8SXh7ycJt/Y4Xw6zpgPKWYyfam14sBm+H9F/kGHT4zajGzNbIibcGrr/E
65FnMmMeaP/zoQ/zgMBUQArIPr2YAjDAUCPidR8j1x+5wuYG2DD64cFlhwS4PklfgJGxjrPguxYr
+1GF4K4QZIBXEq3Mw/ugKA9GbYRMmU72Tzgmxjjem2Xl+BundWC2ZOdSSfZbSacXw1L/kJGRH1jE
rHFuAlrjZRrnOQMOQFDdYOqevQ+ihy03a7PkU8pSnZiU1QUZmOKCrDT36ItgUxQ2v5z9EqHP3mYV
ExfRfukUdfLouefgYpYVzjRw0LS/MzeOGwyQBH4JByzM2wDZgb13HJHk1p0csbEP6evrBRrdZnQh
FZhcGCre7xig1eX8NMT2MEA6JtXKZTYzQEgUWItYe1xwLcaDHAlLNEHUDPTTOSvJL6j2eHoTTF/n
sqZ38Jb6lgQSC7cApihccm6TZL5cEoqwEU1DiVPznq2weukW9xy9FvZx2wqTq12y3wCsWWhMZ0Wq
pt2MaHHnDlsBu0hSHPYorxrR/xUdSptjgjMfbOwrnt7B1ZresNfH9ljv9VbfKTTXegvuPzKs/ExU
zKGHRE5KexRl7tdj70LSwiQFSjYhw+N9aWN3ReOApPfTSLPvQIQMHBAwxGIPjbmuLdPMiG49IEVy
9scaX770ZZal50JlOCcunqbApxvgfhvPlL7ZYJl1va5HUlQiZpc9GC01UPaW4M2iLoEDzHxQsNA/
nhF/fy+ietAt2O80H1Vgus0Abjf2qOF1Zu2QlLIy2m0ycCPXyVXsQ6SQT7MyG7ddplZjJLcYJykC
fIljIUgWn8Fd+3R41C5z/jNFDHDrD02HXitQmYOf9QsNOS78Yeb0CLyZwrsRDMOoFr4p8YibPWKl
/bag1iwOzTvhZKKsGPYWGhzs3b9wGrwra6xN1LFEdJS70PdeXSjvJvXc33b8EpJLb9XoP7O1xvks
ZLD34J4zMG/ewTfqn63RP3BZ2ZrCO+JQK5MRz2uhpyASnC462u8YqJfIguT0yQnX20dnoYJfcbST
C9p/rVv5VQ4y/G992wsMzbcWki4r7hqmX0yz4oy3wIpwrTCwBJu8ZVi9Kqa3RWehswK+VUeMN6LX
83WYuGIOYQAShLXegX0brySxaxzIp5ZE8OsyG8x2olyEu2XUweYND5z6Q9UpYuhU4CJkGSn7nUkU
kn6e+xHu9aDqOPRjsqI96Os/Rc8K+kkwDW8Cj79eawPEEtN/Jaz0sFlhZYcyt2LQgRnVMPUPl/WW
X6ZbdiXeWTFa1IHOP7tWED2age69dkK+owtDoQqo8mu/yuYFhD6eW+9StRpiAQT9VSqZ3KEdh37v
/RwqISymuaJGAZVQsjhHsAYwOOZdLC/nufSdOCeNS74qxvYrpN5WvXaa19jTsKUL2YbEmWwKL2+2
pYUd51EGVgYUv1Pckj3hp6g2EE/KELyvhZDso5Uf1PH/dCUs+fSMDDeBBS33cHFT/aVjcGMyLnik
TuJkHxYspKXps7WVULqCFEgIpNY6tTw1UqKNRr5mHfO/R3f7fD+J4OtacjkIfRxK7Dm4DGWTs4Kb
/7pwKGQN7GIF2RLKBUjWm6GMvX6qgIktDqgfnnblyHJ4ib2lHq7ZEGR4feGfkYpA3X/eK5yAYPPY
7IslgyqhHwJG6I/EEErYIH9wDbmCMZ2zU1qEco6DSkPCSG+J9nJ3SgjNqdNeG4X7Uo+SzyFQpBaO
eyeu4mwZkCT3zVwRZ7hpfYyAdaSNYeH8byYQpL9dqU+jSVQHkEsvcoukH+Qjfn+RAWHCE1cGnDdl
MI5+k4xj9vYk26Rz3G35vADyMjhZBV0w1hKExVA956wJvlRRoK1csLIj2lbBeOLrpN5lG+qDlrb0
27IzJUuVHhaY6RmhEkNOvy+v+/eqxIkOd5i2cljYc4lRiuHsl4l9OXjVJOgjBKUKHjaVwoyBSLDk
3/a+yk58YLdurmXVqiTF8LAaAw3JuJI6GPiDf0ZVll4f01VJJTNiS+TpcEXRzdSzJWpc7yIfWk6Q
17ueMxhYg4g2ymTaVNlsQkv6QnDlfH0Jj5dFc/rEcPLeq8JrY61JRkRERZGzSwCk5hXGOnvzxz7o
iA1ZL8xIAKRPjSqGKD2LrTgYBlTjLE0ANqNu6lUX0jzU6lSTzfYgw8gmpo2F8ibbdfqfVza254HB
qQwWLfJYyvrJ2GEdzoaKBGVXEap14H6eL1N0mFxCsrzIPdhk1KOhb1H4xYdOCgxOEex4UoeLZC9k
M/ShuiupleZPPC2UBVHAOlqEo5GGjvqv3tXmy+p8xcb6AyRGDjYZkYPFUUUw0tTWb6tWkaSf64+5
JeIS48+KF56BtGYo+4JV8EjD9I6qFwBtmxrUKu120tZzFZTSRy3W4fJldjmgcslStxQMlPRyneEO
oJpWZyLxPq5+1eC7uOXdEGc1UCzh3BO2rrVHh/wGylXDpR9MMceUpoKOeEQJxojOuhLSaIRPwLlp
hsB6G2fBscLtSPnYwyEf9uo2qmdx6DWhmN7T4F4LIDWAS/mGAe7qHIoJyp6H2r4AqCDl585W5U4m
796odTCgY+OnmSoxVuLIwWwM/SmMoN7gGcKqWuZiYtQuAo6f4WNz4jmrwxL+KQk4RF0LuH0llfbx
lmx/JqQJzryOnHcS8wTkLNME0B/i3sIZMzva+a5N2Ms3v8sMJBMpY277zyYaYfPfkJtXUFbXSiFW
PEX2jUkzFznnsj9MZKb9J79saDZN4DCsUtB6fyJSZvZnCjDsqUc9/DkiXY3jZw3m3p7I8IyFEkUg
r4Hgubt4SwoIT3ecNcjU2u9MsY8rUYdwIwccQhiST2mu4fRR6kLMGEPn+6GmP08KzoSp62Cnj9To
u6Nhc3A7bIPm+DcCmDWHTxPaOd9fxC3yFPsOISzAastS/z/9LKQdlQe7cCMs90atxzwHJ4yonAlF
DSdxAw78lq/iEgzoW2lvwopZsKI4wk48b4NuIierggyDNRaVOeLopsqh+yTP7KFVwmakCy4a8RTS
l0E6hTuAxBtkkgBo6d7joLwb5hDM7XB2+5UBCuh0VWjsV1JrMm2mpPMxle2HIhg6BAxhARNdnGhB
0rfkuImUu+DG+1r7uaN6Lj7DiDh2YWcz8VTinfSf61Pll5Yr04nRbWGxGJccMOTKW05ZulgbfJNC
Ut5rwkQvj4i2D+hQ7gB7FpX7XuYhNz42t73WRX3NL33XZJLp6hac1IeD+QrfMe9pu2IjyWCLrg8O
k38rEklzSsfFr8bhLQaIgtI+SxGj16AMFyoim+28HcX635kVF5AJd+UfOCJiG2066Rq822L87xP8
z2MnrHRbEfsYsvCm4xxbWzilgBskIPDIoWxbLwQUWhEqcz3fEPVlymHXpxleUcaQOVS2ODJZaxWR
iJmpim6IdqKqJmt/FMGDnfoRh1UXduhZ/b+J7EtUnwyrc+9uR4pU5ca22j9GTJ8ERgf4v7fHaFiO
e1UccZ1DTm4qoFu8+BpUpcn5DqL+fzzoUfvgg53kFTOzT0N9tWdVRHrCS56o8zta5iDzGKd3sKsm
Ewr+QkJAAqnT0947Room/8PuqgunqPB++hitErx52n6q/u+x3hJQar7yvQcK7Or34BWBbRwRGrZl
dKHegO6mfpAntNEELuMycbMilkhkCBp4MQlrjEqD/0iC5V0mlmQrh3S/DrTk2JdUbXHIO9k8QAzv
xn34P/Msf78Vcxk5XgAz5Vqzvqla7aiDeBr4hUerjfU4sM622VjrLYs3oJtWsiEX1q3x2K8gnLet
n05SLY+Fflieip53duZKcZi/qLKqdMN0UBH7RL6DGLRv49yu8UlSBp3qhGy4uHvK6mZWPPlLhh59
BpTtBojiEQffnFDTGwyouOI+E1VLNB3Jn51vcNyJCUCjlpiE1Qvbnhqag+HLSZKkKnmyydkjF7qa
2vt1e11ulVADhgEqqup2ss9nMbgpwPxbWcARIpXE6o3F4rPyswfftmyTH4iQNVCmlhMVmgKeQ+VC
d422qJIn7cnFEmEXqvJEv4oeuhVtEv9SZMJId3hlDvzUKhEwx7t1PSk+c1FIPcBDdqZmN0YH0125
3TcRHpfJJgG0Flx9WgndvfKbbTn4tCyh2/raw1rLmbn4l4GIo0qTJ6ojR4qEIwaaAyrTMIk6Yvcj
aC3ni4fa6eIIoLdCqVtx6+1D74O3zFT1AI2JMVPd/NaACyH9sACSPR/7r+v52MmFNsNQ7IsxeDHQ
cpyv88C5JLed8r5Jq/Pj1hHDw0B0E2Z089imb9fJHtfQBMK7LxmF3Ys8q1Ir7R94KjHywop4yvyU
hJQxrWcmfLmizZyVhOG4qS7n0KRBdHTRJFIqFmk24IPZGrMxQ/uYMAGJzppGcPJmJ+0EutaUN2Cz
jJZs0+yY8ah/cFNWHp+HMbKdri85cyBEthKOWB2RMaF72wxJLBgml9k/bodNy5E/eA367F6DVX4K
tWUPORA4/DjZV7/78z5SYeWpt70/REoOPUZPXvMpJO/a8DQkHmRzPDBaM/jRby1jbkebjLwWuDY2
v8Xj6AarFZ8ev+qvER+Z4ITbDlByY30TcGPNvkZdkCrab54yijQzHNwJ+6BGNSS2Jc8wNUoHng/C
mS+S7Vi2zv5m86Ck1dMoA3yJApEkQQF13+7J4RMoIOr21uLekh5IiuUb2kBkH18Fiv3w2RoLzj4F
ypBXjO0Myv/c0hm5LhCte9YIcuemkOYwSwoeLBcdR+v/o0VUxiIMJtFurOhcEhWUWd2A7C5/Xj/U
3Ozf554cTUINnTrPWp5z2cg19zYSJy1fuDbPRme6e/pmLnDYsUjhI6EyZr7Q4OOW8uBTs6mrGQn2
A+CNUfhwnWgzWEOnTlGieQ2VP1vXsSGjK7wTFC8CWERUxlOpd/OxdNEURSxqq14f4xOw7MVk00eq
r/v7ywyRs71GSkj+wfBCKHgt9pBxMbZlKKFG3Ay5QYazKFxHdPDYg0ePhCAXofVINBjchNf7S5Z1
Bu9+uFIJZZ9gs2QpA/4QeZ+0/sR2/84e05R8lIwbK/UAGynHhorP2ovQyNvUPyezNOGAHFtMvOJm
w83VBeuEZFHR6kQKh2iMK1gHBOnFI8y3uZiyULaozU7fRQoNp1TsLmj9Tl0jJV47A9SVoFgY2IJW
GJAx7blh69156vVJA7Deb4kDW0LSHk1Dn24IJkAGHwFRq8NCc35qO2UkhZVQJSg71CdtV4LxFxws
Kyh/rj7xcvi0VOT+AtWF5OG56RvENjqsyrWxgY43Lc1N34e31Ps3Ke1UmCrmd+C7GvqXADSjh6I8
2QxcrBdHUZqSm4w26XQJOeeSkWBUOp6U4jWGWN1wj6L7GlZ8+SNs4lc8ZroPxSkUKj8Pzfqrr5FR
UMRAB4PGizm3CI0+L0IafNXmISsg0f+v8W5kXRexDLS7RpnsProIDUl9CehGSh5gJ8aI0SpGUuy6
koNsKks+vTNa33exjmUlaKXEJfTHMztRAat+mZMEaLkNJnYtuX8XUWSuEDH7BfOWNrvMcrAA7YpS
m1Hd58nLlN1M007q9el1bDaMwZ6b38J8YPnlXo2kX87Ka6cNvcEci/3kCrUc7Boiyq3SLLIwUW0S
JTWYzBQEPjx4rITnS1zOJBV2sULpJmOB51LPJSLYrD0VMvbB5qSQDX5xZuCZKOyJXOoHK4MKuFtf
WfKNUnK/bmYs2/tWyt8E6bN5r/pl85zBfGdQ2Qb+HlU/J9AMRhWiOw8/vsRZkyYGmk99oW5N30vy
h1o5Gmq7qEBqYWdSjBD3QJzqfLwmQyno5t9fsSuL1bDMH4JEM10wCW3xHaoUekyuNn7xXRcpDBOO
nVxhzKNBnOmsAvDZLlN8iWjcKyDSqgcqHC/c1fHYfsQhLXQFtp66OtQbcfK9zLCl+gMBSV8BL5rM
j+GXdZuRS/NVW7GRHG4d8G4jrMhNHXuMk8y7fezQ9CsvRGSmdBBIM/JNk1+EUIJQqGtOJQbG/PGy
mfAOFDePlLVoZjJCl6AKmdRJHiNde8qcL7iPQqMmGYQU5JzVhb//bKuo7pa3zYofXOiJTwx+ltZZ
eLUuffXlgK0fmltXQpNoRiIYuZ+MBpgnimRm6QiOusxOQdKjTDZowGeWfSW6QLDOiA6ye2sZvm2T
O717WOPQAjz6ws92wjXyfD5t7kQfXPsyhs6gnNyiA/VeosKsH13boSDhHP2RqkhwMdEyRU1lZXEK
TL1KmING/+EU4jEHXq6PuBuJRaS3/geWy0ieGlbSvSuuEHZaLfifPtmBe/fsZyaYMq7RENoRRsOl
XJEAq9QJs4zJ4QiPbvptlXLeJGbMil5wdo2hsDg5BnB6Bg4KalzMQZH+dXt2ymSxg3DobCj7CoGl
gBk2yVzyXk2Bzd8y5elYDCFkwJPKERhBOxHsnx7vR0K3UmHCj4DjmFOpTFSg250cmHMvHlh2fOs3
Nf/wdmpqwnLhUhrQkwUicgvloUJqaZqhrqcrXRq4YiuZ0Gpixix1+C/KixP8LnxVbB5urUbEDYTj
Fv3fmfof2zQz+rPH+DkXFanzMayakLdv340F49383ngrRDiAPgHpLRDxM5O0mbWYcJAYzPeTD+UG
T3TccrijrSRXFOUoagy6OsVp07WjKGUvufCd7vaLDVFPxwdxZ7u8EnSkqAfEO/IX+QCgvfP8lAIe
9kJ7yqxVw/HW7o+/TNCOZ4FyUvne7d58UScIl/q0xjwA5qBfzFzgm4MxarW6mm5VWke5KkdiSW/j
TpbQJVS8fgW0eIpPKl+4pJYgnfIpnU/AbdjA0nkGuMw25UFUHpRc2yy4mYHvfc87NsqUJovrNAnn
fBJeHjIAWQ91mSN2hNa+ytBAgRjIwWy+Uqf/Dq9T18Y9j6v/J2aSwPQwJnuCsope3O2azzraCf2Y
syCEKC6QK+szdcGaKSRC4oHEBR767psrdgXha0U0ap5+kg0UnAK/i/fdjT3H84C7ZO8oclytBY0n
vcXqRahramKuPVS+h/viHCcrK70Nq4NJEwoqXRm+/ZwzM0HPqYynzHwwDTY2TJoQjf8DWo0b+MUJ
s1beDGawP4MH/4RYMIWty1M/lhbtyHzvmjYzWRxPEIxaZ20D64ksn36friHdhKzORFcBzV2+bDIv
6Cv+C16wn6loo68QYsk12ZrKTM8z/M/0CICpEDi5mI3iwbA+SxK6qv5zeu3patOdDjSviPB4yGHH
QPYXpl0yc8sVEQUvY68xZRQ2J3IejXQF3B1zN6TZWymZXDFVeJSisdl7ViTk0yH3hS7OTrew05Bw
1uEBEsDM2np3MLa6X0PUrQOaO7qQAXGWV8Ld8j9oqgY1ayWMbTvE3g+5FhU6JifeKDnIAxVx3Iau
SvHiZjhynaVRmspaeGndCn9I20Ibjb7AFW7tTyKPRTaQf4d2TPrEIAKlI1wpWVFRsqFPYr7W3pQq
ewsqufO3dflBqBLvw3IN9welyrre/0eyKp/rHXVQ4Ihe0aY3WzzLKbhppegXKPyewLrPRWlKAwxl
+fNQvt8xAC6/1AjlM3u/ddbGrZzc65NpPOD7rpUFyug6Jeh8N0+9dqsXS0W0JD1vTrr61pfEXM1P
kSw5saYS84tMJUhmTo/GCecgzikRxbqXl4UROBoRWse8U3ROwRpkQn49/ZXF47mAZac4Qma24a4g
1X3XA5LAoBEeRsXyLfeoUExBG5ve0uHUvawWk+aRDG6WW5nCkXMrhr26jo2CKhUfGXFnqXDrkb8v
0ykJ9uP3Uz4SkA1nRkUFr73DadBbVu8qxzTjbN8SfgnIlwIImael/AeV86kTgiUtEIh8QM0ZuB/y
ggii01AeIJC1ffUIb1pn8wsmow0GZbG5kqWfU6e845rE0N2UItfHLjyiaVj5zEvQwbDXDWj8mp8a
RhpmqvstoWiR9jVphltNMiN0ltZIDHQeaQ0dbeUmxh45dA9h5Ht0Pc8EUDp6/NIyKcHVTVR3Fhgp
TEPzaatmPC6M1zoVL2O6IiMOcdGbUeUCQROl3c3MQ5ZFP/5+QWdPRKn9xobLboo86tLctArQQZrb
ImJluFN0ouUKJXf5hTWVbVEPDZhcCEHKrR84ZORA9hrQkN4FyvZ5CPpbEepqX7Y1X19kixK76BeZ
9/dMbnwfmvO6vDgh6qG60KWhYJyAVOcMtiS2oT8PlK9TBCVxB4/Ks9IxUhTHOc8y980KnSjSiHYe
V4u9MhsRS8UAqs4jSrYIxEA8Uz+fR3HgykP8sQ+0b29ZDHXg7auUbfxJKD/F6zzrbd4U3EVgE5At
2QoiDdAORiMV9FAGanpQdaWPjl9Ipkf61GGuN5df0a4C6B+7lf3LBSIs3l85ulnDAsDbYRaQR55m
WCbU4euSTq71+BFmHvmty/6kvfnA+FYkvawws9ZZyq4fQw/EsNp2/EoW3sIakVrR7iCj/qL7OU9l
86lR4W9+LZS8GmTkObEoGgyskuLE3lrJQEEjFnM4i8de3Y02axGzrpuCW8wc+J6s1yMasAgOjNLB
KpClKj0xL0ywL+VBSTSLa2JQLgH0+0kIBRAfzemOYX38J1CwxUTCQF1rdz70MCCEfhh9w2shIRvg
/cnb3hQ7XwRbNHTHI5OBEwp9tIMkvtqTHGKWurF3Lo+P2tuav4rObJnN3nSbcMyOWETCAA/lWBgb
8R10Z9Bso0erqUf9K1ELnX0kWupSAcvnNqyVZ4+C5R+qY14INGn1CM8AlLjQ8KgO06mABxr6eIH6
IwUk+wGq7NYOT9TryAum7LFzYEN8Ih024awvUUGPE+YNkYFAowwFlUYGaAtUjKTLReoCAx7iJz5z
7FMcQXM/4XwMt3VLqNADHv0XUuViXtwLfRnHft2sD2imf1rcsuQVrjOy+43OxzadOM9e+bOvymeb
A0Fi4+V9JeiRX05HqTTlJjRcyDO+0sG4F1RTc/cpCy25HtrC602JE8xqgHYHgTeDQpwY8BKefyr7
36Y4fWDbDF/Ruoau2bGQFsjQIG4rCIpb2vVrqxxShPI6SFVcy9epATEO+QCK39MMskCXIs5B+jTC
qV0OLiXCjaiTH9Eo8r3UuCUdn5qskOGA7jffYPe42j87EjkduIUTsj6z20Kt7VwRt1JRy4WuWtum
ZN1tnR1qP0zOE9nEnMzCaPtYgVwahfZcSgveID+6It09hd4FSbJBGF9olMxepmkV7bo8mlYMcw0n
LzvSW0FsLiJsyI4GwhqRxey1DpS37r4hXY65NlMzkLj0STsnETJIuYv3hT01F6naCtFJqO6wZn/9
4UH+apGT4SpDp/nq+wlyss65GCsh2U/OKnA/nu8S7Qn6ORzrC7XpC/qUWf5w2yb0LxG/pDAhifsm
hmg/tEt9iCQo6QzCLA/OqakljSp7sbA8FzxXtkCahCcVeGqU+EpMC2oPbfDGOIOA863LpEBFeuuB
r9JpK55dQY2n4kxN5ZzIdzctzDKgB1Rw9exDjq7DBsb7MfSNkpPl2bbZr2u+XlWUuI7pF2VmF6cV
JOOS5dy9EsG/C9AsM9CdAOvjg1EmKp6jYDY90qJQlnOPTqbUjNKYb+DyK4/Nc27QgOTHylb6JSTl
vof9VsQYkVklofGQREdJyp6Igg9HIkwOUDOZW7iCy3ZKmyLISTmAiLhzj8gteCOJ6BxNwwfu/E3D
VgQPExnUWqVng8FhfEUbdmej2PcmoFyKqScLLv+yX0cmcf5eSNgWa8R9zGPi0Hj1q5i5vN6HcQs7
x4IClHec1Nh+/0PJY4m8+mfI+45n62zOkt4/smSZZXQ63Jj1XdV0nFl+Q1DwVYbQjIwX3LThOtMS
ZEmz+L6/Ay7ls6J81gNnDBqi47b7bKCBEv5Z3fl5flALe9NUVuoSQBIJSTttEHXHeIhzXn+3Ba0a
cE8CZw+/ByuW5ZI+SP88VPgBv3ckdwUOR+CTxzM9bFdUKk/u/GdWvaghnnmOaqX9ihsNDVizv8nL
2EqArQTRDROa2WzKQnRfL3OrfgI5jGzVTim4GRkV+j3+axVIsXezdstkeO67o1ekeXgELOB7X3kz
w1L0BOtEgfvyYHMqY90GZMcgKNMzrsvH+zOD5FPBsdKYPvLf5S+U3ad26GbdqcbsR6MqawmijltA
VOD6ARlsDerRSpyc6kKoBCBmIErw+swy+5VYJQP0iswEuqoBkhhYkinOTzCI0PsOMDCzkBPFyLmo
oYhHpPfTg3g7R2XnfbBd0jvDpdVTi9Ut5oPaEte+SAMyjdyvSdIeepkdZKk7s6HGGKkSMa9vd8Y/
eDlQo1VBRyjElYUXTk4epOfdRIuR7hGVZA/duq9ZnefYoJ9gQHQhZ3P05l46Ma2DjB4dLEUpQgMT
LopvJT3esqUVQ9w4aFp8tBhEFVXWGG04t1BUIJiFqOFxqeR8avkaSqozdXR38asmOgJWI359AuKb
5xNxBJS4CPhF/tYG0b7BgFKdtIBUW1oZJ7BtP8VQQdriK7k31lQwFcwN88NjWDQb9VmytF2P3uJb
sHW8pJWLc/vuarZyJAVifn9V2iz/tcOsnWdrzihPiHm5mZMfTWFa5kiM8u5L/z3Hi0cFsMWwA29I
ZCzbaIYKpAjjnfdhECdkCwTsOVj8wEHptmp10xBmAX2e6PU29LkhaLa6Z9133X7hEk/zIIb5348S
6micVj/z0qHIgKz73xgET2R926BGRR2SjTJlmFCHRs6t3kj5OClTOcPKk6raI0tYh6bdAT3H809d
VmIu5k/w9/wkmkUD6HsDhnkhmgbyMFxTAgqsrlLoavXec6hh8H2VIgnFmIco4rKYlL/aDXKxOQM9
7RWSfgV7HcGgXYXGHDGmbR35Q0VTTcZs2JPyV/hPoFVLv9d8OoDhkf4zQ3ARfV8kJIc6n92YybUI
aYV9VcwITetfTs7pVFnrPXfQttcDvMYXW1ocTzG6iuwp49YboY1ckmpJZMIil9zFBd3t/AFDirw5
vw7h4MFZSXf09TZA/UkNGQN+kVjUFkC03EAbVvNGzlptglZSjleS8SmjBCiUP+7zL2MhcI/Amr6R
quU+nf7Nil1FIhHPjKXUxgMP6gLGrvizJfHq/zjzag19tYCfANtMLsxdcuoSZ4oIgJHJv0oX46ba
M1KGUy9iDgcJfWyTx3A9K8oP1FMbtIHbjPHdFt6LM4y7QZvIYOKpMPPSWrJKLOzDWk3qd+5b1wvP
fbUyPzMew2JgjywNkf0YZPME8t1MHHBbt33GrO+pBVFBUh5LNuoCGSxUGYfJzErmrxmhGkf1/cBO
62n8+hmDHYgBlC8fJ7o/kQurAw8QH+sKHoObZvdC6aR4TxxaeG80aXcft2B5fFFkF3LZq68ffxwA
PQuKm8JJpGPquD3MPnR38uqD1OSba9O9cJJfa83KSjfP5wt7zkCARw2A0jiDLmR2xkFLP8nPQhzw
Pd2XBrGVXAS6PDcSfnRv/5aEgRyECE6+/qsXuH/BbzrhS/QaeTgpT5cODpnzjd8Eza4aKpMHEmP8
rShLLK41jVpXzOwIKVlAST/BxKwIqT6Ww0Sw9sci0e07ntJ2aZKFCNKhHmkM9uwefaEGei28NG3w
C745GgWHqwtBOQwA4vPBisQwa3ybCGKHKoKM+LM8KXtB79aycyHJhwf9vg8pU7peU0ryq2GUlzI/
JsRY403duq83uLM51Kyus7o7pSqFFts5bLPoUwza5dknDh9xtpYQ2tIunZV8801bzLgVl9m4MpeX
Gd60m5AX89wePqrZLd2kfw54ngOPowP5pgyrdEmmL/I7kR+J8W3rQ2tJdfqt+Tu62MeKHhLlyAQC
D0eR6HOpWYuB2LgldiNT+v+OK6bvdLrg6JorJ3zEOmUutqkLtRvTK4kOFJ6QNY4vMolWCp62fvry
BT6dXFvFitOg186ou8WZXU/cCJx2Y5kzYaoFLknvxeuKA/kJptJpzvJNH2Ck0eOZuCyOSkn/dS5N
A2UcMH4nYJtGqBjuQ6OIo4PIfCBGRCZFalq2iaJcchorJa1UrCywb8LmVT8rrfXYAooW5g9MZpXs
rj/YSXbowuxuQhtqN+CjfetRB1P51gjV9Dqs5UQajD8NHj3V+2LHf79b/wr0fJX1AtvkAjRPInMy
jJgexjPUeCFB2oAOTD2PAyzAa+XxYDb6EfZ7QFVCPSUVksPruPd2a8Eg3jeHQI/UlXpaRgqfNsBS
uJc1BAp16txT0KWQ/tJSAhgGYQoaaR2TH6iIUbaWzIsFx+WFroYrELrnM3ahIxghk/vn0MdC6PFT
zXiptWnZXqUhVdGvPWuv4OCyvZGPXGhutlOZk9iAJOW4vi5G78oBgQnNEvjHBe9n6Bu0pU8QS1W4
H7icC93/hOfJMI+qDsljt7Re9huOjwN1IV70TrrYt0Ek4PxLxWRzBZzY9kgkka061hSeOUenZzLh
meUfbUbqSCTCsY8u4UE4jfuGQnhZuigkImileiPkoijB15lq8Un03NEkb5j/yBuvQC7m2i6zZhi2
CYbhZdGFqZ+OnVmgeRVgyR17GaaK5UXBpQhWy/XnPmi7acbwrr/NrlLOW2/KLWpP7M+OkJWKpAoR
Z3qMII688BsQmnORp/skBRuczLpOUKw6fGyeBedvRQZEXDKkx+nva5Qni6DdwWWAXRd9ry6wfd+d
ri3Pt5T1SGHfQVHWwaDgpMETfcvtEvTiNcTOpJmODlWG2VNzVYtmfKkje1zkfPNdMUvHnRt9kyx5
wikIOniUhxGzJto5rBrn9cQlQnogxYPfVzm3+Da8FY1DGw96XNf9nwMClmPdjUd5n2f88u8+qckk
VNVwV+s3GBv7M/etz0ZyWAhEysoePoUztxtAppzqwUVIYfHx5OfsfqUYbiAxDIkbpW8tXiG0mEJI
TNdqo2fQc8MQexMTX2pMhRnvGYzDVxgJbtb841VaHf4xms5TeCoM4M79OJGeu8vJHMyzcEi2h0ZZ
YVWnmvWjcOfjB4LarXzmUiMzEhpzXFSmRXwzkW8aDzyrZ7LSDGQZcYw0tiOJazOW7yOoHT9BctoM
r7XmzUHyfkvzgbc2KGzkKDKUwrxtApaUYfAcc9iUDyvyuYL3cLOLOw+M7D8MPVn9UoxHSGgV2YIs
6YJkmZOBEYr2pGVoJvm3oSFPs4PbzIzHYE+z78ONnGWPzWWMPqUP1WZ2Xlk07yCa/VVAAlHC8hVH
ShLuZUY5rQxU25tsDMjZiZIMKQPHPTbFhMD7RmWW2g7eP7yYTRERUf6VD/LTBpd338DM7IIRIHil
iUwy8uURvN1w39StBqHLVDPvaub0pxJq3epBQiFu0lqdTaE3Vu6LxtOQLYux7O5oYOfvR6pIG1wA
d2kKuyvel2tyTH0H63Je9zKyI1+hiYNN5/3oNaQntQWA9afBaY2cN0gZM81BI03GSflDHuZtggqN
cti8eFfaqzZ6Sxhau/vR3HlzM7lk8sU+WxUqv4SCIZysuv9IqXAxQiO9vuv/NYjqs7V3/Jf5HG5j
2vZelrZcwMPJ4/icPMfAkmM7KCsqQuhpJN6o7dHvl47rsLmZXW0ikifxYGArSqF7VkCQ6Mc+EVeg
y9HQgfRftaz8tX6FTr6zSt9lRBRp9ZcGzNO6yegxxM6kH/cB1glq/vaUyMQELh+56NdWxUdL7bN4
VbOcXnvo8L5CA1b/hS7zDjepSjIk395ZJi16diaeMhksYVkI0CqRkJq318iyIFqdDnHz0CMnJ1Hf
riBIh/ew2QBEXGePfTWQ7YwCFKdhfCIHu4pkptyQQrS7BzcYg+lb+TpnvPK5F0Nt6iskA7xhpcZr
724rDueyM+tuf1y0WaXEUjQqwWF9IYos6OR+xsz7YDfUpcWnfdxbY1UOdr4NOCZoQ0MwDeDGHoCF
wZU4rcdvTc9XnTJdpYcaoH0pM6/CTHOFiJq7blreN83W18j6Bl0GSO8BL47cP7U7kbm1QozRAcZX
8ddt6uhffyEqNdqjOf5BOTTDgxqUmvpvx5wVjiyRt9lXx5cjv9/sTPjbPT4gM8ddP7S0wWYp0KxQ
VFxe0ME7dlSzU+sFyEf6kprgA8uHb1freaDP4YEwNQEVj3Dxj5pfdhTdvlBDPoQlAQZ3DkdUD+OU
HM7A5M9QpVAbc010/G9sWBvrg8HlXaYpUYroHOR67Ul8aqUM2QsYWr+I9HYjBLenA6EWXinqxtaG
6CeM89PiPGSCrHYT+e7q9NGVctX9Wff0TZYRO80VWvJl/SOs4ullOCvlNLbthfwNaxnTZCU8niq0
FLUiL8GwNOwQrDsd+11iP+EhF0o6AOCmfFkyREcjiE/5gT6WyS2JDw54WfKKYXDW8NCLiGi3R+GN
LFpA29xuOojtqcFXEnnmZTovnX7XT6tYHHUOZ5Vypv2ljPtEetT+eH1Oqhi/JHMl+2HNhuUKBh6K
KLKDVOCEyne5KYmus9G8PMzy7rqp4qvWSQIDdtrsX42K/9vE2pHIUzJMeFXgeR3/bxvPkUc70OqP
wBztSVpr5d3FViQi6LXI3VGkE7BVDljhe6W19496ehjVyycaqomWefI/fKOH1CnQs19mFsQdh01N
+/RCytL5SBhiwTMy4F0L9+BBJmM1aqmO3wmJ3QjWcuq2pkWhHQ1HIPAxN5o/GqxZ+YzXO5y6yXFV
cStkIM8Sym9/A5U0OO0BoqiBTUFM+QiZQcTvLCpby84A72aM0hKYerM0VNHxCHpVj3Hge3uYX+oI
T81ZmojmoIAP4RPtwRiBw5TT959vtJtBfNFyfIgCftC+s8j/3AbgEetHInagdkYlGWC3+a1uvVFg
iDwzMvsGdGrMUUU+oNmp2Q2zuhi14XNr+62AJhBKG7F16fPj6AGSaDhW3dm5xpnXZD+u4JtDPZEI
w8l9oLQCQnQi2z+gZq+hpZ6Np88ieg7IrRVtpJEN/F1iA3IT3MO52qM/TjvevrTbMb56jbAymeSP
YWigGPxbjLtV6cQ30oFyIRsHuH8K2Q2dubquk9VatCC7JCq37SxPcwkKNLz1Z1AfmMwBByfnxkTP
VMf3Kalbhg82amHGE7FeHExt+41xWw+gar944fIKdhOTTbpuBOROJiua2BHiolZ6uDrl1hrtlh3X
hJd4IhGJ3sR1+LZvcFC7nkPEoPS43aq/QvAbA6VkYpearrU8+5Y4Q78PFlECXVJBV69eYMrFT/cS
Oka+ChSIGsyRY8NXWwTJCpGPpQV4M/YeSCAcDWfFSAAmgB1NzoKYuHjZyBH3T5CjYIkbb0fOpdUx
zamVyolI9SZ+qxaSYGGnZ9nCS1QfH/8cZjRb8+un56RoGSt4kDlyzAHNtpMg6f5LHer4doS0g5WR
HXr0hQtaGDuaxZ/9B5DBpvp5qLr4rT2mTj4eoyy7sDrNTrroCttHKV8L7QgqbFHD55tmRd32kdS6
vU7XpJDfd07P71rpLAORyG7mR0c783tk4OuIKzjJ+TFVYjJk3QLcwqBaazMPgi01Xph6N3YNJwJ/
6gSjifww/p4VVVyn3xkkDBnKF3s/EWi9R04Aqu/ovOZKJARAKsrp4MqxqBD0XAe+MBA9SoQQ9Vdy
NLHYX7fg+EDNRDPczE2EL/HHAa4+AIfNsX1VMjuK+w5TOLa+56/FhZmchWTzxlnjkbZmMZIuv0yM
A2NtKJGeEVKZvBwHe51A1MsHKxSVEltvdcPctg02ashVenU2XP/D/Aq4xvNVgwSZM4c17Db1EtvY
+XXSp7U7zimS8HJ6i8DvwgzCx6UE2aSOamLhZB40iuxiM4Ubupp1SMKFtvOV8jYsu5kqOeekvdDu
aWsLw1dqpx/n8QC8P9dekj0w0JALW33lfvf5gdFVmI3BNyOS2A6iuwluYfUZ6TPq4xJcJjHVgd3r
yYxeWxcgqvY9dYFT46pIyaFBps0/xgcxyBZbl6mWPxxQwvCu4Dmb2a2RmhdXIGyceQ3AygrImcYi
9mWX88d8bbQlxgTkLGOa8MhshhEF5QE7u5t8shbdeuq+26u5HiZCApH5dDosoxjkPN/TIqTmntLQ
U0w/fCwN7b0EcTar2N6a8L5GeQapJYJ3qdU7EM26b97Aj/Khls7TMIOgVbJxvym5z+WWvdzkgTu/
Ob+RLJd44szZ3qpAx56BWaxfNXycbnoWvmVF4NU7rwGnmf/p0MHDlm+qOqXzNLgJGfCk2lPE01yV
eC6yz0PMzCQzZ+fB8DvCc3accr/mhBqu1QDoI3NtewmOhvo0wXT0MdrcQYCBRi5uFg2fz28svZGu
me+fWT8KEhLNnzIgIizcnYsUlLGjCbsxxQwLRZLs2nKJdoMXmi4On2PEpX3i/ixvehDFDfc4Js51
RfPnQcUGNnT2bZmBCvLJ/Xq0ZDvOvhegiIhqlf+sz87EnNJ1b4WeF611VnNlbCljn4tANvJVmgER
bvXGwjcIyuBaw3ejE7hiCSPehkRH3JT3ci9BgEPE1y24cNAF749ohK5cmBawFReJQG28LIE2qTI0
Swv1dhdm9GajQVfa+Kq5iqG106nzY314384wJ8t1QUnrTVARWvQ+zwQ3jv7exrQogARU/BF7uTLD
Twhfm3s9rrCxqqptfnilIqGAib9uML7btWwsTClIU261bJvpRYxva5LkzV2YrTOZfZFu/ZwcPfpZ
tOfvmSxE9aQFtzDjkDRqE3wwCEQ+dTyG3cC3N8E3hYf5FNILjN6auvKYVu8kQ8AHpwbj9bvcVMeN
Y4R0J/07+7bBKXWv8ExFdmDUWtwAE8JncKiJYPnCLtpKs2YSC48B5tbBvcBgvhIJjPc+F+DFNj4T
JS7oj1sdfpBUvP+t7S0iM8pcpKcAYi9aYwQ7hXak9jfmE3UbAb8ZBUhbjBSRItjF+rI5SBbmKSbw
a6ALWffFC79r33XmDHVQ/v5Vek5bWfqlHJagptVDKDqb4/9DJhpAe5Po2pM50HyoGTfuH/eUBfSD
o9CtgRMqXCpHbd1gaWcxxKNdw4ZmXcIBxYSL8/UUdC/bxN9xfAd5oRmTs95W9533CthyZh2YaYqF
i/AErsHxDG0nUGIZ8OUAsiUIPojcVzCzSHor6ef8SHfbO3Dfncs3XbGLnxQAVCuQJH7UeAIId7UN
TPWHMS/fh0WA2JY/5ZPoybx3wMvZbrsIRb0rVYHigTQ121YXb5cthqNInfJDHUc8Gu4TyTrKq/oC
YzF4WcDpe6zy4/NtSTBW4VMVN1veujuFIv1ixYa2FBrCIhzwC83klsAl720pCJ1v5GjVdi0pvcx5
eVjcTUOR63vcVKK+CBGwWtsSyqd8YZsz/KM16G1FvbkL+LGUGFSACmnrIPF65YISrXtlm9ZfHDPk
mdHxAES4DDIawx/KuQ798lPDBLGivFubeaed2+8lEnwq4woK6atuAk2qqFJ//caGoFVHmmsK4ggg
hbR7PBl/RFc4OP4exP18/i1e4QKDy55GwDpU2TNhQ6aFUTX2MIsYDVwTrCCOKe2U1pxZNnHpYEcL
lnC3QNMenzW6GlInMfHQx0SevLKvK7UwoyHOn2AVwb3RxrtonciXyNetrl7XhPh4RDI6i8qPx4S1
W+kRFOKPv3Wo7FLnf1F6MSc7fyyNAfL8qhBNPCamb0kr7muL8k5yAtvVngg6svrJSZ8HiTfntFzw
sqBeVfvCwo+TjmC8GKcvj3IUOBfAntZ3hNoqg1ag8rhtfTjmcs67c3VBbX5F/tEoXTCA0mAi38Xu
EEFDagcAQRnuWu7I4e5l8E7TwjC8j6iExqJBd9vHxdYRwwO2wLOc9A1XHgaE6n2HAUUVdwNFwDwU
UXCCSMlQSG501GVtlxfFKU/K7JIuydFKH/UDi9BrJvmQhuAsdZ88t1UZexeWzfWzmCZbf46onXAb
cjCSW/v8hH8vHnZkKEWDCTY5Zoi2dChyudTZptnZHfUObczPscW0ZQvuPQigG83KK4Z87UA5kKHY
fAh8+JVBdkJa+a0MaGZvGaSydZGfuRZ4e8Zi4y3cTEjvC3EB5wAs4EdSY5cxYGEL1MD8lKC3qfPH
ENEvm7SyZuvzuneICE7YECZ4YHdvfIRQWouuGJbWErcKkPo6QLngFyerF83z4vqDhjDi3HGt71ie
12oXvMPlzz0jh4z1QW3KBwQ37iPi+sOgsBXHgrBIE6c5FZij/adIxmmPFsdZC7ZZOhmzmyOf0brC
7qtE8gEeydfjmiv0/Clp/E8jMXXJCUWI/4cOY3i8JoT9V6QbTfHWXj/eKILdZGat6c+PvpM1PepY
iR5QKplpnqgfDJFyR29oiTwYpvuH+K15/DF7SiomzA2Ln0ZPexPhj4EqcfHK1OkMTf2XXeSqJF12
AuRwFX2Ke2AfO1M2P0JDY0gVB2m67h2h5sUKbrA8lQ7OSL/GYWQDCTGo+PDl4OxFgcWJZuI5Cyq4
nZuk/RASuqKL4EfYhb79cJSIVvnnXiAbyRwtPSbdDX7XkywrvWxwjhFy9/0FsAHfd8oGt8mXcmn0
PHXYfjcnpXC8Plo09XmJEWP7iLLCk/Rr/E/S3B1xLTpRsHPfZXe+R9ZeBBI30uZASowbvgJ1FfpG
wLoW6h3R5s53Je86/+o0Xh20pN4rDHT40n0/d7FY1ZAuR0dmSSVlGX+OG8TxqOT+NsNj1npf/rJy
Cfncz/uA/Lv048IuKECwZWOSwDwyK+HWA3iJQjDrQ19fCDFso/K/zBdBSWUaqpH9Qpk2lPUwyFlU
YXjmsooIYLGckIJR0UE53bfIUqx+NFo8q2fYgkuDXZUIMCjfu4jRNMl6O3abAPABGh45lw94paVI
NLJZ4zQYYAvj3gEB9ILZbeOTRGY/GHCx//OhFAwuydvou6Zgc7qDbeapGSpZwpQHFGxRrDZRqKyp
TL0O0Pghg/mPVwfNT/dSuT6VHeHxzF0wcfNIvIl0qt6aaQPZIysjYd53cmQR9FeODI7Fjfvkr1Rd
V0a2Th0hoI9Ya2Zd2nD9TiQtDQ4UGwXp2r0+mrhpbzW0p6a0+uBP2XXcQOE+X6qaWPwml25N6Maw
Bs7APX5z/H/nv0FDuUK8xNYZcAy4cZTLypEEReyaLhl5jx62OQWg/No1GCJtYaX2V0D2c5YVGlA/
6UVMhZapqWhOA/ByST9q0FxTIVDUPzupcFw5hppqzCbI6Jop2oPyvV++FVcb7cQuMOioGitIwbn5
eZztrmRm7756YFUE/ddopbhjcJz8X+73NzywxMMinP5S0f2B4kKZlFUqRejyom02pSenwU/d6VVn
LLjzIpOTWewHetQMPgY9L2pdrVrc9hSOX1BQh/G5OdrKT1TTaKpVrWXOTa9HhKAYpAghEKMHI+/i
DcDCVjCqtPXdEebMKlNKGdgh7fNLrTcYYx1el3vs+Bi0O8kb1YezAAvWmNYXOCUW1JmhH2/zdtcn
FMFctcOYMHbPmb+xaGEKKgrryo45BeTPqlRlV3JqUPh3gebbyeRZlWBUb3rXQOfXPhN4sPTkfDki
a0ZlpDZNGgctQpHjwISQtP5pTtvmI6/H7+lNfVWAvchQuej72irZLaYu7C1XKZn8QKuff/lzuiIT
o8tIUntppRyk0ZisILjwK5Opgo+bCOv6MLN3iMvHUZ5WdkP4aAI7WsIMqPajKOF7U+boe48vODaj
pY6FIzQ8DREqQOUvD2erRhuTB8LAz2LI7YUAnZsL3R23/rYWej3lnkrFkzLcBJaRVmWwIhHrJa5S
BjcyDxvDrNoN1RZbUbVKD0WNmiJGijIWrZFUySMiaNIBjgUWAxeT3O/Di22HUI/T7DF6YtacYvG5
E9jjiuK3pATpNpFszx+Jwe02s8ZrE2cS4QTAgzWqHtH+wuJOwm6lGIyp1dx3BDS3/5ML4S3NUW4o
ypdInoiFNZjqhityc4gAU3mt/WNfA44Z1l6cZfE6ck34gWe2ZhdwpOcFySEys8eOfMHKVWv0Tvlv
iCxk3m6IksapNWcjLw5Wy2F78+QlQatmgGv5WmsT4HpNsINjSdf9eaK3bTJr4oHzBftgYEJDN4GU
kAQSsUKPvaYXXKFmiRjL7x0DZkMoDa6nb0T9I3VCd6OKdVaEg4G26iDSGPcTl8ApTLuJQ5X4IYgG
NJhX+ZUPmOIwM9fhzNxQRocvP/uYNqKGJo8bYMOonuAx7dNelUq8JnCL8rR0k7bOYtP4qJ1U8XcY
NZe0wozSPb4N+uIny/Rr6AQTfzChOgVrrrGHF62HLSZPYqiOp8J3yhLCi8vES2CXm34cI3zXRRuf
ISUcXoRUCI5BsvhT4+iyvC3x9mUyGSbZebq/szuKIpJGMv8KyXPWEw+mErRN1VUcZUDwz/Vob/VI
D3IHJTDsJ5xnJ9UMJhxamH1qb9ZRW6F/nJckDCpLj+vTIMohkkKpdZPVa7H2d2bH4sxQbY6ub79D
kyHyKVewn5IRpnY/b1Wo5cic3Bd+20QZwZFdw0Umks/gxEX3HgfM1xSAxw8u+3y3PW8jIuytnINg
xpKGvyCugADPz3fPZ+4Ctwaj47sA1vlmdIsk4tcVhukRO9CzFr18crKxEBLKtIRMOXzJhIMvBerA
5HDtQpRAqlS0A3NhOb//wYmj36LvFbiM+NCcGO5v78aZ+0yOL3/DMbOZa5i4U9OKvjMIIVx1ch4r
oKur9+HAKralh/0RbfI5mBHIIoO/VLYt0OKoYOoAo8Eazjro1lDTcPXFar7mWLMjAHbieLmGYNqk
aCX3o/tvA6g1tS+mm24Yx3TuTQ8a4lEIkTHMNjeEyonwbbJ88gZpfh60UcBSdFVMlMd2Pojo9tN2
aUGWKcQ9wk9kQXa+E9++xq02cZfVjvin3MZ9Lnjv54+jcMFCpt0yqQVgXDuQr9JlhZN7VSeLc/wN
c9rPC0bvzG7lUAAaKolsnYg5oGTPv1ob8jYZrIU0w3c14L+ef2lmF+EL7NZdV7woi90Yc6BadnqC
t5dSe9yq4jYKlKDaC9mI1WI5wEeDExRCBPyTOZJ608Jq9HKRaEfHVdgdklFFSjEhj4dBGF/9TU7q
m/NN+ZV+k2MPCman/OX588Tic62sKtGzLBZ7cLzt1Wkrni+5ZidoyxLpKbReftrdq+ME2APg8Iw3
zleDU834O+3qDxPwxyrec6YaQmZCwQZTUdFsx5IwoASxrvJKuIJPpPOm7GimyGbw1zkOjiVZ4F5K
TYRfVnm2TGZj6q6Y2ndR4klGP32w2bziP2vsPcAIB0+40v95m/bbfWrzyLKq1uKN+2jThfJdyVIc
aNrWI/Wy/tdJvqID9WbyscGGFIaUYfO5FWU18cJXzy+LoT3M5xTf+YBb2ZmBcOR5ySisgMnUt6e0
PpI5KbhfMmdJjQqecNtMkGyZIHUcWgnCy8G/L82TZjt8J+DL+Z1R0m+oJZDwMsvaycx8xcyE03hO
FyajWxpXmeuf/UaZW5gJCZ5C1Lu9nNz4pxY6d3J9Qb509ZATyjeIAdpqPLSYCHQvQMi7pCgyrpnF
2LabmOnvaHbFstID4iticKlkA2Ucow89/HxLaRuWC+l/+tq39kpNtjuRYbuyR7/XvGtEgHiZJFwT
QAYyLCGHt6n9wgx3Rpl9mB/rzyW2YwgwAtJxAnQdBbnyRHn01EUp7LSfO6p+0t+oNJ+YIx5mz/pH
CYrfRt92JirgF4MHJu2PwAy94CFv36qYWi9pYpEklivkGYNJZh914sbnNgov3y5IIvgPIqMVr+0J
lWfrCVktuH951eiVqaqj/DQrQg2gXafX57rcRHU8Y4bDolmtr2DucIG+MD5tOqhG79HE2UqZSz7R
dnLyRiyI7OjMARgMJsZlj07SzhY+Ny5k8CeTwLhkbc4d4X+n0f96/eGWJ3Ydjh+/9Yby1asZJlI1
8IQSAHkmR3Th5XGYj1aiEtF5T4knH2bCEbkUipujR3gmSJ75RT5RR++eZ1NRIeJPqDv7eusDoZsj
9E4ETGxMQqzi3OASM5bXfm4OmKyx7fTHFRIJ1XGpRkBxS+/+XEkiTUhtFqy7I4HF75B0WBnjRlrz
o1QNa8543yxsJ6gzz2KTMHimg6V0EyiM6Jt2qsF/xmh0UVaW0CHEV6euI9zkJIFDZISAcnOQvG2g
bzRLzktKI6fCml/tBUB1BufWH6WlWXm0XmwOZ3byJGMQyuAnkPJ8adkHIcKlbjWgCDEVfi+0livN
Y7SRwyWoHpxqZ9d7TLwR40uv3q2JxTBrI8r/6RTVR+P6wtB59wyiJ0W4iPGrG/m0wHcLuWdypC3h
+IAnrl8UwC+A/KxKrkOpkHHFRmWsvVKuv57IMuk79be6FQomp5k1iZoNXGtzQWIAX/7kGpziPylH
2qV9u7QfPPma1GThW7tMiilXhcZOGJNho+qiUsS74kuvtC2v1lYLbDCF12gUK9QvGWpt5WqWWQo3
Qz6yXPcnKxx3JMxmQuXdNOfMWrE2mwSgGmkolAFUDP33ZGkIwBYcmQpe9ssLZIQeGryy0SUGT+q7
XwAXoD+4QPulQEE3tsZ8ext3QDD+1pmUpZFPvdLm3fB0iZvh7eoAzX2mXma0q6pAvlY3+WYIou/8
sOBHnqgwBxtKc8F7ms4feBwRKhkRrdWpNRUyTVerjB6eN389YcidzjtEkYcPe/yHjwCnoOP9djKC
0Xt1JOZUspF1pnKF8Co9YLf+CILjr4Ol9NOD+5ObbCHpDnWkOtbsfG6NSlFxaVf/u0APLTi3ljmQ
bC/n+tYYeMrx+gERJ3Qgv2OuULJwqdowHF668IOX3o0MQOLovqk8gMXEqvpr96hVQybaygXl5JJf
XKbtVArnO3mvT6jYOrVVtbNX5dKPnwe5lQIHhpULH64iU0gGCEQUcNGXLyomTsBx3rVtB+FkRWx9
HE5rFyy6LnUtevqSIiO3HMKkRSvVsDurvx7azJ7RJHI+xB5GCQgpMISyUhcIBptb7e/rklmnqNmi
5VI6NHzvetouNZcH3YV3AvAgbuS7PLbDiLco5+9fZB82NWMCUZD9J44zUoFMm8ianOsuDMLxXMON
w8Kk0JY8l/WYTLD3FHreWYfA6hwCZqXHkySqmMa+KyQnj0I6nrhgFIlpIJo4UMEqIbFiw0w8zrlA
oNsJ9YmDSCIxJ8EgXSYWz0aYJe5BKB7i3TjVjh8YD0gpSiQZ1EU7SUglpNDvOndRs9u4aFLNFfoE
21AEb2CqrP4Sj0ZlepAnZfVrcznyqIHYJw+6iq8dzuZUnu6PFxV875vMLkc+fJYV+aHW2VjjGlKI
iOWzzDqI4f2ptuhq1xLDmGMOrUFXoaSgOGoCRh9U2ednxF8LTqrrueAcvZ3a9riJetAdFRONyHz0
x8aaSP9cWYED/SQqzEDntUmpfkdMED6Tr6nj4t3ynvE3y06T5G8aeRuU+DAp1W9lLgdFeNxZGQS5
zbUgkO2g/1WyZMuVL/rfjLXmY6pxBX9ymUTDdRZ7bx6Sxfl2S1NwuRSepX6+8pIfxQOVgrULx/3b
Pidv60dHrUKp35MVsFm5rvxqnGj34Qop1dIXulf0TPNIhhGI4VRwM9s4PK4t+F5e4ntWjHvFLLE2
tUdTnq0artzrqSWOTlt41LXn9U78eXdr1HnmGooEsFORxiYmvBvRLeynSr+/As45Qnj5rp5cWuCr
pVX/+s1Ema6BVuXq1xvZYROlQSu/1ZP/xX6QazPdG28jE+SSWzYZZ+vYMp8mLZXg6ovttbEkwSgL
Y9W+RY0hwy9fvZrxyMD3AAft69hphqGXRs/rrPCJ57Dbq5YQ97sCHQPkPLS70nRx/DFDTrbQeHq4
z3+LBl6XRXm0vp6ctxG+AhRLKZySTS1b1r1EMkZwxiviwcReQRsUqmiZtyo+CTe3KEMKIEebV0xY
WKyo8USb3D+zBQl7dM4cSt4txdR3S4oFao3AKr22va9a1aduDyP+f89xDeElFV5SQzTwQoiUMsiE
E1Vqc6BFo9mSXawcD2Xj86D/KIEP3YAQ7tUp1fVUko/s29djb74zVItZo8QJX26HtLqEtdFxMBHQ
YfesBosZ1jo4/ztZ6eE4tLDYgGwC/m9P+mISLZLqf9IPlZDdKiQPENFZv7cDGehfwKei7drEXvt8
Gq9A5/fsTvRhuvFyWxGhH7fjIBmLqtxhsLfsVizwDEjfwRtwaB2QbUevtfw7NRBDuiQlBvglvE73
U3qdxP2aT4ohXgjmmdU3P+q2Dgq5EFEvgRWKCvMUYYKbcuUstAT40xSzTjQWC3OpbO6PHlIWhqVk
JTdRJqsugXWzgO3J2tdyBYc8Q5niJw7FZF57T6NXlW3GiPU5VpB+ShBzaL+hc+4SIzaX9kTPaGlf
gf4ynPQrA0Id0+4eGrlLIOm5Efmzn606ps1b9dI4rCsJ4WxJyYlQ6WCnFYKp4oXo27PNF2itJtlP
oiq/4ne8siMq0Wf2Li3+S5UQGz+BQllxuSMzAJtSlRC9LIPG6lK5i5Akapm+qQ3SGOQZU0gFIMz+
wX6pHH6Y1EihcUIkJd7H5l4KKlyaNPWC4p3FZkHKerpOFqD+Z001gzsvf5SeiRuwklG0rhYvMNZA
tHp9+jlU8DjKdPSYBJ0cSyazsdll9mxAxs62ioNCljtlZv8dGA1zOdrH0uPtRS4/0Iop8MWStj3a
kTC7WrZ/Q7g4N0nGNujwvF0Qvaso4b8jIAol7g/zGzYV6mc30hJggbB6M8xx8kQ7TdEd5yI0iPfo
Ln9RLhozsa5JUhK8epbkiRvpXXzXTlyZlcLAldzhGGDDsyMyqNufpgBl0hfpw/OYDjN+FOArHsp2
ZwPh+fcBtVdUvhmPT9KhGHlyr/4PRq7B4BZyaExPDD0tEbeM0K0G4CHSRZm7w3dSdKo1pMnn5uCu
TKWahx0WsqlZK3oA6sCNti9use6pWcEAZpnWmSnT2PSxmupvggB8oLvJk12DCwxYdNzRuC1J4tnN
DLOF6aPHtyHFKCA4KcY1o4HRafkPHnuyPnHASr4SYIjHl+UddtrlI0EWuWmdUswFeKpDc1BBlq6W
/j0BbZAqzDt7aj+TZCKzzjfo9ZpAyGQatH/vKk+fJO+sgjSNU6xW202QUz+cIPEOm6zoYSibTiFe
px3+02d+2lq/mrQmzubYMfvbTBUbM1CwhtcOMiFvzy1pAZu7pyjB4uwLBZ8Hm9yGVezlckKb6YoO
yvmPJV2b/umffeA558NuszOf8Acp75qqxFIVvH9jBDZhZwQ2bYaU6TZLfRlwHesr/1EANQwi61uR
hH8gR2jZdcnyTEKyJE3QM0diEimb5u9vQ+yqzS/nHXpo7zll6A3aADwQA9mvx8G8rSLANFJk3Gzw
sTt3ux7EzTTXwAhyFgezjPwBGzRk4UdoNtjOH61l5V3rJEX50jZL5pbZAOfKq2OEKFEZmYbJ4Rw0
lYX27rfrgxOiLpalcV2N9aJeEvQh1teFV6932Xy3dbM4Et0K8ZjwopHxLZzeiBj+Od4xpeuXGCoH
f8+r7HOQqkhvsnoWDLPXL/h5kEYlN1XCmlxKKFq5sXYhPwCN2DFPIC8Yo/nZseOg6k6WhxsNMiTa
LsMw8wcBPBVAsv2PcGrsOxDG4aJwo0d1kQPwbyaRmmjthElcSYUNjJ38xZZSCimxaKb5TqSE1jXa
z5bf/rnt7oLwhVuZ6QLcw3do0WdT4BAt3YIjT6lxCxxrsSbDtgSWRvOGiUVPacRwBmiulQhKAcUD
S7NJoiiUr5tAIeuRw9LGt017f97QMe4KZN/6xUPIuT3BGIVEyVDRCog5kMmnmDQof4QF3VjOdnWn
VBq9CTDvNqNIj6/4U0GCcb5C05WcERHBUQfzdlo6SCCR3P/bpJBfc4LQTxmd4IJNbIsAWmEvnQXz
zmCv/QOuItJXb5JBx0O0T/nrb/WUhvXoVRcTeAJSuuDBIWS6rWmM2kEePInY3Y/BNtuGGTfZIoNm
IHsh2R9VqnUrJioLZd0HKS2xsqCDdhNTR7MaJ3ra/NywHbl7A5gMcoP+/14U9xNPLzUm81qncnbw
XM6ASIH187wnNjM5RQ9CvGL1YFfyhuRRaAHPoX+t41Fia9IW+wP4sgo87+WEl/5MPS7JDjrBVZMg
VLZiM+EdtI6zrHWsOJZpd2HtfRhJnhrjITSDldw2qs0usctGTEp4RHbzWONLSDmTDkTaOUsspHqX
zX6Uvxeq/7rh28TL7E9TBFNR9VgivXVje7QhMamDGuKhBM0U06uc7fn7UlBKTm+zYIiYnVW90A7p
UQeHV8sbM+wK6TIvGJ+6KBbFOZRPDKYHJ84cl5SO042Fs1rrtUC9dwC6cact5ClnEyHRohGr9UN/
hW8G5yhjjAhi6EO3IGOFltm5MR6inuLBqT5gwuITvTpkbHgeia+9ME0mIyRlhQERL8jimirvGK4Z
TShdocs13lM62HA3iEr+T9lG93KFbyj7Dh/iSjJtL6L5tOsBsOuwXmN3ayZIQAy1w4QuBfyanLTy
fxyYWummD4HTuEllfeVzJNnS2bA+pgLerNyIfTExzrzG3Kh34dRzefc0j7Hf6/8W+wM1ASDQu/Fp
tXhlYroPg+Qu75Mrw+sJ4PEOiS87U73Y8h6CRKNauMwSxmMObb8hDOEz8AwQ/3RRzkz4fLwH1gnV
R39G9IySXKSguCoNjtOIrHkKEFvJMOyW6Ml6Z9oehy27ceMmfHt8T4SDxF4acw3ptB3XjjimUu1n
GkBRCvIq5va07nHh6M+YKbkxMj1+toYqt1f1vBP2/e8ST7bnd3bv1JNYtg4qFGIfDWGt8F717Ja0
NnpKkuN2qaVIwL//BtRzr0WOgHVP29LZacHB7YuJBSCI6oo2EMou+uRNeo6rIxG+h+QoKwa53acb
fpdF86JLZ60D60EAlZbupkPqUwUgfPr2jcifydIperpNwtWAtT7eXErw9U3DsQU0Csv5jMYnG18D
wb6Bj8FWGiiM4er/XtvbljG4DZQIgNxzCdZy6z3z100tEEGe6u+rtzUrQcmMFKaKz3j6f7oPTqjS
F3ioyZcHJphDa3nP78qEnm2aBV+BU4v9n6RNBHKWo+MJKOZebIe6z1yNYZjEvkkQeh2vSISV3Dy4
4z7F90aO4HYneU3a260DJAOtiTFfmlsJSwCxhBVzMMfoRzHwhAs6Wg+joK9FQKdAdvQUgp1lViMu
A5+P21MgT46kOKXfDq3/yMQkTdFCOLxdcWygPnTYqIthRsrQYXOY63eXauPL98FpUKdbdSD2P0MT
9cec8y820Y9+aM6KZfWdnzt1TfCtvpyv6vJx/YDGIjKlu53Ix7ev1aeZm86p2ruhRg9AJFdf4rVY
xx5Ob/om4g4ZpPsUmD2BS/rxu1XFbq4j6sTKW49vrzwVRdbsmDJtvwBFQ+DdQWD8XcyKXetZd3T/
XHn3cEyyW188yXsVsEkdNI9AFgya3n5qohJiQvGsvvS9/QtkPVh33a8R5KUQq24zQh3Ru/EETlw8
R+ZLqnmlAG6YWK/OBCEkDxW+Iwo0XBukQ/dsMQqmL7hsu0HXe9N71Ri0iBFtEs9R6iVLCTCEBJOc
lVWd5Pvu+po8m63D2V/wIFNrhC/mwiKkh0m73zGh5xBDHaSH1OaFOaJ8sW2Oi3mbPbaL56HIr0o6
CluJv0XUP3mOnNYhjM6OZA3LYqXFyh4eAYAdolJMRimXAA/I4kI2eEEJNSm3pzU3ywr5DUcFnKGj
sIceroMgDFotOkjinoGhG93PEUmo/pAlSEniHmsoDFBFD7ok/vCLPMYWgDXcymx6/BUosqGTb1rU
CWbD4688XbK0QZZU44YH5LftqHpnM1yJ0YmPKQEfZNh4zH0aPdEKwnzbR2RGo5nIJPxmURH2sn8O
Q2mPnoMFzbqGS4Yt0O55Luoq2/QCUnsVN0AaObGd1dI0xi9tATj2e2XgosskqSFACDt+k8iN3+Ka
fwuN1UCiar0hgHN3ct0QgSVvpDcMs98N3t03ABGIU5jd2zQMokwvcEmP/gyjs0nLh/seuu47KKUA
7moKoo1snNzt3H8AUI1l8VJbAkoqijqdxMdRhMxIYke0L/oEgScRenE2HU/s9CLHNv0KnIOzYL5w
5ckQdugcf+4FzCPf/FTOmOepwC8/cGnn5HtbVqsMT54sW2NRla+YaPGHQE2+AbdcRo1Zm23Sn2gl
N5fY5lK898oHHTbIgAnTyc5AS0olDY+vjR4ALuLt1Suc/rYuc7eTO9UroecSvsZKkiaVDKk4PByS
aRgAVGtFmScBCNNTFZXHIWhTMZ1QVriaJv1VmI1FbW4i3xMjzgofWg/Nvw/I2lj/fq5hjjnc1ICb
V+kg+CcmYsu1LLk9HFPVqh6//lnUeP6LNfzH04vFjGXR9ywqwUjuX5DzZ5skHmpE81SArzlgk/re
PdXqZk+ZxYgHwEElL8GGAPaGjJMwES9HlMV3v83Nv0sRXxFV6q9n6Pt6ORKEuWGB6sglFQgpgZq+
XlDSBOo/38LrcoPkmuTX5AAuFzgsrzlx/23rxxuqs0MjZGqIkUVNqFOC6YLuYUS4NIczCioSU8vO
vQmpOhAZH4H6X3imTE6HJhjfbxKedbco7dpd3W5QHHnc2uTXzNaJ+8zj4G1Oiu0rV+bWX4jvLn61
ZUMzZ4WsRwDjdQahhZfY7NPmltdnEQGk9EF/45glFiLBHE+TPkkgIz+xk10Fbnt+GukR5P7XHSWu
O6wImkSdGiT6NRnQDf1U/ln90xB5WUqH3xHc7vBysMhMenBNMY+enWSaaSOfL+9HUYC2ZAm8LUFx
7/230dKCer5i4tLalamtYbHOq2efZlRRwI+ZArhi8tgbBn3Ebf4Ouw0PFe0OBW0axj2e/zItv5dW
s9o4/4ryFbEsnprV/D/e4JChb/Yig/DDatLVoNrG/4VshtgXTvwZl9JlM4Tl+LQdx3Pi1HuCFAg8
Q2umQqbxFKzCJn4ZbnEUxpWkSzEGv9yOZIf1vy2vIUv6oeFZ6NInplB62mUZCn/x84bECWfnnCfl
BH4fxs1xLWFMhtPr8RlAckWAMPuYwRVfVaTDMIsCrsFNf8K6n0Mt8rxGQJri3ZC+FBhwBMyYxfk6
ZofowpK2iG0kYwopAIcUiUFtfWc35WqJIuYcGcbQGenKJ7ySLU9uMspKNYghmaq1dcSbtUlA/gVx
AV8qhLvdRicfeGcRJuAJyqc2OtDgL4cE2kifpd2Y7UjvTmZwfVh2JLEMevCBna6JhhPYUC9UB3aI
U+hG2rabuqdxpNshY0ZSdCrVOUBoOm2zklVHPJE5Ps2lb2I0XSGu3ZyEsoVDMfsk4nWDi4fEMeKb
D5IeM8JkmJ3iU/BGcmQrToQr+9JRJT0mo6q8OTy7CEHyP2U8XJxcMgMiVrugpmGYjDugZgtRPegO
H5UFtCbRokNrOt29sgYB9NXULrvrGisM1ELNa9WASG5cS7Sx2bClsWZ5nEz0hKn5Qtf9GAI8a96a
/Fkk1WZrG31bv90JwC4BHi2ZvUQJnN1QNRDJfiuctCWblUUHlTk8qOxUgrSPV3oT1IDPwIqznsKa
bRUH1MLaAU/wR7LL11RL24WqEAI+WA2bEmreuo/jSTe8iW58mbLJexNiiBICtmP/3FCNAwIzTexc
CkVi4fNUyQhWTb7R3r3iX01qWz2stm9P0dyrbERNGSo3dwDZF5F8MmV23eD6h2f6EXP2G3UmYnr1
FeeSgEPqf9bKuY6kuWQ9gQdu14s6toEHOlEr6PUa+1JPV8I25lGbcqqHUrBme3wMBa1RXrdE52yK
U4epHps5+UYqrNcYzabGgeo8VmE4ckOyRY5WB9PKD2S1kOQOUFKjgxvSwz1Uw4bf1bkCkSBJr/d+
G5n0QE4oYb1dKDZsLCpmeiVYkDpa3EfG+cRTpBYeQGSc4+WCcHPG3OXrg+Xsw79x2WhXUv+cn98f
2872b0IBNpmEkOne8rCwy57Sa9sQhGX5YLYidsuK+bRt65H5XN8cv1dEX5KnBImN8O6Knob0a93B
+4yO1CacPhIG0HHgOuI0Y9wMt2SbaYE5AM9+CAV1QY2TSAg5yeAdf9Iq03htNZm7ndGnwPuoxZp1
prY11QcO78HBOqpC5aGJ9vjgoiHf/BEXUQmM31c5mgbTIWg/L0Y6TW+n7xFCWHz55C9xgsvmsZuS
MMgaALlJ5bz3q61XUyNRBxa+yUrXjeZBeqQJYJhXvyRRh2QRUpxd7sZZUz1uEyXf/CNDXSknaffY
2l/UFTQ2JL1SuYcVXEJ8c2p5fRxoBKmqrIBZpFBNx5KkaLIqFtNcPTbhD/GguwIw4TFnQvrTTfKr
SJP4sz6lYBDTxvF653Nx6MOlSeblQv7+WI9lwj3blCn4cDGGKUK/5lP9741EWDRTAJ1VmP0ameFa
5xnZ7idjHC1pd1onexMH2k2D2HIJkMYbSaIm310PnYidrzCRe9FgZay5D+WlDzAz5nDyJhI5S7vL
K7E04Z/th3INPn7TkiDhixRl+5Xo3T+biq4xnCpn7/J1V3UaSw5uyfSjKtB9mfT9py+VVWGWt8J7
Lx3Nd9A1nvaQ6uPGqSwnYRKuTkxMC5ukGrEwp49rQu9KzTA9OAa7ZyMGXU1IRuV5Qm/fwCEu+kZC
hs+a8TeQX7WypUoDb5TbeQ0/gJsS76/7LaQa0K2EAE0Yq2TBeQL8h3ZJ0iP/mp/2VvHo/+BM6Pny
KHwu9mPJtTlH32ZEG6+y8loD+Gtn/jsFQjy3m5pMFQtNzCaq5Ly07UcLOaKuBuKAsBrr62kkNB3s
q/h5w7ebOfE5p2PK0HaDzKBUrga2WqdZOXZjZiOX8tsOoOVoWfUjTC2CXZa0wUNE9t3DP3wIjYvg
lVGPbidj7Irao0vVHjZRz2xuKPcul4+asAuj5U+AlnX1ZnSam8mXpR2W9vGMS9U9JQfbqD+AESUC
d+9H5LzOgCQ77VzmL3+kpMs3uv2KUU4dnsG/G16SVM0tctOg0AAb4Uc4+mx2d0w/HRuGabTg0qa+
p0cFdrcEvLtGxy/9A/iGv8opMKe7mZJO5wtJme0TTKH5H5FbMupu5f1nEQsZU7u5+w+rkqdKf7hR
ktR2BaR8xP1qkdWdx7GryjRIzKuR4E6dbDRkqC2y+bZ/aIw2cSJQPCfQhykbmkJYsGP5GG/bO52Y
v0dEeHKYoKVMqX+1Q9AwTU8898849o+NVOxrTkrejTPSBddrfmMxZSkccS8Ca5G4WLFzgqJ39W5e
vnmOpTWd1FCyFV/giXoeWyQAjZtpZ+7ogpNohiM+D70XmkE9+4R/qL8ugE3lqIiR8pzgxo3+UqAo
5Skf4zy3Yi7rpCJI8YwhtVvPDJRCYdnCA5WZhaM/V2ALiMOeL8mnptr3oQFzz75TyUwehk8b7HAY
NfbQVDccvtUvnunyHw3V+ajM3PgPy2eCRzA3Bnho5baH7LBhl8p6n1Fbed+EG21yPoWe0gdNt5ln
HwYtLImwfoahl8CimN1d8gfPlm2v9DDSiDLG2JIJdmdIKrmomZwHdv6yOVi2cJSVl2QIiR5OgL63
9Q07UYHvbQcPbbkCgu+pMjOyMZkrju86aIdvxSPuGF7fXhKUcrn8BK33JRMa3XIBd4XAS8gLqF9y
7bQqxqcsvqVTX33Yi7a1yuMJuOOzN0+g2An6RRNCQbxKmNrFO44Vj7ZqDM2XXd3Z3B84QmUKreLK
36HOp3GLEvonh2+XbPHkIvOnO4XunXubvdyJ2K5/SVPn6e/89qLKWxyuWLLgG1y6kVo5xPFBft4Y
y+Q0IPWYfMSR7iJsWIg1ecpkqHSvGAvnGCE1kh6ejDt78I9HC6kQ957jiNdlMh1Iaj2YcfXJDDrB
/mx9tV4RmPrvExOj/7RGb9+qHyeNpoF+9NvJj/q/51X7Hrcupyjpi/Phful6U35Ydbv4NDbEvE3B
QpMLg8K/H0aKKRBg69dp0VTubnLurfRwXG8YdvMYfl3ETLVCSQJDqwoxSsH35oD4JMLRcrtWgFIC
dVkbApGmxG0HfEhrNc3qfycE1e4sjeWkiWCZ7oW/nPbspIu6SlZUOAwSQgOCRC0wf8t0UYosLolH
d3m7xduUJytCHJZ64zQq4e8DLLGQHMuTvp15JMFpzjDd++VBg7GW8KV1i2T7/2UoKaSCAXCf/ax9
shYeV6bXU1SuWO8k4x0t/ioRv8MKOPpzMIjSHuoS3uHNrMuKR2U6jFMUGqafJLciixbIRtI7bEas
lhTC0nWNa1iNsxauJJsn5f7ehp0f3jwGQxEt0VoyYqI+1goMkxzSENFbotuZp4A0uVkIwg+FWbCn
JSRuwu6jtRJl/OXsyTn59ZwSwGLlTvpdu2DGxpRe3YRTi+c1CwEwgsppaZcZkCy5dSJhZW97p/KR
v//R+v569NORTUC1M/widRzZYHIo/rLoaLBD8cguedIYXKEDNO8Wa0jqvQ/eXY1sUnefbCM5UXhI
YcugTorvd2Tzy4HOToQXn3blsA3Qg49JC3F1OxHliAfLVf6scoWYPCTy0UFVa5/COwg3fk7/HRK7
qdVilOvxLa88u9RCZ2kHwSRVgyGH4mb3fQ9TOvoySv10xbs3GpMwmBK06U69FeLUXlhQENQSL3Tu
/suJWLhw22yPOEg7qlYmfaMft/q3SgrGw3wKVG6lfVR6L9bFXqUnFxGezVHHilzoNrMo607bjVgk
ApwIe8KkrAyDShcQo6MZL1ISTRDWwr7Ftqm3Qei69LhUjWnMXpWUKtcNveK2t3NqEPd6ljDkZ3PW
KChPhodpNB0N8zQBeQ8Fr0x4q7O6zzR2RZsTOuAx207/Xco+nmhQ0EfES43xbWV8w37AMAlVCrnM
IZhGmOqbekzrv+AC+LfPcnuvmyMenr/JopJ9CAyYb9YJOlwiOPuSa2EPksZvEj0v7KcotTJEfwG4
pksEc2/w0QkxO69z+jSoDnOrLYFu+IPWUqWVASB6ff9jXwMxsP3sz8Mr1R/5Q4fBkxzHh+b9/gzD
nHnzOhHAAtI7+QBUKQyePi6uVWyJC6FQMb6dgP6DO/LrYe9F389ZAyVc1JCijBEEDlUf7JFBUKZ2
QVtS6ZW9RYGo7MjAIy6bbwcCnY8xt/VN/Ps4+fAAMFFk+Cb9BVAi4tEU1/YP34aHQ4APOrtaYjtn
fEejCWfiC6Y23RUEW4181mWHPLnVt3C1m/vvmkfrJV0UCimoSUxOpEMxTEKG+Kp/w2B5Xv+I2vMy
Rj4Cl5DVgfTOwUa/busvaFL+qRL2E2mnHBpuqmh3/aCQtTHp+Hv/mZVZnpPXwj4JPH8SF6AB2AbD
M+P8sy/dvccdYk+3p/G5xsPhSt1fjH3eUMgELtVFjl84oMAt3chxPVMb0RIO5aJuJ+NvUzekVyCA
wgTfZBPKARLqniBOIrqXDm72acRfWZlVFqc6A1DD6vlSBu/lgx3xydsZlIrNmjF6OF3sznLShvxN
SgteE95JYXihQg1a8e0dL96W8xPLvO1sQjP5uAnzGu4D80q+DifnBbcsXC1WVbAzetZYw/kIcGEH
66aZxbOIOgF+1mMUxZzh8+HI+TrA6JHnWUCuhQyuze4UwHIEts9Urakuo04fnSuYwDDhYLcoJ6TI
l8qYyRr/3y8bzEaiL1F8Kx1XpkqcZ4hCwjbQskaWpSoJN19GRH31uEBT88HLg9XhqxL0pN1JAsMe
VKNooZN6cg4co11XFtn4+yzvhgjtqW+4CsghVDpypNqgsJHTUpgZqY5dhfMfIVNk+DNUtPxRWQJk
Js6pXW8oxQhoHFlTau6mGG940YPDp4RqvZEgEKjie4KHd83978uJbZZVv/Pb3J8Vx6JwFCGfVDin
/1JS3CIAHEpDVBZ9vynebDHVfDmmOvJRROwT1CPDukZNzLR0CLpexyhMmvExI/YcBevOb/edEUKZ
bssD7fIU/pmfh26fdqrFY8hqrjP6UD8eB/R9Ma/cryb9a9HFH63tv2B9gLoeP22eDLeVDA4+9QiF
b8XJXVk2IgNEbnXEy39UaVSjoBQZTkzt9R8CjehC9E/2+Xknr9FJRFYJDgGNEONOejvmZtc7iBNC
JqMq2YN9VfMgmvfXrkpxPC6V+Q3wsPLnAwYW8pFrnkMcF9Aevu/84HD5x7LY32BSVRmTkqPxFjG0
/CVuX+y8xNK5HAjtBvD6W87B2KGE6NzpIe8lbuGa8coimyWpERDD5agYdk9fSznWCivRyzEbkpDv
8VRhy4hnvm3JX3AaFU8iggqn0y5Hrg/eqZAR/vNQ/NGmivu4ikMym5/VLZwu36ZaPQCANZtfZVqz
6Banbn6RDjSlQGBuzoz3YlBdtMYAZzs7uC9dedTKz2KBFXzgPSQ897EKM4+SxB7xHr7Rtu+NQEke
rxjPr10dL9JBD6OvwZx3t1sskgaH6KnyMDmLvXRL25iqj73eNVX6jkn/yrwdAjMv+LMA4gNrCwiJ
Kl4lD9n8wypL5gFMTtYbQ79IMjtTwChceCiJ/suAu1f9kt0gn71Ay8P+XB9a751w/KMqcAiRu9bm
9vqyWV+1eJaZD6mm4ZYK+EWMqTWumiV8lSQq8OmIlK/TDxb0TQXlNzn4BcW9PRML6EcWF920fWi0
1HssYwbhLLykmLibaxErK1IQDwwgFSb42KG9E9J5et/1RhLZ9Uvmdr8NkeJRS/ybclZFwK/UIjcY
U5IRgz7TX2gTlwdixS0HnSt7gzOkfaRWdfDr6mY+EN/kNoZ1P/Xsg4QPkyRZHUXNaq00uOuMT12A
euzusvtPPS3OZIp81fmY6BF8PAVy/f+VukOzMdnOKSVgNIVVbih30Mt+5mipu+YUBYl6Jlm9LV0J
aieG37PbNSoeamRcnrSz/FQBmoERZTjDUsTgjqhTDURBYPyj8nsPXmxNf1AwQdHsIgEutVvoQDN3
VsobIZ0kitgXEI2KPD0pqZkoN4ol1fwIwEJs1Nkvo63fYJbMzQ/kr9ItN1pbOEq5uwHC2aQ6gIAX
hfuq8PTh74e2OUGEt2dJCsoguT4ivARZpdbb0u2j8/Sx7qXWIjSsWDd6naoNdCtz+rm2uWTtkbgg
96pyIJUcL3mBUPy7MvwwbTzBFHtXIO9NIdFphR3snHkUOr0anYpHtNLQWvAtOGoHUswoFePcPoVV
xibelN7Vrxhf3GP2VqkbuAGZ5uBueeX6Zs9ZNzdNLL/uxtk2cwzKeat/Sq7e6fdMQ3UdyAmJRCyd
gKAwkbpgX9nILCZ87VGb/KcfOx3Ld8/OswYWsJXSL5ALA/LkWBA7naKRZASNdkfyUsJSR8eUIJXo
30wBKIz22G+xQMI1VVb2+UG3ZosVnL84vMWl910mkm9sn2KOxKHz6Xt4+p8GvvOhUMWSAxXcb0+M
2A2Jubc4JeWP342h1GikS+3Wb+jTjrfhWMioFV74y4xvtgU0CANb2BITGUpE2vuIOeEo81xoto9y
bqoAsKildAe1XUnnFka8qkWeCus5dEPus8tY4o97cP3XRBSJdxr5QoN2IkpFYMoPB4mAj+74dGsF
KCNTJ1VZOq2Z2+S2lGmpexFtjsBYlnRXNaYAmO7ZdqTeDeGCwy4UG1lMn4KhbxQV994oDvL2Ga89
N9z10ZtN/6NJ44WkxAFmvdHzDPMZ179SR4Nuf5tpv+2CDr8H52xsOrD2IogSbSF84u6SAPjvRpNu
2ytxSNhwLgZ/vgiF1WDs7hH9mq6ysFx7YfUVIseOiYzxUHUrgm8NyXe0jBrby4AQeylMrjrtQROy
JrnXm3QhY44TY8k+T8KzKxEpXwg0EEua0kB6SKYdDgj34AWMTCJFGKAlCe8/Ob4Yo3XG7F2DmV1y
DzTV3EcdWFmUYCA1EdJWxDfv7rUxw52JsxaUIscu5BMW+hmgXYP6Uxkc4UeSotmihBtlkJTTnGTU
7cHW9aYEpMEhCoojIQVsABRFvY1Sx+dQq6FhkElF79k70zy8U/xuro5SaDTLEnKRC1bJraUml7K1
77ZWMODpIBIj89fwG98eatOwI0js9LaxN/P6ARr6oJwKBGA6XdWsbTHnYTOvspu67NGRTHMJmMbk
7FW3CRvwknRg0yvK5B/7W0y6X7RpRzMLnKp+taJ6JfToHiWk5ycFkiYyOG2gGrbcZi/i7tGpdYM6
kL4Lld/0X8ECKrqQzpFcpSakYqKZfI9TnXwdRNxLhsTB15EQgoo6+1dEa2arTwEQNh8rJAxvh38c
Zfdea6L+cn/lcFj3SRSuDXsXnHKeFEUIlzuUwY21FDLGfq/zT85nasQ4FIhDk7L1NKANETeBpXFS
8/OvzGRcmJSlVY+pTuSfRB3ykf9TBFnPpAGO+nUyF5o6ruZ1XxL+SEWMzflSXPoRC7dagN6wqZTn
fbcvBQEM93RIAjDZzlOi5h+vqZQTmxWYprYLo4xOtX9+gMIdYvP99um0oFKl0/DL7wOcrsop6+Zd
oEvNXrMOcqI3QN4Afpgwkbu1wAn4qX5onLlYFT3Rcq8UTrFpCeXU/2ZLxTWR2M95khodINETBeRu
rK10qhA8bYEF69Qw2sM3O2U0Y/9ZVTmEAJIUXQOmTMnnog5gBO1WaJCmIqaVcoZ9UTUy5tPnXEBq
VY2A8Cbx+CEJBwX5XEPI9Pw95x6lNBsG6XPgPdB1I1r9TikellZQP8alSNDKmYXpqeUWefQ9FRAh
hn9/S6Ty5BP7AfymE6BLiT0Trb8K+o8zsePmFucyxnviV0QQcklcR9B6lvEaa/Y7AKq900iYNJtO
53rf9DtBkc/S9/0Bkmzbs1tgU4mi/o12Ft8GllDezQGXe7IBDyM3Z50p4aPUPH2ugZqxP1CvD/gA
+S+slhuLAEwkB6EFVtPfgezIuIWUBh4iNxoDvv4wB+8AvoHG6SiktakUqjCTL1eMx9cOVy40NWg3
ASDLhHTOjg+eS8dhIrr9oswwZLFqItsp8uEq2+PE1+Ebq/Tm/J0Wzq+FuJafaw3c9TSjCjz540oo
M4PKVAxPgnYAHgfwJ0uio6wrzKX4LcKrRxvDx01vpOxR4LX+B9ac3tIxBUSdtf6uLAr2VGohlqh9
5SwaOsihqBBV853N9UsrXFUB8aChDPTQyVdJP3Ys2wjdP5jPhNjg9ZNk8Kk1iP9kJd7nMSxD4/Jf
N8I7hnpxpolAhEdMafK2POfgBD5mSPBdcnnf0H2yGpz+jSnCw8wKFHzfrQv/Jgl3JU1pZp4ReE3y
8wKfCFyqk01gTxJZ/fYTiCCgMd10x3FTze0spo+soI6pnnoJ9uke59gQPDvOwGNzX4NEG0SucnnX
sYNVBA21aBy20iEj4NBMv8nMf56xx+noZrrxGbpA7aONKNYDk8GSvIFS3oyFAdKpS3AD3Iir8jAn
0FzksE/eZTmJaHgYcbkdHI7rXmpCXd+h3QTeiQmWmhnTA1ya8NAot1V9O7OVEMpZBEO5OncTX9SM
bOOJ07m44ktt/wp1EldfQuAXQicvx9NSOlUqou74dFDLqxVVo5TMcbsm/MxM+l2i+9WEhHEk25NA
EfYsHb5G2juNFES/BguYmmnkoC9sioYROXFDm014O2hBBiKTvKBYWk/G6DlDjebb8kPoAeOG5knT
/kTAQej22BrbslokY10gujV55KEFkHWfo7rQCHAz/mAuEK7GK2S6SpvEklZVQbOmu/vzfxgd5fN5
ZTW4cOrBI5iNtJA+6iMi0PPXhEv+TxiWgJ3DRPToZqarewuSlyQwlZ/ifF7990N3o2u1UTHFFW0+
m6XX16L0c5PBID4+ZAtdDJHFGewe7XNSvV/gChSYMmVM0YqdFtIMyn2uTRrZCXEhxdS6mcKbBq7z
2xvONX5Bw/UhQlicmFEOk2NaV8DZ394eqVfGvNeaEXb3JdEseBv2pY9dXDVelFtQdHocyzfOtngE
wyOfMOowL4jsnI0QEGaUgu8OpzCJf4rhXSimR7kQfsQbDe9TKNDe4ZP9ad/+LbUSKg9asOGDOBLK
fiLvPqsvokKg4C5mRh8ZfdZfoQazERtQ3L3ZEJMFW8raCJ7m8WB0TBLDkYRFiSGYQT11FaLChgn0
LyNGHk5zaHuiAWU8ifo6vGhVmleNPdiy3LtyYFJIpWZxZy6CIeyJbOZlGCh4e9PdQ2gUVyy9yg4I
+lnfCG6vXAqZEti59Lk/EmiVC2TxKeQiK1ToHJUhN/Hlp1apXnRpGjjdBBMVYO/fP1iaBRpv6R8D
Onpv2FdqjjkaajcQoLxmr4ibknM1oAxG7Q8YUTJEPJ9VvA4qYO9YqVDLha+xlusb82JNQjQxochl
qWwjFHvdSd39Oy5kTiOIQZPbyfE6sNHQcfY/xhdQV2/1gY8yUDR/9YMLLsT+KmF7OhmxMQMTHLRL
nt0l2fy+/5U8vZcB+TNeTejOuUoaPvSIZSjf+d+O5nis6W9+9rk7rPA6QgKipyrABRLDEp8XGWBN
Ol6UR1UkUe1oYtMm+qwyBINm0lSBz3ATNP/u9biUySZr5vPE1K9EyWfvWHRjuXm6xI7nBU0LtD4L
R9uONRPvH3bI58l7mAQhOD5cRmB01cREaOy0mKluToqceD27xL2CqL0DsRDy6XObuQAYetrH62NS
U8RBQJBYXkw8+kMO/lBRf3xMc9v9isRp0EJE3bRLcMUqNfNvPAY8TC67k9sTZjvYVBYlDAXC07tZ
8AvAXdFLHsYiJTXMBv+vCiLQQZgoeObVnSvuvmS9LKJv0hG/ShEUOgLwBkZVOLrTwDhhK3irY27J
b1GlsTHGCvFLk8I9byYxv6pacrDmdsMIK3hE1UqzeQ11AP1cDzYQOd2xjez7iwyippx0PM0tbtSa
IYuuIIxKCs8VQuUk0u3jwdneyn3BUdQnxe0I5wLPownfDDXjUgxrp+QF+CDBlLh7b0rNvC8FwHW6
rtV33qfvRH+xxs84jv9D9Ftv20P+UzddwN+Rd4QOWIvDK+BTqf78oy9rEOb3b6gxhFPoa0IXM7qa
UVPlq4YG0041gXPpwrp+LUcfayy9B0/bQVKD7iDSV9Ku4hcQbq3zHTX9Brqc6wrLzdO3G/4fkCci
4tZnoeC4xcWjM8V6az6P/xrzIGLRWxVExjW0t3bCTd4dj7NO2D8L7qc1uXAa6S1FemBaSThQHCrM
DM1qNANrje3AW+HU2JPVTvOayHZ0RWc9qSEcSMRO8IMDNGhsiHjjOZPMY6j6hWm3gymwtVw18mHw
raivK7ao+j4TXZ1jfq9ywxrYP65PTuy+B1on7lZhADUkI975L+cWwyOk7ZN5/aWpXiqEBhtRDBzi
wcgmvG+1pd5/mF4hg+bM7gC3kIomTuGHfoX4ZE7D8alZ9yjvsuAZKhnxgje2uV6sI0ZrhSOTIsrK
gyY7KSnwKzeKzA4fmd9jvAP1Jr33aC+6LMTQyYaLhAGgLhMTFw9UqB5KL2brnPU6b14TenqwAvUr
DpQRdMKg9uJwNTupbAO6Q0jNrsjSYAiONjTLtQanTkc/RJtGt6gxTvX15rFGb/QATctGz4XPSj4N
wOVTcUb/lh+lP4rE5DvREg919PCBZI0f3sziYUUuofUvJbh5qeMts7wqvV9UkDs2ofjg02WExt3f
ZqiuvlEiLQwYZr7P2CB9ZQXXJJB7L0tNfJv8TRW7bqi+8rM8+s/8T22TBeYabYFmwQGhnenqcv0L
aQp23QSKgDyZ4WIi2A7wkWrjaOVp7i9QEUBvPltwjIgVHrwXPc0BVxF9J7ZiEwqk2AQAdqBIy74t
Ss2thqKReKwWdfSV8iltQvBPDT9s6afGBoMlgKeVw9h8Fi0U1XbkxorObQy1rBOgqf1f534euLjW
PyT8UyNslk5i7pY1a2m/xbjbLS/BvSW2UT94kjNK+bYLgPcONwCcEaqnZI7EF5zFqbLyl6/eIYAT
kvbtwAHL2awDUj/XajgF2uRGUhXk2oPz+XFLWTe7liAHVfdADJjEcXvvbFwDjdJxmJggWCSV1+et
Myq7CZ2v8l+b3HscPC6CWeLA7ifqvlILY5iVk3TzlXLGJQqG9b2J14HrlbT9DQOfGoQCHjTmYZQY
8ZTxiPyM9TYPsa2Ft350nkJ5gSOAdralH8d5LrUYGv1yDtZeWF4D49aOJ4Vfcaai54RwsSJwvabs
d5DEiU1BjjybLSnhB88NgBkbRreS9FSjYJ00okffBmgdL/EN0r1dwdEsNCniUqPOOysERFs8aq1B
PhiMvcsLFGAuiXRFajTf+SAJVO0b5Uxn2X22/ugyMhcLpKPTfJkZbJETN46/pwAlFivzrJJAKXAy
FAEq4AJVxvmxYpFkcdRd5Vnu4tzFgVPlBSqacg05Yjtl0AekptSMsbdx4m8Mc4GU4N5PAq7x7LgD
lKC+bY1jfx13FwvkgrVhRihIfDK2bWneYNTVfiSI7MXSogx6x3jJOjxiM6SvnSOBiUW7nkhA6hXH
aHCHJPpNkxaPKh7R2XnB2nfNt12D/R+MAZ4qIviyPe1pBdBhOPYRTw5u/113OeL1n79u/PQG7Ncl
Cf8DEmcsRrAR4RZDz51a87KgVP5oE6kj+VCmLcnI4goThAaJIQCxnc/xgPF4b+6yVicgcbX3WL91
wlGl/yR756lhkFizktrwNLOqomzz2lesx90Tql/Rh8ZnE+QZI6Ni/ZjBr/TBvQALpKWqzuOgLW2j
fdUE2f5nZkFVWH5QkHPIVzE/5urWKAr5TL7GpoHUlyYqLalcRaARVjq6T0kSvI227OR2xjfz4KaO
oz6ApRvvhH6J3Ubk4t5UJ6gss9YLzuAYumFS/xtRE549MWZmc2hzNMJ5JZG/tmSSoU+N91iwZPAp
Dr2+0Q+330VNVh/Oz3gG75pRrab/610DAJZ63BEMqmPmvPiN9ZwsRa1O8ubX3BBs10BwZO0W/67+
BhzebJjxuGcAm/30OAN1+Uy4pr+tZBSf1TKgFuOrPtVa9c5Wz2H4oJ1Xb68/fROyaSa4L8KaHtDv
00PJDUvnqfPIlAxGIzmyLiqaRyU9ANWfxzf1wzG6/QNcCqp+ycrTHI5F743BnSWVToFMjw1c/YNT
wMi6+9VHM6UljfkNp9QNyZqUSJe54EJ/RnJewVyqTNcxs2pQTY643yac+rHql21FMTHdguK83a7a
H86Hce7egsmTlmZ62owDDluJ/VnpwXovsNgL6FW7rZEYRKI8zCNbGZLSBFUZzWPJTa142YkHB7FS
BoSk9D3Jl5lu4oa2btEiRskogSK42VeDSZZa5qR6lsNfkx//SDFSOxh3C6Xyua1E4LKULASJF8GV
F8kdWW44DEqdlXxRwJnwAo5OYabSR6+zwXCgToVri0h0JitzqFBfQi8pZ+ZWTbUDH1HxEJkx6Uzw
/GgMGNUhep3NDv3sqUnuH5xa1uRlZt70oB4m7DE2RkVW++y6ulsMfwwDnokVvocVHukVFt/Ojtcn
vHjCbUP+9DW0ulGE+b1E+XlQ/H5zX8hKK0Vuc1e7nyfIW1dci+0SwLqhh1Fkhjqf6RynP4T6seh8
sRSUrCJwB0NZdQRuh3CCMmPtzIKUihFMFRD1fx4ymmYxsyY5Ic8rOVeBcvBOIj5uKuphlA1zpcpL
J3ah1r6igGBe6RAi4rJ5oOLxNwXWC+1cBfHyGNARZqDoSCps9TXB6085FsbiSor/zOTb1juBvNuU
g1niyXyXacgMmQFvSQHnWG4PQrCW1SelBRpqy/yMq4nGfj1yWvaq2tR0Qp/bAe97AA4D4D+B81mB
P51FlQEG5RPldwgyUbxFfbgz4ePbylJiM/Ht6nbq6BwPAx12OvARE9b8nYS5NPh5m+127lsvUYgs
tjSTpkmqFljPZzSBDhTGmCWMsBtu5oU6x/HsK83yuGtR/838nmKIROjJl5/pJiYrsLZ7Ann5l4AZ
AILQGoLiSoSl9JXNEmrKxfMyOb106/Ky3S+x9y+5kHhQ93RL3fAeHjjQL7FhpADKFeytZTe5FIq8
0VKZPFiPEmE9Rqc3fxP3VyPcmzM6kTPHgUhalTN+IVRabhZNi/omjEHYXFBJLm2ka1tsgps5Zike
HVSXFw6cXZsUzolE2k+PhgYUhJwbIrqG5JFaikV6pDetYTlNAu5nuxXfaEQWhx5Vo4gTT6zDw/w4
al1qlnlpEvv0VKX860XqXn6CpI0zZzhv9WU6/3MbgPkFeipTlNFlWtNjmjmnIHOnwJ9U2Sc6qMMb
Rh3t3iXuzIdaKflRpr6UAdhMlCtJ9tDx6LjNXJn5s6gP2LWMChd4Nholc+/JdFjxwldoJEs8DwsR
UZjDX7WGHuWvtGB29+tjUPcRdtcB4JCPCogKj0ilsM+XXZNXUQ38HPlfmLUjbJq8isfTnQK/yn3a
CFqjy8wnt/bduOVEn8vpmfLvzAZo3VVnZyCY8HJdASowUl0o6QYmdRpqoLpSxuS82VuMcOLPFYqM
Bd2Gl+6HwVoUv2SJqRhIMGsZtQVU29E280oF6lRexqzL8MdVCYcT7EjDoO4ed6PRdJUmpswFnWQc
2eVX7DghtYrPbarQ+3BztcslFxBvGxF8YugqXBKD58UwlfBNMcCMQYQpL34/syM4BwejO8qER0Dy
ejRv2NQzHVGpuQlRzlIkcSMhmG7Ki/3l8PxHa2mQULPYbkBb0EMW4nvEatdgpRVJipdPmfI3KQj2
kES98WkSYgbuF3ClXBup3yQsy/orFAz4g10+pESVUHJzu6HaJIypFdoJ+1UBQhMbB01s0nL+IWSX
nMt1AgE38GiWrIbTVILJOEMm25Zq70a3pT14wuHcyjWMQUf8pnwbj3+y5/aDq/y3TqoXvwcl9t3g
2XMPtBaXlWizx+cYtFgCJyQu8b5MWgALwgvGOhhvMQX8cMQmgV8ot9/2RxziUEjUOMbGE9Nz8HQ6
LlYO1iVp9P6MDkVLP4xOdoghtFRZbQa5NWRUD402bjFL+qH6Pdulklsh8BEKF1shvEAj5M76C5tv
3J+GEr+W6QXBWh7wyIQL2/itCEFxpo1xc1rMlZ0GmpRHtGdB9K3hgxJZsmENRCbpGwROsuG3UOC7
82pCNfuzAqTtACvye0ORi8wPib+stEnellAPf02I3DU+I5fOkA75B30j8Cvc9nEaa+juPYiymDQH
b/D45ZSaUnsXAhs6p1+I4CS0Q6Vz01vufGdOyE7y/Bbf7sq8gWAq+bHijAcwGCpyD4nE3PqiMVYL
lbwhrJpGlrQ+mFShNS48LdExhRV+AfxIEdLvM/igd+2DSeo7xpmbJ7g+a9/A/1AkGzC896trQwyp
YztoHT0qwj1BvasSrkclr8IPbzOFdu6Yr8ohEXfpOrP8YpQ0wHPWRZlc2PVQ4qzSOlkJ1KwxHHX2
0SVi6ihqT/2IqkZomfzuNv1WRtg9C8lLW/Wm/qWCtzgDFLZkYyJSjR9xP14cCR93ogelqyP27czU
VuKJG2Pv7YtrRXSKuL3y+TbBB3M6zBLNFJaxUeMIvnvwqfuMxFngeNFA8yABsE2Gq7CspZ/rOMpW
gU38xsGnwOeMDw2fHr8sv4Zp8fC5kIMqFHpR/CNkItjzT6YLMCoBQQGU7s10Qu2b3to4TB/AMBIZ
BdlIx0CQSec2vU5AOoVt+g0++xNBnRy1ovpfOgEASIg/ARLYZ8afqkVzr/KfZpsu63gsgLqYQ0Uk
F/z2zwrxNx5DfyGj9a6hbsJxbpDdcoQDsm+MibtYzA7wcgwIXIH1JCDkdjB2WhIo2zXrGYUukWK8
oUqElCQGXOX1K8tHDoWVKWmX32JmIPBoRf+G0t+ZrP/oTGhUbAeYQ8ZjzQt8HXwYIF74v65WgDP0
Vt58CqNe0B/2RWPntPEymhX740Kp48JsLmOWkHDU0wHq+yDp9GHtB02YAVAm4SN/KwrD0Ygv5UQi
scGPo67o9LB7ZCz5x/VecCm5E9kn6xT2zeis9mpGbd9rvM723Qr7FCnj4XXWR/voslgMnl2RxXyN
TtsLPTCGhv/W9L8VEARe2qsqqkcRwXaezsbI+QdPfL+eE4WVswCPH682Oy6pY7QmNnsemR2aOBD8
04pBEMyvgWUb58YsyIcybk0/G8zCRujib5XRoqgP3hmUqAhzXiMALUkm/GdKSYkLOsf7IQO3YdTq
TEPsXr34j09PsJkHPdZHM6xcwpyZP1i016MdNLvH+swjqVy4e6q6uJGXKmrY5+VFGwPAXNk/Sz1/
LzNGMH0JjgO1Kj5+cdQyrzgzkdBUPbiR8A7exNCvEERby4mIZ+AKk7K8axqdyf0MZj7AuUe+9vaO
7lXIyOyDAOeSzi43l02yBjChb5hRQZHzHImm2qKtw9MvCoJPsKnx+bQuXGXy7kRhF5BuD8YfdPzC
RwzQD9oICOTSIw1QEb5K+SFBwNgfOExWYmOzOI3ymTD2+Qo9P8yVaL4DPz+xm9m0avzTSYtIdfQv
eLG9pU4bEU/3TMDzZV3ckL3jxefm15TCRriigJb673cu8eGYQDpfmRYlchHrvEvlks6a0rhycthQ
ZD1u6YVMTaXuwQ1uyf7TKvzPhrydAOsRbjqCNlSXy3AQIi8k1EGp5XAIPdSg5jSmEGBAAfDbMgME
XQ/KCDKNp1OAZ0GSN3PDf/tTdMDcJik7nKJC+ZTXWSs4/mk3tW6+hvJxepRhw5hnbXpNCRMOXVxj
n+1meXtxEe3xqPg+8lLzE0GAvjbdCnlMB0ZLdnEjzaCG2uIg7aIEuygkSLi8LAv/8N+sA+yNbw13
TRUWdsMeHhQ+GTpfM/2GUwgVhZqPrTCSe3I85weaNPicPoA7UPTnfXlohZOg295jz9z0Pg+A6Wwl
ZKFANhJHxFJzhwjlw7F1o78gvqtrV+g7s/832nRC2fMDMJIZP+gDi978BfO6RRp4z4ito4JNoYk3
cu7E2eBFRba8Usmkxn/JenXFuidsqKQ5i/41SFZIQnnPorg2TZnc6vo29KSEQJXx0vA9OWRD3tOB
2/W7hyNdD9rpqoLMmhZK8JqYVvxLrze1KP0Q2SRie0pBLMLA0OQ/z/Yn/jD+PbOQ6U56BhDLlEaq
6p0Z2h4N4tWikW/jXO/JlulHQM9HarFRKFgPD/X58gISZdhEk53JhtDR2QXB/K+pjBNwQbpm2cRs
pjU4VZCKeDdlekbVnghwvyaw7V2W7MCRcXqidTlvLDGvI+I0TOMHrSg/Mi9m31KiGY5OFG5o47Ah
3PDbBvQc1Il7TEq7AlI6KuER7ayGnVx5lrggqShOqw88BuYiKwmGZ00vV1VBVOfdVtrhjZ6xoCSm
SvxJ/mXuSNaLuSp21ftwcD+Bl9zg3p2vROB64HmhtqTOM2ki7LO8W3mx9KsQhIMtvJR+Db/x8iFD
C/A6CVmdiaUm/1Hzf9xzKlxvi9bU0SHIrnkRqIi6PSafQy9LVGJKYoWeC77eSQ91FKdzI5NzpDnM
4Sj3BtjhlzBg8fhWf67tzTREw15l3fbJoTrebBhPnv6/M0h4nAWw1/RSgLVr5Z8L/d8NYROy0aiX
CY1FeLHkoYjPbZV37/NedUuQXgxm/zqv9TUdgrY1H25wVTQsa4HVLrRqTR5VqrKou9VQPu3gV0de
RkHUAsYnu4ZR+0um9de7tsgEwiCC7+aMPFI0RISg5FJDEj9Q2qUASdfBxh2qtUy7fFnaOqL6mQ2J
HR108IYjAMlOjmarHYulCYSD1kFx2A89ZYfY53VBhOj374ZS2B6UctyZkN8CQaF2zNqmyjvMdG7d
U9N9QNrqusr5xCEpQwxGZfC7XTbBV0A2/KADewHNPJKwenG00dV6NgjWEX9LjM5jj2c10llHWUVD
za5dgFGdlg/uJ3IXgfj65jLqVJUtufbdMP1JxSWPh0zoQQdNMDLGAfigeJ2wUjesed4IwVy9iVHF
qndwJyCGnEp3es36cxmfYXICdOX4WEqpMTNNifn/NIbGqpCw0Jz8VrKrBb3XXj5ofXFlVioxgX4a
0OCdNQI4/OsgBxIICQYfrl7PbdBANI+x8eA4ryW8sm2y1T7u65n/hqbqJSdaPbhMkVOB2FErFFG/
qRpbsh1wa6VK+sZApofusBak9x7LtvfdeVMfk6xeO5J1SxWI61LhIASVeKXmdWCPHxaJj8qheWDD
yOtrqX2Y9gwze0/nKyKnYCjKAs3Vp2NqvSGf76baM46umAH+c2Scj/xptnf+v5pvekY9RdT8q0Yh
20p+16WRZZtlIVwTeAhfUUUmf/n5nOJFYgJXzc60Xcl7W5SruziFBFqxtxDU7IXiibLAnaJRiowd
xo/9N3KKFLGqMysnMdtgRRZDgrfsKdz/Px1w5RN8vd/5BlJfaNwsgs+h/6FhtdhpTW0TsGt+9ZSA
xT9W5X76+d221hCeM0BjQhW5OBCNVHyVF6tMcivBbyJQ+g3+vZnixWM8KYsdO+cXOeec1YmrABxy
UIlsblzeCUJJ+H4ZpLbekJkDjFZbJ7QWokwnuwNtbx7gk/Q+YH4K0NAOce0dyT4kSkWiiEhvr6MS
RlWaH6Ryt+nlanuHqMqJ4T6aRV3A44PXv9DbXZsLzIIXQ1GMIadwF7PBYa67bCYXBIbgDrs59IPe
V5XUOvo/Vso3Xmzh0JfsaPlDYBh/xtvXkeQGfXljRuksg96kEO6o2qFCMR9mbgybHNWY33NLGMFR
3tsMVcAj7VcnKQcYM+SJtTvy3+BT9ta2Gb+Fw2h9X5yBz3pvvsI/fw4tF5iv65CRbTGi3flAjZnk
FLhPbjnUtbRBwB0k7Xe0r4IsjNMQsDAVMDGNheH68V3fLh6NN/5V//BzH+9FWdPLnMNe+I/qf0ny
8u+VL0JIyU3EFaYzDzfFRW0fp9vZFX4dl0c4cHNHu/6NMoK2FB5qsKGN+aAVXO9InmOntCN63/lD
7a66sxHpyYNET+KOqqVLqIitKrebm+ee23Zoc6wzL+s2w44vNmUFklmEmnVh0fmsNhH3UcV4hDuu
MbLL3rEFsF8ZV/DfXuDivtVUleIhRkAElA0Iwhr8zWsOP57IXGBUPyT7UZ/1Cb+lNcx6pfUXvoph
hVGK/eQ6r/KawWBLNApuN6thfnhm9x5vf9cpb1Ebr+lug5qm5W70QOtxVkKocnxtT5wFJyS1WM1h
2FnNNPP9VCjoT3KJC1Mxqqs9hwpuorCz2CcaiMUcwCrJCSpP8CV0DecBcVmqcxj7ZsLwQW9SCBxh
ZRzhYtGW0T6PeRgz8VS+oI0mW8HlfBhS10yhlrZmmGwFQpdoFqBwrCcrmRPHHxAfVVUVuaVBtRyw
zLPfpmxIf67nLMZUiN2BgeBjlM16m33xMbsBsQnWsesQPt6ycLqEtTGISoaSy1UKD5JRqLkTTMpM
HKsaI+ex9c86x1eJnJSPyPC/E+gkBfslzfcMXp2z5wJ+iU9vKYs8LY5XmGpLalDXR01kUHXAI5e9
0eAWRtNSVF3S9HupCG1BgZ+Iq4sa87WW/0ZpffSkCBcnI6gAXg721bc7PvAAKUtzVb8tspWcFCfu
41Lg/e17leJx9WaBHMHJQdHi6AgaugMzlfiQ3DDACCDbMNU4benaPQ+KjpgCyVENVAlnUh6oNx4H
3OCtHTWfSkLIUm82ZykE4+v9wg12lfbJduKefd51uc3PG9jTVVDTDe2YAttw/uqQx8cG2u93KiIX
aA/1QkHeLcpBSPLxFGcpKAlBSn0Ds5tA3J8pWqd3vOlhTee4vW315z/rIOcFZQkZUvQOp5YlmNMx
Kri5AQBmXxPUZe9kptgbdEpCv4w/gwR4DrC+5B+sMqzFGrN5n13hycWXWuJMPCGXPxMITpB0NYfg
kyIU8mZiD9FvnFXE0PurKYg10aob7TaJB+k0qmoFo7fE/r43ajFmd4uHXqSGC/WUe1MCmtimJebj
9m+y8omXd44XPkTwE/hs3gLXXrDMjpLWO4ms3fiOHyETnqVe7Dtzx2Hb7YaCP3kI0xql17BQtpS9
Zj7GqFnngx1TAcw4Q4ZB63XW1q++NrTYV3VUCasxay2YTFbSULkLnh7sylKs0wOuvkthqXk44EpC
Hj2/3/nJqFi3gbMPHJM50s/ulM/X/ne+cr2FLk6zG9GMtGYG0Us0qG1Vv3uX7N2VBgnq1WXVwtJ2
bHXbfiQS5AZMf9t4hSoy5z0//eGegUnPuENMip4G1Qf51/Xi+19boxpmRAy+AKmn23fZG+0Z1QYD
zddPanLJtB1Lors0ZMZLLCGbd9Y3Gxveq0zWI1/j7P9tu8D5xYKsqu7XG/JcHvG0qMdG6ThWHjgy
E0Luj+H6ATtFIcOyAl7ThbideITW2UrcBDSgkKngNLPRfJLYLKGzuyF4lGi1K2QVMnK1Adqn2PsB
YlpSqzwWQt/QNX6aJFxioTmzR3LHltwpnIf5X6qTEYQI3yygpDqdXdDlo9ZS0JTnR3Mp4BNI1gBu
M0kC6bJOYN2XwjpSyejyRLNA+nnnK4Yb+ir+ggDr17zyjzeuKx0UFv+rNKyoNe2lD2Qzcf0JgCyb
EMdkevHKWjTNXbXcxusPyJOkKe1DHs1ZXYEVAFqzzYV84Jnk8UmTEMTsYp8L7YhvcmbGceBZ/pTd
+7EAbHVm80CG7nLKLweCEOled3XnchrK5eNUUcd1/+NaOXlKeKFkGzRrxX3078C8YYFs6wyjNAbm
mTMcYwIrxQP86aQoz211rWZeDEfkrl/w0JDOxhpOxabQ3fspNQQLgaA7mWnmUub3ZkgMSwVCAs65
oeUejIJbhXK7yjA4YzqW+ZVsFOczaRl+10Zyl41gRA9UZQJjziPWolVtc1IhK+3BWZxg2MhBOvG3
5+zYkJ7mFeOKIhqEvUwhtseXVdVhIazqcc4FZfgn/fbhE+cN+yBumR7a72KcB6VpiGhh8gMtD/2/
3hTwWMJI7ugMjFG+CU105nAqDxRXTHYl9FcHIDiNDwfEktuCyMenMNi5S0B9GTLHwB1L+wcTgpRb
xT2fJacXDhbUv4tPgAs9HvXuIS/1Qux2htp0lpSC/iVFkf98MgCMKV03hi/BF4oevGymNXsl92gc
2mkPpf1MrkToMtaCLuTmc7/8XtFn20DMPRNK2WxaOtSeTBCybPw2cHa2ggN2Q6qB1YxbnP7VkAyW
teM9aAaptRYayyEEfsKzxUzCK1eS4EKqLPSrSNBxFra9M7k3VmmK8ShOdx1BSb0R0/bOKN81oBZX
sP2LXny0aAH7cbsYaG7ZakuuzlwruhGmYV7haoAbH3rw8/j5WWwAA24CGldI9LY1URuQnZlZOL9p
TWaFvj8LSS70gryLglyWtz3DRl7s6PtQ75p5cAyjOatJJqdhpAQJ1UFWzEpsYll0ggxPTqDTNIW1
o0VlHxq6L6BH5iGIVNDoYBWKzUMKja/IQFzBkYclT0VBBFjJEgg1WOaDTHhni7RH6c2Gyn9ly4Ua
gZj6xIrcwBkF+UlTSXw9tZF00BcckrC1ojBwH8jClkgBuQdlEkMLhZBu6DO6QwivBd10nkC62erS
POoSswkde8QJehneMo6dgKncPadNMSmJGIQWIxmx/gydA8KPg3aA/ZKoBLDkT9L/Kjub8Z/3OUrw
OkDF9wJOmoFwLfcnbkouNI/nIassC05VNRLB3P2+U8gM3wx35iG5ZWm4RHHWadPhhFm2AmbWsdGo
BcLXUhQ3Fg9/A5zmqgzR1GWEughiQ2olok7dX4cnLAwzYZ7QJX13CNVcmku8fSQ8FgsAzquEcgfL
FWW+lDy8ALPsYyVurc3XVV7TObk1RWZKEHjvvHr37+3Q8PNoaPuywkG0Kc9OHiyFrn3m34MJzB/M
ZaV9MB6mhNCehlxwkO6KgjtA9Rk2kCb48f9xFwD0Bsgqqhze84bH87pGBwgErXYaMT/PKjnSUCjR
nAhUgIdfEY2x41JUYSG9Plohq9PIztPHhgyZi+h1hMlp2Tb5kc1M6idXutkLKsQzBwjO9V6lXb5g
CW8ROhmn4HnLx5Xt/DCeA0WIpQ6OSkQa/hIxJSLDuSUFqQEV1xZpZr0WZ61mCZRChvZmg/4wDOAu
Llmrdx1cUgTiTlS/EhOFjEG41M16+RO2LwRWqKT2y53PA8ZZarvg5xgKqDhnX+UO4OLs7Ko6i8Pr
mZ7Oe0IeYdpSuRrbKi4jeHydZSRAE4J7+Yn45E3tUTkS1PQFsMniiwsnT7HViCJFXqGoopp90nfi
/0KAMDwnkAINjNt40RweB++hjukcwdmDbWSpbXfq8Tf5kAWQABnCAeRruchzyry6imTC0QwkRQTH
I9UyH+bEYgTvRosPVHQa6uEplKUVIryWXisQqj9uu/KgApfybmajYtQnsncvqI+bF4gQOYew+/SD
QglLdypf7A74ZOm+wrOsl7TQoQNCZn+KqmSvwa1WJkUmNiYcxUBer4FZBxtiburVbQHGPtAHqYOE
p5rAepaZfTR5rWKAmpom0BJeAkCRE+JH3IT8VA4LIKC+FMO+Sq+ZNqpgh9im9ea67nxzZXiy3TiI
yXry+NCFG7cb87TBADHlm+s24urXWr5rqoNTqaaDituBL1aHNCmy17faEteqkNno0wbjMI9cu4mY
tvWG058UilISZAVwvGNRi+zj8WBfZoEpn6gnNlremRMzRhxa+e8CoNfYN8qHVY6m6nHSkH6qGt6G
zMGH+uVFXnG+eawvCdCRsTJXz5XGkJeRb4+snExVfpa1Tp7XMBChboKOgalSo+1Tks/dreldW7UN
zLFuJ6BXUV1ENJg4eBwtwVjddAyH/KQaVWZL+tv9sbRiKc+S99SKwN3c3f+kfSGOAgwRc+i9qh0y
lzBt4gK5IRTBE7YfAulixZ/uxwxUrQ4ofw5738kStY5u955b1ELUkF+pxqTPAnUTNeTFTVx9GKvB
YxR/tZPUaMvh0YSFmngenFwCsdMk6yebHnae+EN5/r1w4MMHwAExPVGPJzuVtNaFbmOy2vnQ4+Pn
0KxCuK7Cte9sm7KMy4mS6A97HK3QHlW1cYV9D0hawWkiETJDQos5hfuKUP+arKeILfYspm0aBjxg
6O2JGzX3grSRfwF/OAVrlABx2tm99APXmUPyZIRzxScMQ4BEowM5AuKcYcIdW32dJqTw2mM+Fvbf
BtFhMG9ZnaTmbYb7KL63NsyVb37jSY8IHi6lSwMhUYYe7DZMWUgSTMrph8QG4Si9FAPECjaqM8WT
7nOcfmNyuF/8B1Wbm+ddEoGOwF5jHpC+afelijV08qJ4G8te0JD/j3daVTk2yQZ3teDTK4+nOZ44
lbXuKa8cPjDK5UGYTH3OSsqdq/iwkZO4jg9vBhGTrS7qwHi3inVjkVUF2mPDWzsTPflywBjRlTls
C23/dyZaTybH1gRpwjiXcZUR24ZwiVOksV6DkreIEfiMsxcerLGZMIjFz9j0V3YLKb0tbQOQIKYn
ClCGHeBnDlE/80l3h3etDfrbSP7P3g7Dy0AKCMJhzxpNRcXKK2KbA/+PLEwdyvkrX5ZmDOysgocv
EQf0SlurTtuOBMiuiuzoa4LESDb47EPnUUOplbhpHxznhFCOn0VZX8fFtxrQpzHI5ZPwXk5fFi9m
Fah+/v/YbmFkEfJeVSMdjO+YkmuwBzpMwk1LGGNlYm3HalGMUxydhmNW0jiYKq4+tCE1G5jz88NR
m65cmW7UNgBq6uQq7UBO/gE7q3mZAqVYMAlbx4z/pmDX3GBWw28GWe0zzFY3Keng3idneyCw8h0K
EnSaJbgm0sItu+E7jNTDVS0qQReW9/hse2kEray9XicZ61DJXTPnjandqiS4yB065M60SZ8S42q7
RzqTpUJpY2dC+6LXH16Z9tth05w7F4/+Y7eh0Cmj4c8eun17vXVwcbySJ/+KyvBZ8C2Jk7QIZsEy
EJs8MfYgDRcpA3mF/YJ5uEFKPlwXGLCU3xgn0vgwY+UtUer62JzssK5RXTW90ql5awkTmqwkpAl3
K/wynr2ErD5psDWZ96a8O2jTCiykpEgaIu4PZEgODH7pYKKmcnrfb5eUZw4dNosgFPZWkXDTzbSi
tqptBoYp6qy1VyVLN1orMQXGR2Byoqlfl/LHO4a47N0Gm5HYCmQTw6N8lhJb8otAPvc0gXdCEFTs
aqRd/XYDDNXo1nGB2Axy4oA3MjgQp+9nD7L57GSPLiRh4duCWSKJJFKJrCWjnU6GrdKacQ/tlSJZ
vcxXx1AJ7F3r0MIBCnJK4uaNWaEna+r6/TkhXkbwbyXYua4yVNutaVby1xIc2K/WYoBC+v/nzoeH
2OORV3s/cupXae+MUMiqmFqAHnTYVZDi1k6QYy9dv8g2wbbO70PNzJ3oVdcxV4LbajKbEqCehmt9
ZiX8RAdakXJWwC1B7y1j3KSu5lFtOitJOxsOuq4mAobOPczNuaoHPjRt8nMPxqjmrUiz9NBtJ6kf
Zy2s74iyxPd9GuhzyO8ito95XrUO9nXKV6a+Odpu1Y978aJyoC9P+aWVHi/3ZFEeqM2PSNr7ERnv
wVsKNBzV1kt3GXzDB2t2HJfnYo+2vNa0FKnsz7Gqidi2p544GVg9ESfPRXH9SPr/iuXCCmBfBLhQ
vtrTtPh3xbATbIybAU57vk3RPOjs6rdWwo1tH+pZ+87W9xTRSu+B22QqvsC5KdYiQEGtsO0EnxyW
PICBBcV9bucTqrV0kWZ3TUY8e9+seXWi64MTMPCict5sHvvqbZuHpvKUODAtFJCGmoBFELRZVmtu
uM3BHpdrpBrctbujTdvvBLYuocBmRxnT9J19FlpnwUj+AJZGXKTlmgSLSbGOL8Ss6A+B/pM3qU3Q
L/s6GAs9m4B5a2MCSHMB0H0W67fzjV9eFlZ8XkO36QuK0PF4BE8gUanN+eofrsOACQ3dFtoi/xPB
KoBuUXz2bqULS+1qjz4Ld2Vw6+k3yFb4I6E7nYUjbihZTYmQ2h5SbSaPS/LErREjR3IKcxGB4SdE
FmPF4/eduZdLEUZlzZcdUMGJSCnDSt0kW6BiDbaJGk/hNKOUXHkSamk+ZU8G3a8Mj+CbBDlPkE4R
hZZ2ppcS2rcREXy7fTFBUIT6NJu5PyFebJhBVq8zP1+cUZ4TUxCjYZ00rILe7vLW/v7MQ7pjqK/X
itZLglM53KexZ9NgRTpN6RlHAQW1TBavRT8JX9/KrfrzytB7N7LGVG2E/FjuY0GOLvBOaACsmuWo
lajb+dxsC9KOew7/5erHGsFDfV2AbibwM9raMzpS4qmuRwlNgxW3H7byPs1o3zZH9mUYPV0jZFOn
k5gmvTCvYERCHDqpaNeMzAlAoNjGtOfxPDPQ5zNk6pS3B5yUfEKafg1cNKJi8IGh2VP1tiZVGykO
IthRjlZ/UpyaLnhEtzEU0uK4Ofi9VWMWHxXTi4fVhKC0zYmaUIDEw3vnaMi0JXDcPv7chGfvdKd3
ANtC8/GwfPNFYYzgWkznBU7mKczZscVj/biTMZlNpabRdLIPcJ9e3m2xo69i0xW9Lwyz3q8PrBLG
a8zi6Sqmqq3eSfQo0A0py3XMY6lK8S4XJK71N6vQyCZ5upHLCjvmuZuj1FV7WahxwNM5a4icMfgR
uSVXB/y6CCL4eVmeenUxc2DcPxUPlDGoeWHS47eFJlEDwL1y+1dPELb5K+HieG/YrDAqmNAIJIUk
I0CfsDKF8OVlb/u7p00nbIvE3WgeNdMxpiAN9tXbv65Oxp3Cctv1r/BJzbkVxwuqTxuOOUccwBjp
+3o++M3jv3imVigZS1c6/KO49uGsbjlBXP9oFZ/TyXC9u+GwFCgxT9Cq3NP4tdfC5/U77/vUmOkR
YYHt0obI52QHIRG/4ED+HyjAhgGjhqN6OmMEFW2EVx1qlCEC0Nr6WFMkSUhOh/mi9JFtcSM4Slp+
dQBnIhWOXaPwk7uPH4mFePw6v8hZJ/Rf20KDJsbBdj6mBVaakYuzyl6cK5Rwq6narQmv0xI8F5hm
0FadOQXU1VV9hAFebv7Uk9z2GDUovmAp7Rgf6k4OgabsQBJnA2bkzemzgbVeFiQ3n70G2m+5fvo0
ArtZZeqlln++N0Tgo7rLXTXgIFBPzWNUrkTc0A/8i6+cGJnTs3HbTunizFT2j3KMyaPTt6jaCpjt
J2NCX4M8NTl1ao1qoJHFJ+f3ms3POaE006gi+fBLjSwwYfshFbcNHaLt6w2QL9i8OcZw7pxSOwQV
+c1/Le6KmgnRHwuE0SSzpGW9Bjd5SquoW83x08vEmwe99gwM9kSFK7LZM2xX+y57FkW3N9EhaZzK
x+NlnOvNvxMf0lw1Uq/CA0+B/AlWQhw7g+Mi3rx1+Crho+naSplHM/KVyTAsmFZPR7/GUwaacEUz
SmQ3njw/ScpXUMMLf5m3M9ZiO8PwanE8mmXxdP/TaHLxqcFKyngVjPR1Q2zAttMJ6lnLLS2XEgrj
OCwc/xiHj/1uRTtkzAUGjIqVPbzITPsf3ozQ8XInMIoE43/Ryd8hWbFfLNNV3NkKcTXRyVkNEFpX
JG04J4/5C6D4848OBm36MSK0tzMrGxCbxjf2NgJeZ8UFrfZL89GRBSvhGOKIFtRU2JMgC3r7Iy6o
BMIAdgkfJmFf8SecIjs19xLLmB35s2ebMhMd7nyPxLq3XWqFEfdCminoiWTgq0z1n8k1fOVftuhu
reih3FWelvrHZgfGHMCYP918eNPy/F7NegTGg94hw7zf97JrSqx9mbF1tzlHFRuLmxA/FZe+rlxY
FFu+Em9NLYMXqnWHNrhyG44b8RShBn/bSvgoGlWXdQKsoAhXDC7Im+Lt71nKzEsvTFaOHWqtLCPX
Bj02i9dPUDi3jqAzo/Dju5oq5g9jHTLoFjYbsVkWL46wvx3wUmpX1PiiNpjYNbYi+nt/cvjLirQh
Kq8Lm61Me9Do0VqiAiKETa2GMr6tUBw1vC2D/eBvjMusT5tq9c6rAV07F3/5R7eTq2Y1uqjLc9OI
4Kj76YZPMiADY7YSZKcMdFbjoQgE4NW/Cj03o4TaYix+BNVC5yNSYkFlRYz23RuqCzBAkEwwGgmH
oVV1axVDcTIwPp7TSj7AOOoRmierXTumpnsjgC19U98xVWjRtZIyIQaz/eWgkLmfOkmIhOflbMUg
RXePDs986/luEtAt9J53Xb3s6PMKDA/Fh+zAeVmNo11XEI5nmXYkiddj761KMLQ6H9BxLFwAa91S
wDuFBXZjIy8AeYQ/On6IZRVs77MrkM7TssHfs+M424iEk60/7zRwaXrfoE2JAPb9hWAJMLTETTfw
7AviOQdqKKeXDRzRqrL8y03HGo0pxz9+erbngzzs1Yr8W81idilXZgr0blPs3M/5s7/MrSl2q/KW
N9BvZbrOlbVBygEGnZ3gH5BieQOw+lEroX7lMXnENBiuMo2xeOdeg9QQqvPN9hcjwSlMn/2PmlGh
T2t8Z4HOdgsgU1ZM/lWCcv+Wda5DoriEBpaA1s30XLhbcRtYNHWiCdrSzZ2LmYP0CUJ8H6iY+ub8
8KIDJpRsvof45yy/mhQEoZIc5p+V+wAOCbYZlYcc1KB5srbPj5Fsl04W8Qv8ixMgs1F1uip7fhps
Wtdj65B/G3+M+olbJNCNy3ilTUqNZ6qaylgPn05psqgce7tl1x5+4NPPKPchlXPDldpNaw0zKeB7
rvYXjq6Kk5+Rb8UgtaqavBS00kCgi55CpCuJ6evt3GIgNuI+jesugJaXyK+pcalKKeZ3pKSk6edq
3PFss8ChKdZuX9/LSVrPLYXjKXgAAeqvq/oPFrZR/ZAB+alqXUn7amKnxdIXDJa/IDqc+yvmgLVd
2l41UMZwjcIvMELW+B3oSMI/mrEesJTwBcDoBoel9g7TrLpxIJ8Yb43WFhbdAoeQRWLyRK7VhsMj
zNdr5wGdS7jjVAW8dyAXIkRDoaaUwUjlQzcgk7td8hQwVg1SJXQ9LfNRF+p8QpweGf7MEzd0xLWC
n4FOLFfAUAE0xi+KksmUhOOzsUmYQMVgFyC8+Et2SHnqJ9YiqnDTDTvsmjO2hhlLK/zhK2C+exlp
Q1Kjlpg7xBIZ9MIz5jFDRfde+C2poQuRm7hGy5+6EgT1jyvgZbv2e7lxB42x3yJYWU1aeyFAtpAB
B9lxpbMHYPFm0Hm7g5lktLYn5uQJBo/Os3kTMzY0LWUvZcWH9hVwzvAmk2sucnekwj8FdtkA3S7M
mFp5l6rVmByHuBi8WJ6NVRTTYN1boTLf1ZJ6FyhRySeEBwK1TOsL99RbyXJ1NllXL5EUyP7IATFt
IJtyxzFFa2FuODJ0G8mwXuIImuM0Rbik4vRqoxcwKSngLp6IWChv2l9IbNDqarTDRrmbGjvY/Lzd
K82BA4ig4O2DjDY+SrruXxFKbEOlkwVEAlqPGfXpc/13OR8tiXt2hEYB4MNkMxT1QY6gr5EG01Yr
HIqf9xUB5ZntRgwM8OpdP1ZxYmRRB+wcSiSZta1Y2OB4QjSlaZKWNfqVHdmo3fvEQ9o705NY4j1L
asKx8z+ndzh9R1vQdn4/CkfWk1gR3tTGdSEV4QvqITUfMzprb2ZGiqU9j2WsPB5QDeVJp8XBJDIh
D+GnX/47NuQ/SpdUEIr9aoAn8nBWmo4fWwh6pwbi5tfrfDZgHgmEa/j09cd4XGPXK24k3+HWi+06
J1l3LFDZnGxrNx1JfmZJ0d0sLzhNrIZ/7pIAPG2liovmSESw5BDgk+L3za4FBUQIjW6czCZUAZZN
bY7NF8L8kcxxTqOybO1S7zVYtH01aqDMtkXd4spOrI4OeEmobtrW6BA9J/PKfGlDqw/qoVd6/eTW
HKhfKOzHuRWIuKCRd+JLTsMSZOBaJoQJPGF+GYCXwmLH97qeyVuRW8V3GUZjE9erI7CZi57zDVCj
vr6cORv3zkd2I4dTz8FSjzPXdnsmy4ZRLJcmDZ/g2VjWgHRtLPi4f6zUHctJMtO+i1GeijyOdME5
yoGUFa5CynBE8Iwzd9AkdrVKflO8Mgpu6R9igDshgLls/Xj7959JMF3HROK9DFJ/ohu/9me+u60v
VNBWvm/Hqq9hShfH0DfcXGTtlVMiytUt+Q+5oMKe4SUlBKpY0ab6IssNLDYWnI7xOhhdPzVa2U31
zaSDkV7ItH2SY5qIm9kaNaG6vMgy5YfdhR/3S7iYr2091/2+8nZ4XE0j4IweoCtUqJcTPyhPCZVy
zY3HoQh1kk5KDEm8wrQshd9wmoC2HGbBW7LSFZoeclgMh7b0pbeHPDT0Hksk4uUJlph//lOvi1JH
TQu9KHiERA0sn7iOXzGlUpePo3Zj+8wzBDnfon6kqfBINF2+e4GfKuC1gWPmlEeJ1AUWe7Q83NGQ
6Ooh89hWpNUSliO+/B3IfM3/iqSkzpsgOxEg0lI6rTWFS7ubokfSdn3Zlf0Y0Q4cgDcZhrCJh0n5
buzg+MLUstoC9e450N940zeUckn7VeLP54UNXk300fw6sKuTYcmNABOyBcZPC3mibS6L1zhadvDL
whBK/fcikb7Zxa1k9tbMbHeB9fT9YMCeQtvLR01Jztufnk8cDr0SukXbm1SkEePhq6Xka9qzxqDn
wNq3PfhF/6hSui9Feuc8+2+wTKgWGxaF8iuXuDplXSqRKMuakm2mGEgMWyX8H4PwnjZXiKjO28Qp
jwiRPIPQ7kr/9xvMo4nOl3fpbc94MHfdoTNFSlajChHF9AMbCPveR3+ie1RKX58IoTR0aphrdaiN
DsxJNkfXJCrgBNQIDciLsk1rGn5YvyDRkMc7pqL7BJvxSbd04dL3FiwTpaZ1rrNVwklY6Ubs4Vw0
nEjp0XAXLO8EhEk+WIGqWH50drbUuybRXmZTr02ggscAVJjjctghjG5Xpgz8EN0VDRLj/IWAbt7u
Ev9LMwZSS4WeU6AV5lYhwzKXBbhzWCH/h6KGv6Aa1u43By77OhBaTEL/YPLEqujNn0az5aBqmrGd
sqoIQgINxYUrzdwEVQe0JClbCpkqRDjpXreznoOcwi4tCwihu37YfhyU9xKGxWHaYdJuMkYwpYqs
+SLCpKsEeUIgHgwIpoJx9PhKL1BAZuKctp/Cmt05Kit2gapi5cpAbgyzPfTcUiRwsGjePv1cLVcP
BG/yHJ45FOZvE9rKOVVYOxQhu3xh1okacVww5Xn2tuiTq5v1Qv9gpm+Srg+8FaV6BaiDwOVNAcwB
f8NIV73rg9d40IlwHZbr4zfZ+6bHSqnj6YdF58jqbXIs4LXvTjoUGt289USTWEtDmu9UMGuGPitN
nRkpoxVmJbQgaxIAvitW4T/GonQLU+l+wm5S2Cee1X4K4uqGatKkR0SIA2bEc+3ee03J0ipdv9kP
gYjmEpg34e2OJ7Y1yOhlMHNtz9JV3p1Wvz/mEb5Nl+cHu5bkop0znPUW08jmOBTYVLQGumcqDwYW
ku2IKr81N+N9vbTmOrPgPVqSsERHzwp90irR3+SxXoVVfXgyrtzHxNzatK/k4jDm+snYOZxQwo9O
A/rSMLaEJah62gd9wtCloO6B0IPdrgHojVhc7CxK5P6SICINRTdpRwBNyRoqbuX7dLYw1ghtqwaM
odt2bA2nlH8gkR2vF4103/Vla7hHgTKagarkpToNX2FHyAgTbzj9lB4lG4J876oc3YMd1LHkJq8H
wdd5DhYOb0+smm8Z448TP7dRfhzjoCu7+4PhRsCEcKFx3QNVPG+qOy0ttAFyvhmwVZIWIUSf9SFP
MzbqLghNXgyKDbEzugHgviN1KkkWDthL5IkcNgnXR3gW01d/Bo64WCG+YldsnbfvibPwk2er9Vrp
MQ31JxDmXztYeQk727iZttWftOZxgWQNBZ8k74MK/AiRAQYOOHNz1aakGZ504n0jTepYfZVPh1Io
DeVNiVlmXvBVWWfWjakDwqaynlbJAD7UhhGMFVrjqLzGcRmzBZyCOeiOYdXkOGKS7fQyaNOP/4Bq
GxWlOVKf+oND60KhT2hSfLcYovTSiAjyDMHBglxSE4slNNqIyyC2RPfU9WJq+g5gm91w+BhNWlqW
gsGNX4SU1R3GyPO79pIL/ZISAUkENyuhcZTu5Vj0dVzaFWaAhCVqv2hfGe4o+kC8G8SWJcSY5L06
pCvyRmBAhEvDCBnh5xLOHiKz3c6q4jKz0EjJRNU2/hklVFUVPZyQAbSLn7czKqZu4X9AIPIkCyiC
+0anym0G/nM0AKKU01AOjbb8iSGvLtcDetBdyMzDLTyKZvM/lpxCXeiaHIq9rkTKSCluHWHqNDbY
VINaTaucGXEEXMsqeAQ3O523aJIiQCo4u3eJBZJP+I6wKbkp2Ca4RDnLiInJHlpn6jKS75lNYFCI
fJkCPaWWbHtyZJlteyRwqL76CeNhKb3mQG5wirlBGJXTvMDrTRq6IGRBEQTY60CQMN71gNWvHjjA
fU4VlchpbjOBOzeu6YZaEpmNKLMTqnUsAnGnHpTmz72FqEdWpXHxrQc6CVhUYwH0P+Tp+nPEHGuX
q1+jfkmft7C3oOGs/BZbyCwq6pWV3VNtzAnIi6TMHLGrEU4RU/MKZP8bvyVPMd9OHtmJl77u0Cc8
6lz7wIFRT29o2mc7neTktxbJGwBzHGOk5NPayDf3ac81seFFbGmFTF42z20mw3t0QJEJvuRIJsHj
JXKva9t6Y01lfe+XpjKT6nMz00pFUzTTPKnnf5chSsYWCxw7+EprbO6WLdLAfLhTtDUFd3mdqatb
g0Ue04Je5Wy9Tqvj8+EFF9DLqmzNKxoEkBLyJZYnDduncr15ogriOEBS5Bljv/RwBiKbqqWNHVSa
gJzWSl0fIBXzGgf3DE3xHGaBeK6VZ/WRw3FVYAEIq2c8iEuqiBCgl8uWkEJoF4XjZyngu7dMB0Ev
N0c7IDdcL7bHADHVU9tlJLjf8ctH0zDBeIUNzyMlie2iAmoSW1XHCk/JoKbP2nITFoCDcgJhNXvh
+w9io0iZeZHW+T0h96sUjNJYsr7/6uwcYzDZY9b6VrJdzXf2krgJmqTRmwryzVVirBjOYb7DX2YA
wdS3AfjszdMLI44iklzPW2nryIl7KbwSmDKbnsfaELRdPlN4T2B9N9IItcA2WaprlePgsVe73vjM
iEk+ep+NhHSh0jlqyBTq76bOSY8bQim3TboRF0uuzeT+Kc1VCnvEQ/VawQFw2Ih/gtC72CKWY0K6
jO0xaZZWv+eGu8fvXIY/o50RtSJ59NfY6XjBfR+BoFPS/EysMsh5kw8h59UIVe2KoqHlOLl9+ksk
iJ1uGKSdBy3a7mDYttQzr+7hTi9pbgpGixvywDmAsYo9meRLj2E4sQCWIeIUZ82lIAYOUieB+6iT
X9aZxED4WnHbQ7JHT3vqLEmE966ZEyPSpC68GogzSuZ4T7VyPr/JuDC0DHAcdLaCeP9G+umtJRlL
H6YGWsZBMe+nekIdLP935SJx6fPVwtjxbmko4F3OrSLbyNh+H0UrFHXuqSYoejeUf5/T5k9e/6km
RFDQZOtmamEPjeuQnNwYE1sL5GNYlz59TBmBw7tID+U6kX4y47cvUbP3//ooAfmg2mI1qUWkvKyH
fkH9XN50syPE6lM8BkX0gzKJxGZHgXu2T0UWO0CrLTgglSfEx0tlLBV6c3w49xiNIQF5jqez1Oo/
8UHQ+hLCMZ4f2MvLLEQX/2mVm0KbzpuWexIrVvmABlXEL5ik0m7kL7EKpzHn1krbBatQ9QnB3i64
yfHk7i5YbjlMCcx4m5Nl81f6cJWBNSa26hNyLu7o6naQy9VD7swf2QYRKFJ4XyIMFLFIC9sUgHSc
imyf/q1kzIIXOg3r27fJxgj7ZvFI0KDd7uaR9Cw8lMmIukMEcNWRBgxA5sd6NOsX2ICdMFqdR4eo
4DPYYmmkytfubzxSAKXUhqnUd7yiHRtrt61xDQ1VvqhXPE7Cnx3I2wRmh7Evx52jlt28vffreFP2
Mg3lPxYqGh+X4rMZtE8wRDH92fN/16aIQaXBneG1zyhIne8hVU1Twl9ruHQcRL+u1alW9Bn7cXDS
UrTypIsEuxqN72qu0s+FMKac3P/Ov/Q2+w1WmG4RhyPY+q/Z2uLurkP5ql1ZyG0k/APuE7Jwjp8y
KgpUHPcdtZ0EX64q5Fpc0mSHwDBtTxRG3aJVgCSGGv/tz0qfo0MPLkpWZD4iiip1MYljqgnMyPTV
UlTlZPlQlUxhu1z9MEcLioQqBxAAZBDFwj35qqQjAAXMKNuqQyyY2N6zHzL55dzUtluAgMfjwLu3
LYwbwBPFH0dSNzV5MgtDHaDOrk/bD77/j7Cv/XRBRWZUlfACRuamkwb6y3x8Dq1q30rMiISTxelV
OfO98qb+iAb8zhUHwIENuKe8DZeaEYwoSVApW5nYgGlHf+UV1R5VSWSUJb34pu16PvTPt8183zE+
HYuusXR7SPVk5tOrWWaK7mD9BpdbVUAB/OPZFgL8doRbMdiiCGxf4U9N+VVgZj9/IUeV+qCiAIAM
lT1z8PKeIxtTTZpnjSJ1gcX6QD8cBSDDtjZFLurQL4Wh4CNO8sTDVUY8qRM63fLGVHnUH+UWC4uJ
qhQxlhFY9RvjSY1ZdblDkTjcbxeziIUoZNhXhVOYR2CkKX77vB2KI//GBlp4HMUBOCXMAB1tj73B
wXGPTvqHbiH6uA7cPVgM+ETQ7aS2aymW6QiLbuK4cPKkSEFHqEeopPUJdrZnLVjqSbrWGLAgjRwy
3XrsnKdznEQ0SUJwE/IpFfmVrxnvgufQUbuFeo1ky5DbeJA9fxn+MxcQVI9ACR7AV+jtFtSlHn/B
JnL/RMOWCjOg2sIBjgI1VtpkJ3fcS8ZTgnrkKN331CIpZltqV4XeZf8KhHrrc/8AipivF91MNR/D
mS9sS9knCQrnCikoBD+R+bJ2g0v7tN04Hp308EdUeJTpMp8UddLJArD/bV23LzcqTTN+EfNzUkp3
kUdVA8X5aOaJ/0ByGs7kj0wpYUhK3IU7h4SLwr3s7IIWw/aDuS33ycn7cn8+kNYHCiJzqpIdgUXF
ZYRkdH4HuzBAu3dZoowYLtav4bF9TNUH95hJfY7QSq5VYa6e+Tl4UzpBo4l8zMHl+akk2mBnt7/E
hpL8kAVRLegbRnLELQ5Bktoyd2V6HL6aaHA5hDujxECH1iYF6Yt0Q0V2INXcfTnTKiTR8dfx9nuG
t6vnDiMPxbwHWB8YwaChEOUUJeSuJZEK9ifyxIWuOTAvL2ASEYBNTNs2HVn6gexW9sijcOlpVaXC
ig5qylvXp8JGxturXiTjDbPQ9GmtDiDorfNlaPH8e/UeMBnkUfdiHlzIUF1G7BF27jj2AtCANIdW
RiLZfz+Qi4Za00lj+GDr5fN5vCE4LOaXTaovijFdw/A2XeDbdq4FEYAzsOKGyJDo0ve8jmlH6jTj
TyzzUdsRP0ug350/7HGX7Xawbbku+pTPQJUkEvbxM9TcfaouAHDkshdeEx/Xwa7K6GyfBxrRC5nK
6Hbr0IkC2iCQqsO27Btt+GvZ920iNxUaFE7qHh627FZuPHivS2Vz/T/FNrN0N1G8cyqEdei7du1Q
+LyzCfAbH8ZXceG4x/O1bPkJ6I1mEcvlyr79gA10RYpJHfuRuBIboBxV74UzQLDkTz1EtkBEJbXm
be2cOJekx7vJDSfFFEzNfL+ipkYUnNikKizBjsr43Y+qTO1Qk4d1XBzTu1XABT3ZFt7LqAgeyPrc
5tf5Sz1+NFxSDFaqP1NIw3UOfo4yPs9WRL75VWNSYLdXZQh+g4nW8CyYFTlmc9JCNxL8ZuxrBjI2
eDn76G7eafbK/pL5m0NGj7xG5EkCvZT4eyJUAaKpQ1Ngmmau98IZixvdYIMsrmBz/xksE+49nTfH
dhBYoHw4ULT3zU2kLrhIIpoQnAWdJbALdJ+Lpzp53/acFm1bHCgLE5Gt5hRD3UjpgV1vu+ehbAzS
jm/8Gkrd+0R5qw62OKe5eSHuMzXgIqTZuHylu3rxoRiAvf6Ww3lIYQhgOoF0HRfpKbfJDdrMJoOh
Wy0Kv5P3Xoc2ycexhmdEnKDbJ2oVLOx3ztW4IajHmwoVoPnR5KO6DFWJreJOgEfDYNE/SmPUe/yw
JNjSfwKU1n/oLvXRK9q28kyBg4KdvVw8tWmvUGCqgCGKttiZI5nAaJIjuKaHN8IgaVjeAztK2yB8
PSFDp9CigN7i2snIgdv0UwZzfW4t2XFvSQmRsJaFZHFjNbsXWY2wP3Iov1at+zNNle7ot11csRHl
tFLUFubwJyGwU04MtgSu9Rmk0pw6XaIzfNw3Ntg3v4gIsXozDzSBSVdGpMK/9+mVPpaA9LbbnOAf
Q5UZ3fH/c1arIKDQEe4qLQPs9Xtf5N8ZuMC40wRq7mGr+j6+TisDALs7rM+lZEjwqDz402+kmpaf
B1fADvxghK1+qGh4rke1EtNz8RN+B2DYlMBcpmj/21iNWdlIArcO58P3VlhA3df1gq5ID25x3WOn
i5jeiaDE3shKwVpyOScvPJpZyOb49IMGdLPomUyQ0xqL//Zzwvn/E08P3lj91pQPhMetBD2v9vX+
hUCZXLEdYbModQHrF3E6ZHkAVyXdbyHgqg1Iov8gNmKFHc6UoZeItnNQQ1pzPCYVdGhPdYoF9xYt
WUDCWWmfHVIoZRdhQFrW83hjDa1eq1f/8s2JoUMKgMZKnz7GvTsX7ks/kuVs46sOhEAOsygjJ/ts
Sz4U8YJ6DT62kvZqHocFjTlCyRUAJAjZSDWYYn0DqFNyqLsOg7vc8K+j2cbO9boggOy8gUNEwWao
2Ky7K3FPRblyJ+HMYIK7F6b+8yMPbqttJpe8VgR2bpM85EhCAAofLabbuBSGxrfZAyjC333pMHjk
KlbKJFP/gJi+KVXTzHqA58YxXq3wPsrGqZuawDrs6Lkeum7bURPn2K3T7/lKEnUlmlKX5UpsWP9+
e7jUhL2iZcRrDAGQJOkZOeeHGfa6hwwM6QF6BODpw/g1tbX3P0WtotDGO0Et95zJXXIfYJEcqR/R
UsT1gAUnHsEDs8Tjwa2D85g2+yRWqoJd4ecGgANc2vTdhlqB9fk2ezDMfqlzA8+uP9cnIqZpyjRS
7R3bKg02W8G3+3JbddqprAtgD0Qt4P3WDcRfpElhgo81NLU0H5pFM3u1c/ckfK8hP4VsnOohXvKK
RyJYWHR71+poblx2oV8R7bILqmzTBJ4AbgshNh8RUboIPBwRGhgK5ng/wojr7/MK6bGfJQSt3gif
bWPIUjPXofEHAPIAJ/0Pk++qth0UNHdKP/BxGTslIcm+AxvqV4x+xW2o8/KcBKDZp6fvs2cfb83N
gSRJoa8iKZQ/6NaOfIwUJ0+63sUv699BoORwxZjX6RDvQANSVZWrxF/NiacDxx3p82KR3i903h1h
jv4yiLhHuWxGGIKJS0KJEoAo8ta/LholYvtQXQ01DJY218JLHe7Mrw7yRuASL9f1c+HpAgRUWWXN
/9hYzIppUpvXig24pZbZSyzrn3ChVg9gMh3rYwLKTzWIlfqTuS8j2Digz3xsejsyLFeA7UQJzDrk
vwxwiiEjusUQ80G87zBonSAUkH69TId5xOtr+QyfCNCKPFpNLmh4SlT/rf55nrQiw4OYRxobAbbk
shHcggUFOaf2mu1bm+0YntijYTgWvQ/95Arybp0oWRKYMObMiml7Wp7t6oMH8ztTiDpioZODusY+
4luhZZXWiDjinMwdD9H3bq6jle7pkxwpSb+MMfjd+iVh3TYIwd3WepDbA3nWyLItfJhzmFAZCAi8
vAjBnWqvLsMAW0IiMhs8SI3/mrZmPnKTYaDllRQyuexn5O5CtDD8SbASzOS2ysJ37NwgYnSFK9b1
dtlF56vz5r9WPhxzJ/oZO3jyIIDvSehcDSXqUt8iqlih+oPto+cOEO3YAzPfTj6ycj/A377ZZOlb
5mYqEw8T6xcS7RTtbIZWq/RWMRIoc1jhWK+oBEJh4mhG7ciUZwddz781f7PpU/6GixRoRbHGW1sR
Zkh/vcu47osFYIc/hDrs29qNQICG9xSZV/RaisdfArdTqeqGziY+aqYEIBhEFYwPgJx9a30Vf/k6
KrIUqDH0SAYJGHnv9WcuD1+hvOzsiSr4UNJtIml7vc0GUKbbTToxN53nucC7OQxo5pS+syqWBQk5
14dBrh/+HmHNW6n5JJPsytVJtAqRtnM65jEEq8T9WABTqDxw9zKZKSlQuDQ8lIcvm8QLpC4LLnaP
ZIUQcq8BtuNYv+U7pcmPSWRHo5KPVyVxc5lTUSLbdV+LQRGkKAVr1ZPgFg0XAbBOsQrI89zuL2Uf
FrQEWKd/tMKRwZUhqMYl1t8J4wEO5P+zUHQOC8oALvTv/B6OmKdzovHubm5TINxV02fnsDgQor2T
2zF40QEBWYKDhKIItJnyuYuRrXtz3qh0j24JMipopXWcIWHbpikW2VhnL5ATmcABb2OfVKj9HP+a
CegqcnpN2V7EWuMm9l4yWEqdIlagPGXfiELtN9JPr7JQF0jIRwQpGarRvFEaJVWJyqY/6RDQlD/c
Vur8bYlR1AugqPKvewBQn1ZskoCHbm1HR9qth1OusqaVrFrw85rJ7tzAESMVmE1S7pl0ur8jXnQC
oOINi/HHLwqbwY8TH88LPRqkJr2rZPWXwWkfjsBIY8M7wJ1dEyZEuZWHoRo509x6v6eQMT6rbL9S
6369T4JBvHSGZ5FKCP8i6qVHktx5xZR6EOmM8pRmqXrCZDxzMD6zohwxF0tagDrUIpm2v0euxpah
01NpS7Wq/eRYj+VqJfZI9/Q8u0of5QNMJv6cirywgasZVyGIVyiMXkuttuEx4X37DXyjASMRPKCl
7dcp7gXLaRv3XPcuwlrOX5fZlVecn36y+I8qpn3GD98xybEffSo95xe9FkfXuDK62UY3rS6y02ME
Q3dUCR/igPt7qYAz1sJbu1LZeozJjWpySf3stO6hyCTOveFdzVqkL5mgJJ7/4KyjtweIDv6JwbGy
RgYra3FmyShJzsKhlJcprjDRF2tCCyHHFj1JrMtdNQAlNbTkaF7aGBeuG9xx5oaSM1P/gIE42nmK
kKTaPM0A0+93JCh4+Px7K7kBbShUYCe6s/p3ccN4NCgHxzEI++S+X9jm6lVFpWv+lUukP4r/e65w
9ZgLW5MN0EulCfaj087sciJGsQDZq0kQTYdHFtqNdwp6RTyxTiKDlI9cb+fMlFyYSw8MEBWEm201
BTI3wB99v+Kkd6ryznH1Ze+ZvxYGR2znDBXZOX46iLKUiFN4KBNcUcu9YpJ/EpOAFFe+nYNDdKYa
Tzkei8Oi5796qvtl44lTdTscOJwXn5/siXgy8lv0FgZV7++4rb1SXEyvhuNxYwoYSCG+dsNO+bHd
/dRJ/luWyTY3vlPnhit7dk5Zbyi/2DSJj1gtndbs5leQd899DxvuvNFSJ0QBLIJU1a+UMU1y/MHz
t9vpkbfOw0pYvSVO5FFYf5Pjz8VB4LgXStQL3Aag6ljiqg+4+UVKv7k07Q1bmwrSH34xRnE5QJZU
Bxjh0djXtOo7cCESC1clga3CDA39IroRZYrRsEPOqF4/K9gUxDAzZERJnbPK8tSYlCUQAV4ZMUQ4
CnnQKRrmxw+v43sDg0f1sIeIMEVY1UcnT28sJB2M8EcM/zZIiHBfD3wdztsRuie01aM3uIu/ovuQ
DU42zEWWH40w9RjEEaqg/bNI2gN0bpJT0q5e3BbUErRgX9xC1bK3CnpXDQHwJzokLNcbZmq4/gwK
KoTD6+2Z+C+u0UyVE8y5pberr48PrSqbz4o8CHYf9mDDI9ylQe6N6xWAnhPLWaWitAtd40MTBEuD
vrH7zG7JHLSTuFOXO72NcNS+8oGIKUhFmksIGDXEHSyR0MfAdOP1dFloED8HW2oTLcxI5fyriamh
fmLKR8v1AjuDkkr7faRhm2afQTrrXPciBY+h06HPGyA4hbl4p9RzlNKBqBWJ+rKaPmYT83KCwfyf
UZFh646Rifkwl0YiTVM9TgCfWYCWHQS+MwNQsCDcZG2bhExmA3+kYx6IWR4/FjHm6N0qrOzFO33D
3xRufli7YT8yVgUCc0E9+yvUtpqpiwolZcyWmBvimPclSInQ54Dckar3XGkx7qbfXBAqYmpsU5Ey
skbU2v0LT6eSgwjAczOd3DnDcga+4A2NOe3wJ6V9G9Z8Cusjbq+c0oucBaNuUYI7lH6+hYe6sguS
/bLcX913v5eji89DeIwJQApIM+lOYFBw2UE0CyAiz98DHQoqL9u4jMpGzduUjHOXxdQRccy1VA7Z
q+s5Nvq7OcK78C04HUjg6ZYU9koF6XwOe/ynx6AKd5MMxrvnOeKqFm2jjDLZFaZgVAF1i1F/1bL7
CX6n7mE9mrXcqNrGdITDN5+XtzYq2J0dlA4XzvJhVq5Oh/gpbQOKc5bpahFbjdlTDfCDSskrmEf8
K4A8gBtYoiey9s9ZiQly3IspwwGPAPASrCnZ3wG9plaiIZRGjkFRCqqMnoezNl33BXCI4HrLJ9SD
G1PLvDu+ZZa5kt1Z6nuytK4+QTUQefdsCYk/HfGuyVPZuZvHVC32K9LMeI8vaoQ3X5CmXinfAWM8
TCPQVo9FvWdqsfxmbWaiYi3Kt0AYj9VFQjdzVmtEhRyTMVMIZy0Rv6unUPAb+V+7xQv6wHE3i/JK
DL+C00kqGpWRdd5bhLyy6bbX7KsGLjOkK34+IhFCvoawMaGndvQIqwvGLzTZB1M7I9kt3uW3mIEb
f64woGMPLi22hBbbgAyR+JipHsJZFqCB5xqv5MZnI2F9EJw2um80l1JYa5yZuVEFCgyV9JDqRErH
YZbToY/Q8m3bhJBE38xtH3Ag5s+A3kcQLMOXX5mhFABNe1J718UcnGwW8NqpUfFCp0mFZY+Dedld
HnEYjNP7bDHxstdggAthrkr0ykkVD18rGY78CXnKWSsF8S1QsiNL6e9GDeBlSW7KwUR94aMALlkd
dgycqa3c7uSXiYCryEzaxTB489KtNmkY5ZXJ2rJHQOa5o3ney8RCzJA0XDBkUIfxM6NFH/+arFOv
CF6AhYnSo2o1AvCa+Idt6WetnNNfOHWQYXDmsQJzfvjZROEUU9Cg2Fz+FRTteJ8tFL4RVIAnifmF
R+92fzQ+zLG2HrvmMNZSCahGl0TrKA4IXHvWtVcYwurbQBoNO+bF2VRWHEsdjNm+QrjwzgrmLd9T
FOXlf2FbcHSjWfHOQELG2hV9wWhNAXopasZ5s0vNIdubtdWLFMHPxtjmdnVkG9SED6f8t7uqCieQ
90rtCd+k+JfHuWIDXeTyHW1MiFv7yVdy49dj7etJyiuTN3Je54O4XRHGo259w7/tyQmrwaEZ9PfN
+C3JYvrIS+XXpArNSm0E6G/IvV6ekRbJybSTCoFU7DiK/vH4mPTl64Pk6mjMVKO3a6XkWBtUM6gB
Lec3XTmC1neBIrtQyiOJjMw29+4P/U0RRLQ+USSKoUfhRHF0uJ62T92pvuBsu0BdOjbAVTdpWmMW
z6Lzr2mSr+/Uk8s5YJHCMsYRVXk5CzdJetR6CP9W2Iw+iDqcWAdeZnjx5Vu//QHSpWcxiSKw7NQX
nE+cuBla7AJvTRoo9FePXWdeqoohuiEFd+P9X+r4VKv0XwEuQ8wW2x3bVVt9/ow4wVyY1GT4bZuJ
TElGUuFBXgQS/FcFQREh/V+S4lYfT39XFAMze+CTG46mhZaFXZuPLwh2EnLIW2tN4b2nrooJ9Ofg
mu3C0RVylwWFOx4XrL62qZ03VlYWQmjklJRZbcd4yepPrPhJELQZZpTW4VpZ7b1ifSh7uGIIkYK7
zHivkKtUMys7nqp2sEqNq7apulwpedpWOMXTf6FHdOMEsf59/ZL8ErkLPJgW050vqAPbwETrTIWf
F6hgQmdoniY8DgHJfJ/br0ZJBV91rJqG2kIVTm7S770SKZhAUolAV0LbKFmC9wPjbNnIDbmYUlu+
VuqtU1vZ8s3HOzBP+1AHdFYjN22PkmqNP2XM63JyMlKub5qkPsiZ6ZX568RlEx1FNVzNzhnIpG9z
/aPdwGJlfMZtrTyJmPX0SKnbHPRMMSfxsl7OLJPa1oRb+JFsUMAX/05+3bz4RnLjvGMPzpMVtsUx
CZG47dR0TANksjfKa53G77LPEr5k8HMxnvoxFbHXRYUVja41sXLsrPnLsEmtWvYKjd659zurIQJV
LPd4K8lmrj3Y7vtAjET/nRS4RXTn0I5f52INh6NrCuGjAx2KGPXK7+ZCY0Gec/AeBMFqGilUZVsZ
GsWQpYuBURIBxEc5otEXQ1DmzzCrF43dkbFf5e77zgMG4VUzlhefV2KND0e8j5cPB9FzJuzmsURp
pNjs4xvhhTe4mGV923WKwqKSU9W3biU5/KeAG0PsaliwTntl/TaOm7c4HuWNLELAaw/YoM+cnpu5
Ynqqwp3RQXb/qhPStzCXhZO/of8rCs2jwN6bUmG5de9DWPfK5Lw4Nu2f/+Oc6pLUQ4E7FQtgaeBi
+lNWshvL11OsO7AATO7H8p7BPIRZjKFdeKa/tvymsO85s2gqFXz8RtqKP2Rwh+v7GVtevv414x2F
K8hPaWEhiJLl9vAsV9b+7iTbU8NRIe0NuK1vImwHmF2YK2tc0w9AvnwQJIJMuSYZa2Pxp/TuTM6J
2e5ySmV1mh77IffX213iHBfrkczVT2IAKj9Phmlx8ouglDIPCJpF4GHg5OCYh8Fo2j2wIsPSvBRx
Si0fUILTwwUa3Kk3UGvV2Sfk8TaNY1nnfogGOwv49na7Ya+rlqbwvKMQP38/eOkyGX82DL9xw/bX
WD8xPVM08KxwfdqzdpOp7TUoaKqQcAOAEnLWVd1cm+Fbj19ZRfkwaLaRlUK5AXJMeY1w4l3RBpIb
n7O2wCBhvr5CXBAoY2bF+HriSTC3TPQDNw2xAHbiWwdERqSHDWN/N1yuvubP5XnBvXIh2Zl7es/P
mPmxvy7fzHP8ZA66ZbX5EZDGfP2s0Ru+e4+QjUiZzkHlfmqVCishnwya4K7jSIcztLP+GBQE2x1P
8rx6R1cOgyb/yUWr+H3n/Pp4tlaX3fhP+YD7PMFffKrhtr7IJsWVczQij+vSfPWasysa0491J2oj
217gA0aEcYY4paK0tNoay/WSm3KrBvOLvqq/sIJpOVghQf5GOw9X8toMoqjdy8pEWGad6y2Pp/wK
XvdjIshUg+rMaAs9+x23uypy2u5FX50pWpHukdvojgHZmnoulTyGpJlsA7hz9mK3seqHH0R9aBbx
/kZJl67SD9X6BQ5vXWWWmVGEDz3vfGXOEK/YjsSeTN7vG/2fqZP4BjInT8s70DaFuBTmSVOd5FVb
+G9F29iI8J6wvCocwMjswDr6SPl8UvEuH3fXke93BKlJXky3ja5FCAaPKiKCMpWW9kp1S+r2F2tI
UY2vqZKneEhrwesg4bCFyOhjerRnfa5s2tU26mwDN9I9ON1FO5Cdn4FxhCSH8dRssayclr4pz1Mh
SnOeeW54cu6tCpGRJJQYpAHhItGJYHfFzJJZxxz/Pi/1WvCg544MP16IcWUdn8oI4MRGs9GOsnr3
VCB1gn4yTv6I7DM2LYejaA5DFwAVbPJChUriI9K8vOvqIAa2kOFahaMtSzmqNOhJ+AqIsmnQbAHR
8cDvXrVrNKRtZWLdWUDrKKMpW95P1eiggvTNj6uHmOCFwMsws9TKhUDaZd8MNnFKSCQJ5czK5G9O
7JAIpf2ux5/J2kl2MfufQZ2zrqHzKRPpGKi7muJle88mbeEj/oXgs8yOcxcnc0NPjEXfNB44T5d4
dzwetH5QpQqMmU9AAh0s+LVM1amqF2Z4Fp/hsg5H0vZXOAO/n4rf2KtvloKFNDm4MdLmmIGaFN3H
RJLJU1ewym0IXKc7wngHo6ydxtqQpw/kmjRQ07u2D2NsdpCvwUU3/cdTuAur9IxcrjN3Gj4cv2Jl
JEdvYsnMjS/Eyim8xES5dVuUN5ntuzTsFV9xFYj8rD1VZPM8W5hbMqqTpeKiUHa3vTsqYtX9VO/q
HESd0F0+HUuXeFCQK2rNS+mGJSiMSvX35PjMIwU4LFR9S9AspDiGtUYjEfnIuQfvkggl12eOoIyW
B9aiyvN5mk/Hqd23faYUU9Tuk3v8GA3TzudE00VXIAs9QZmWUr6Delh8xbZRZbOo2bADYR+w+jvC
7vMnO4VtRRrvsnEHjiuffyNR4LbEJK8n3pDvYzO3gQylVHuMWjXBXr+q0dv79bs5JVHJy2fKfz6+
2LYNf0HnkQ2W4rT29gIhZDXYPlxvAUslERryta1/WA9PHZDZLN4gh+pG3w83QKDs/izZ5nn5bF9H
sXSwqm9WKi5nYzQOva+yrsQ6waQlQ/UgvJFHVKBW29WYuhPRBbuRlfGIelpxhO0Y1PnOOMUf+pkt
5ghAaJvCjNHt2uLR4GIEqJ89iN8dR+/g3yLaRBCmyZMBCKHXpG9yDAouhdkgd1HBhZ14Hf5C45HE
FzcHt8y/45+Rb7xQzem7N1KY7oGipDqHNZ8uyolZVXH/5ZpemmmQrUKkCB1NfjZA2ifmBC7X23Pw
/mfuu5A5PLwXGcnLnI929iTy0WU6mWkoWZuzUSKzg8oAf/iv0hMq1uWgBcKEzetcFPUj46B4EmLb
H/ZR+4RM4IUEPu5LnbTmdmSGJ+d9N/9Ic4X9voDCwrc/xjrOjiDj67IvWFeFWoYlR1GAOtdSUbgS
LzQa1cSfi6YbMUL5vRZDwEZSZSKI6MuFA3bvb/QOD8s1GU6bxnUYwcx/feRLP6G7nASIR++dcsIL
b3FWsEu4guEdXMJpocNcj4jdb9Hqorcf9jtk+ufwbUWaBOPISWzINAcTNlKGzvLUz4jc9oImwU2Z
B2r7r8BkCXYs4tJSVA2a1k/uXyPZGuDIkM7Yj3lIzpN5MKgxzSDyyubvfr5yaC2Nv/ju3aY/WUrz
lnzBO0NRm7OKLaHI370a0xj1K3H732yynqh/mT3l7Rccdo1wjeVS5B2E5jz2xYdjuvQRpRx7M/St
3PPjhB+BR2FhOmbFJ+zIE24FUxJVe7L//w+NrUrOERYSESK5/ZRrKf5Rx9vyxIgoMPMrCiJhhVgE
GJfHBL2FR9zUha9jEBS43mXtR6eJZ/alkfX+2ovqGMxs7E1rfVlazz3wcw6+0RjLXDS+vS8Un/EC
oD8Bjg4yhnIWiTWGCm3AqV9+1prIDOuaoVBjo1ZG+SpAuJ2WEvQcd+sF+ZRqAboTUm79AufeUfB7
99b2YJHXXn6L6aZFP0F5+Z4Rzll1NOQ17mI5fiaJP9I1WgKLQDb56qifNpw7jHJ7e09goqOmlxdh
tHXYMrk/OdC9EGINR1Q/ucHKCoNExQhfd5DlrcyIUs/NlyjtHxP51XsdfpExVG2tz7KhVtHE6LcM
Oyf0LAFf93/KKJHU6kfKzRyz+jnrCbgneqT789xpwhKE5RvZ41brNGFVK8FT+1U5QougT2zKonlt
UDYdFxtigO5sUIKcZZBln8j6mgrNvXqH/+RL2PtN1hbecxbb0hm9+SNKgBimvOFIk3vCOaPN2wjO
pwtq1N6OvK0PqwjDUxGAT+ROJp3CPMsDc1ECl0NB3kvJs+D2wgpSLd4kHzKIShLTLXoSH6Ko58Pm
bVT2rLptXy3kw0lc+XkkXwYI6Q2ndtsvHzQgZz1LXXf4S+zrFJAb7YglrGeujMfX67cnZTnHukGL
NqmkSi4MBA8NOzXIgSGgtCTb9BiaLdLfeCCX08zQ/YM3R2jOkciRxYC6zOwhIJZ+CZj1Rb9+4P+y
t+6J79jFg1G2BvOvNG8YXQ7ORHrS707AvM0G7vuAU8NklH9YuOQ+6lKuD5tlnkqQXNGTgdW/kJqk
PfcOgkLs8zFQlXv1kcunPQ8djtwdAbJfhlZcos6uLIadJOa+RMwDyRCnLaihwSCxUZ/b9QbqYXUL
4Uw+MNHTfpP97i01/8NJJeDSeLwpffzXdLS1vpPwlag6Xz6oFj19CoHzyBQ1GGDLjxEhO7Vyxtlm
OSzpcZ/uu2BcxwCNhCRUCDs4TNAwwLmFH0Q2Uh5z6nR3PA7/X0PrVVv4n/ecR2NKxZ8zxbjRYheF
6QVfKcATc21e2L8pZkXEI+qDVrexqqSTk7+aY8NQE1n530ojo5gMUlaHXuu3wEBJlbANSt5r0T7O
tg/AT0M/hrov7PfvSTM97/Jw2mGymx7nFnygBeVvSb0B7aA7Vx5coJhuNlvpC8Le0PHslAUjGf++
FvtSxiMiA0NNoL69WRh+s94ea+BgjFavKSnW1i49wa9KzUKi6kokUQxXNstkHteV5sE9ikrAq8gJ
JOIMyZvj+EpLK+44s5+OUXjpphNs/uHKt9h6amJW7Ill8NCiClWQDLQNFaA1pxwnplRsosr4W/Hw
RhwtojEtscxpG8vw0+T3LQBlLwp4pPUftZ5ZWVjDBCVv+3mPDdmUUdYmCZdam7USy+/1AEZUN1iu
ZEZtSHcWHdG64wHoPV1c8nLH34eU0R4z/UpLZcVE/+JIL8O02rs1kO9fwx1DNjEaQ0xPJ1VhOgN3
HFgCrGscNDuAPbDHM99bh4PGssXHUktjGWuFpZrB+vG9HaLPtMeI1PU+kTAgook42pm7E4AEi+4W
HDsla3CXw1R6QxUq0o8Z/x824VVwp+XBtNOWxKN2fR/ZJUiUyoOHYrAxfmlppZZt94YQrJeObiEl
qFe/1V1hV/0UK/XVkQIpaGuSY+quQd9YbXmMytQaMRpIFJoChKhjpzPAFsUqTGBTc9YqWWQ2QyNZ
lQiVGWU/IHGpan9CFhrX63RbT0/334pIihGAtcGEv+7Zf0gf9q9joJ/RPiV/nxaP0X8NlPMwLaS9
gQ9XRuOIXiBUdEplBFiLE6wvbEduGpKzfxaFbaCCvfZXF8Hverg6JeJi/PbO1UD0ClSSlcDTNgu/
KCChfnKRuJq7NbqaTV/N/zLYF6Mz7w7ywyqRlyIQMav57ZZqiUKjLEkCgIgmDWstzOl0mJSIBU3z
PCfCBvCgTEQ88CS24RKoHbaFMGr7KGBysCR5+B3eposTkhqRcAUwIymMiezbP4B1zJCkkwaQL/5f
tCOldfMJgvhiSDEPkGe3w/4Q/OGpuaS2DuaHW1Gcb20BIdr5KLwxMfUq2+Xg/rlOpLPESMfj90Y5
seSnXc4qSagNKKHIrCBcdLfUEAjMteKzyQ5wXJJ51T7xvuEwnE0mUyXOMrgNaxeFXeLtl+I9tZ9r
bYBlilylGN+fiuLBCmZjTNMHZdDYavR67R2XHS6/7zxPHrzxkjXiaVvITSHJ8s+912J+A81UsuuA
iLV7vbyE571mCuiTiONGGPQLKSKeFQg43EkSwrzElrYTg/YshmtowqLSA0oHK/zSlM6JCPmwmJBd
rBP4VHfTGiYGOPbrcyXx8Ze1rdBuUcetIGeecbuAWMv0T8Gh0na6z3InBaVX5oDCHIebpm5cpYvb
MGTkM2bA68cRzC/4mN47y6s0f0uX5ywd/bBQgSTkSqdMLrAiocz6bjkkORwei33YBOh0dTddHjk+
BgcJ9wJdT2dQ2oOO2Uhi3yf0rjYDDXG9ef6Vav5iEP5IgQ54sy9FzSJ8+VUiaXFBMXRVOlnKBexo
NelGWfgRoy5E2E+Lwy0ewV46kQlHQnkIjTW63jitmEvs5Z11wSWZGeBuO4G35fyPubsOcnWZnC9E
RSN5/PcIqFlYPIxNIPESXxJ638gF/Qnt4JbgVGyGTY5be1WZPIXiGS9Ymv6eLi2Cw9/UP7NNkcwi
ELcMcAhrmaqsX9HnNV/wLiVJBvz3q3YSDsfNQpAeMRTjM/hi8Lb7plPgjfkfERlZ1Z+aNm5PA+P7
ZTSHuH5+wSJXI1O7RGkfV5n3QEAP/s7TKDq557aoGgj2yeAo7+Vp3vq+9Gb233eCejVerbvqlNA1
HOeuDb42mpVedib7A+xN+s8bL82m2lHb6LHTEgZUlr/UlTGpDbejmCxYQuaGpTjdBQ2SBq/c2t5n
cdoiwBDYyun2rGVAcYEmpR0btPC66pZLRD2KQwpkjXXTQfu3dUbGmIKK5x0lyw3GVr+Mwqxh65DN
6vKBjROb47p4h5FXn6yfHjwfKxEiB/Bd7ck7OkOtCgHQ66jIzR5H/stJz77kkVcO1nQtVHNZqcmN
vGkW4W3C9lhsZiMMMGUPSIFK6GfaFuvC71PgjN4mokCN041Xa1ccX8Fpto/eaLYJetuVk5RbW22C
ob8zwGTPdBU397Iz6YdDwM6E4XpN3G58C7eJ1junDm9o4JHWJkx8bnL8YhOy7Q7fneas3NZ+V8tb
OvRHDYAgvwRvv4uz8XEtFKP/DgtI+HwQbnsc0dEd4gTe6Cpy90GXRcyBWAiOnuztQM/07upNOZ4s
FVNvlFZfUbzWf4f42poCUOynvgajTQEqz7W8rdpJ9qT+cva5OjPyWGDcSIyAkoFO5qy0zLJ4JKUV
ODiJ74wuxn9zTQM3Ne7VhpEicJqB05AYx1VBHcqJ5uZbIAUEJhZXnK98fgSGco/N9zb39n2469U1
BAxtJFIm3j1KxArN7HK8zAFyPazeAqRT+cFTGRFGkm2/NmPe6p2lK5POhMwmC9SdLWzWwsgmcDMt
tuNqD1ZeAtlvEYScfnZQUaMJyrAqEly+QjXMEeVkmBwTGU6aOLVftrLkY2khDcPzYUArLQemNjd1
VKwViLgMZxruYPq/aFLraB5G2oNqyYFa+l8crQIbfpFq/jJ9pbakpZMcKsE0hKKMyHKQMjmQgxr+
yiyZzNogvygR1xrDCwZXIOX6/AiOqI0kv9tBFIOf47KqaVh2T0zBIl4drAa22zz8vwrHDX1yrBB1
vP7upfdD3KhrWFsk9CCchUXsOuzFQNRcM13JATqBMUODAolJWo8LxsATLFpxA3/XlTqEcIc9OydL
FidVoQBqPUrRfZDBBXXw3PqvoKCbnMI9DmEzKXqVZ/KE4PYH3evjBrwGrXWQf7fwDOV9YGXy8WFR
JEYoofQvsYEMI5KtlBxxeFSkWBIb0UrYfeqTnkT2MR1/vKGygfFutNHzeAhGGeP4pAGbSuYNzmeN
eRiy3EN8w5enBYY7ND6dG/FY62F7Z6u+vZR3M9AXvux+qETRpsQ+wGpLGpNFv3N1Zu5BqyzT5p8O
lPHEEXjJBhbInX7yWw6CPRtjvjSFrGEm32oQ4GbcxA3bEeqHCc7AEGUJk2o9lTR6bP2U/B4iv0+j
DYVrLmK12+3c6QF4ATKYmdCsOmVXxcqi5XJqdDHMa2eOQep5FPB2f3bjINg7PC33u170zj2FN8ME
QnkrFvXj1ZtAtMC2q78CqAGtudm2iKPo6iIDs6fVFCVx6iqIUbAB4TTeRrx1x5Opx1MhVGOrLrMT
zgLnMIDZ4eNLEgAFIt6flQCjubnxBhRrg396SjJ/xR8MlKyBOovCEVFtPgq2tbThMi36+gIS5oDw
3+WdNfMKYiaq8YnQUkWyJoWXBj+0nshordLByJDuISApEkYkUvjDhUqloyA1AdjO4D1iOS6m9qQV
Q0aSEVoemTMCfm+dCpVqFLuKdJKtVtwm7pysB69jLLWR7HBxTmAvyilwSvniBxgubDkvsLbnyvnA
1CaVu7BbP/8AhFhcqmuCxo1p05AAReChUSS+QrpFBwdTjCt9RECPIu6HWhaMJ9OPU71SwsJym3Pf
Kfe4szGP1Tkkb57IBMdJkj28bcUzutsbGMKu5AdPcJsQTZ9Hkv74HaYVWgUXlT1CwnKb3s5ht8mS
A6r4eEMrY6fLBz8s+V6mq0IZDJj7as3yB5KQkkqUEWXSinmwy4r26oRozl/jMGP4u8xqWXU+MuAL
dB4Fvn5tAZzvXTlsKRsCXgY6+TTQlRKdx1TmZWpqgvaUsvV1ilfI9Pw+rRwtmmk+oZjwW/5KskZ4
SReePG38B4dRB/9fsB+uUmWmu17iRg7zF6raYXzNvzll4AJXYap4bc7Phb0BTsnBpUk/4LDkVwbj
Z1/vkjLsS3Jgc1iEs0cb8X8cL5kD8o2zwK+Wl4ZSXKlRJJW6fULmoFxW5tv0+LzAilp/H4gJaXDa
yU4HthNi9Bz0JCOEcEqH254xrHoLlf1fhUveuks4GCEeG6SMheRRdDA0qnlcYA/GYexlbJ3YTxgs
HbjbrVJA/ueVesS8c/oVk7aEsaJ42J89vwmBuebtg30YivNK1BqYEfGo/bWAkGVBh1bJ7DThZ7KR
xqlxSLVklmdnGZe5ohEY0U6DgmcTQWlvZ9P5Kst6xnFNBZDjHjxNgITj2ptQy/TknCzgCa5SqeCW
GgMDm63Pd9KWm/XP+RV3l1Eq5mUM2sDe5d628vkGNDEpN6j35o15EpLgnkulUW4NcQ22vO0iFmaP
27ClBBDPc7Wirjp67gtI8aqRf+dBaXXePr2xWNQAY5J6xWH55wMaXy6i5oYCIV5BxrYzqTpv6GJf
rtmVDsiFQKejy97/y6yHA7ByfU9DK3iZC9TurpFOreqMAF/8sivygq7pW4FYfXvf87A2qBsxOLad
j/RTiXken8PHvNRO1nNVjxwU0V6sV+ko/xig30BeqgpRg/0lvN5BAGXtf/M41YWkM90h97nK3skH
zpUidTkH4ykpUN3TY2b0EZaeZyl+eAVhqGMZH8uLZVan/Yd/5t1QpJLW5A4C6t0KXRXvuOTGF45Q
ciL2b56jxh8vnQOoDhzgb8YiDAVVI538p9+PEcdEE1FvDvAomdYNvXotQMyzt0bTi84evzr1HP7N
Mv5IPhko2CQaPq21H+yPE+Gk/fpcs+sxym4PUKWY1j8phtqIl0EG8WcJ31FwGFCpSkCELgMYYV05
VKFPQS9wI2QdpbiufJMy3yPbyPL5UWWUOB9ewVa5D4hEQK3RVj36wzdkOm6EO+ypX/kG2WoSI+WA
IGd3kcenCXzaLUn5rlwcbmc3vuOLpTk6CCicFi0pZL76eQ8nI7betXZofeunV+TZSNq0PJWI0mIy
Lh3VoEF3ggU4Mi00r6mFd6QZ0bJafkefk4dkcnfFXzBIXJZgo51KMEfTiLN6yt4K27YL7ZyuoGND
ZjFHh5r8vvo1oyfr66BrRQavoWwFkz0PJLE9Y5HJuJ5tWvbF6icBLDCL0m1AsDHEp4g42XMJw/NU
XBhPD2LjE+veGEg7vaTk9SjGPcya7ifn3CO5l4moZ4P2WxFwRxNanQPJOhryMlEeCPXX3khO7TwT
eMg0Adt8n6w/iSlT4KWpJj07pYdX26t9VXVtpojo3h5eFhw4w+8aEQ2X5eo3jGV1PcKYIetZ2YVJ
f4mZIPLEiI/cBKLGpOae+NzEmRIGuzwW3FkaywOLJCgEMA1QwskiPH2Rg/H7anDgrOwY3BCarZgd
iTFqEfL/3+2yuHC9EXPxkFi8De+HMp49fOsjghD2xzs2eB2MQmTgPn402JKcSEEEN0qE5dv9YpDd
k4kS7PG5HaHbRNGigewka2lcts/cRbJJ5IDHUQ69kcA98s1iZB2KoI8iZDtggnI8PAP5TjEKAXcT
n0b1Qak5yMTXstSqgRB5EaE3ymQjB9YraFUzDDgCxMwYHSNDOXnMBgk4lR4r/VILc0IMajVnqU0n
Qy+2Rz6ixr7ljr0ARu61LZSlE7NLbRh+c0oMiQSPW50rjFZiutEyIvM/rLc6Yyri8380LcTPbhxp
rV794Lp91icVyraKO/C4qyNz5O9yPuN0DwCNWejEjEpnlX9sjTcs6AlNsItKOyF9nv2hBe1VySzO
1RkAVTmAVPRkNO5K2OPuo11FJcPWBEI6MVpOqLgs9VA8fptwWNFe03kZ5Nhu2QG6J0sa3OZFw1/z
joGzwX8G0QbqML8ORuoRZ54zTa05ZEEe/ap7nUTmzlbjbzVR7y58qWLW+fzdEp99fNyNs6VwesZM
DP2o4N97YCw+qqTJKzIAHHSc5njXLOHd4E2jn9QHIxw8fRkO+q0+HtEf4KFJ4HiZgOJoSX8ZJZiZ
3+BvPcCRCQgxA+994sCkx36EYy2cgJ4QmcIns7scGLShB3IiR3WBqllZokHoB8gX1yT+U6LeiGrP
ZQime5M/J46kRGXiXY+zykpSNucb12Zg3ZxQmXIt2w9WAFe8XwQIm7305IGPgQOKcxbkuPQpPtUj
r/M9SrXQIldgDcWevOUfzpxbAI2Hnuc5S1kPkfuKVh/CkNvs3Kk091N+EAg9JgKe4GFCO1qFXShP
JKsMPUGZrfkEfYxQ/5xdcJzo7/c7AJtV3rLbNtEQLeYdKl8RbJVVsywWZDsxPC6ClO+pfgnNytwy
szU85Ve5kNP16rLdblflaHxbQVay5RmWS7b5QxeYilJFgAftdLU394d1TuBsv96KYo/Xyoti3py2
7z7hY/yd94TJfzpeyRFsrAFs4cW2wnnZfyp7E1DDLU7VBAedYEBPNhyLM83eXCM4tIaAYp/TU0b+
Qagj9xeWBae0diZ/7LyZwB1u4xBlC3loHqIJHE4bkU0xDxGWQMnlDJWxNsr3QTXMeKqix6vvv9UP
NBFqBVzvtLgRBPQFZVeqReYWNk7JkprOuqqMVF0GaOttzcoM90ltIRpirHIeqAQyMYtCIlj3vUnk
oaStsktYu6U8l1QXhDwnNmj81lDs7KNMVozbMw14zEVKYd3HKkermQzWZ5HHRoI2oB2+G9RYtSR8
sSK/sC45J92Rgf1EZ0L2khH7M1mdHkj7HbRUBQMgDIi1x8v/jvpi9U9oy7Ra6m3GpTZ2WbA7OkaF
b5SxoN5et3V8NY+KLk2U3LsB+g8dVmBpB1u8wiCNSb6OynU61ML91hZQ84LvtNQuLCBgXQX7kQuE
/yedrUECz+QBfz2eY55DxmHOLDRBqL9GQudr0C8g2qGvVXwfxqv6lyUj2R8b2yxXY6K3xeR/vj7K
6D30MWdchPaEE51Bx3hKdPSnBwd2CFxBlTIQDFEHFwkPE5aUj+qb0mPdn2a9rXJjuekLFzSuLf5I
edwGmNuXf9uuQ1hkOIWP9HhIAkl60hn0DKaAwfHkEntnAs/bFBPUow621PZ4ugYRYvXKC1wdomTY
DrsKgg9iEaC2OP2NGXxfaN0bCp/LOwYADYBWJeFIBQKTpfOnDz8+xKgUliCIIa9DNEcsQx/z4vwN
E7y+iCz7cwMFDtpluEGMOi61Ji/aCtKH0Xt15nAVxDhBqLz5psywF1XlfDqT/cX6eHXcWNj27oAW
xbjKFD8AwHqlZvNOU8vvTKrN0nc4ZI6k4smrH6rr0IoKax9fkvAY0+Bb7pcQt+eGKZT8CLoqGqSN
4Pqi3RB7DytxC6PCy5JWYkJw4yB9vARYX6CCRoPsUnprnINZ5EFkPcwgor6e9GUU1S5aySJ6f2y0
tmEqD2Z8ot/nFh8JkwvIjmQSIVO2lS6Q+0RgCA4zr7CnHFziYuLvAhJvwwIJMmZC3Sf0qIDHrjiW
HyQQ/NDYH+Su4BrvEUEJofF/5hpYmfmYH+qr/LRzJgWrbKvxQcSVPnYQ7HyiOkG8JPlex9pDa0XP
yytui3yUPLJsktZ+wMD0Qm0uilzFLpGIN3dzkRv2R+2M1R5nhGvPdLsF3mDGrm1IMJGD5hUASZX6
krfhtwcMKIxAxYNeydRkW8X8+/sIdVLLQqdFsIL8TLYvKj/9gV2JuhNl006g3zm7nHxXKJEe+BEX
sDTDra/jGRJ9pxM9PYs1Z/yzVGLKwkbcwn4jYHAzLGIiVbCb57CeGZblQxw3QkZELctj8C27Te1+
j0iNQ7Sr8hOssObd7RNg65/49vJX7QrsCHjGU6KDbY28gILIP8cjlOqIQ/UVK29WYyuSLCRTsKaa
8OGtMrriqIoMR8AMouSaP7c/VMmtuBCPMkLDaVdt/8I5O7SnuXEqWhAlYLyt7kSJW6I6ehnsy/Vh
dopo9PV0Irpz+s8ho/hgja0c5OHUj95X6hAKjSAzbq/xA1Fhsd9FX/JqsngKrRzwfi39WqN+D/3o
FF+Z7Kt3bHMnYZElH1sivptiU5kllTVwpal7rrbxBKbBbMgJUF0KI8TGdlnsU6VQyGMNaCoK+lQW
d4wKWbYOZwvUHtkMAPA5i3w/XMGAI1i4b1gjTIaIInB7pKg5J+QSccojndlTLfC2TKUFNK9e2d83
XP9mhywhba/wdKMIRvST9z4H/WW1WRgioEMa7C2tbCf1c/g7aaalD/U/6n7qPawjdbh1knUQw92G
7f9uCakSYuMkm8zjDznvB99NRHpPV/kAbRLflD91zhzrsxD1SFN9WHUzrNyAh+z5MNkI95+Ss6Ca
B92Yf6/ksZasXH4NyvRewBm/imq5qvRBCq/FqZmkK5h80xAvhlRMyrBIdougfo3t0UkOHuwBJLe7
u3m1ToLDpQjdMM+ks430Wsddp7hnfV1/gel6m57pYWH2IQwBDht5G0LSCVfxnOO7vL67J5Xwh65S
6KNePYRqu7GSVKOztFfbLIrcC1hQ6O23cf4FEDCVlwvmCjH6OdOf2oBsAPKZf0YpgGvjj+ElsbFj
e9hV2vEsI5i2q+/MlziAOm5TrVJ1Bj6QPAzSijdEtkHBlWHsVCtvHdadJacQ6W/X40kuvvfh0oaC
S0ZjNjhTjyP3KZeSVVwZXMYmd4I1IeDTsySSJ6Ws+Q1IAWo/jv5SI5dog3DeoWe4FnKin1IDNSvs
Vz1ZH3g1F33tZ5wK7Dr/bDGGRf8Dk+juM5PseeZEirMGc9F5tAWUEvXtKirPYjzFNxyBz5oJLyeO
8HdVwzWfwt+1KHWvCMXClzgqAUs1wTjoKfn7fncomfHmjhuppoRUGfioaoWPLpmw/aQTG8oYpVDe
z6LBnpzK6VWAih4hyHbetY9snaJ3WXi29uFk/HD8MVJQnsOwHTuLD7XUY5y/CLk+5/iYVrVhuCad
9mDfEQDD9ZorvwTglMHM5CVgVpSkvQtlL3iFVfoY2ZhGh/CqJVh65qsizqznyFfZMz1xEH3lvBVj
qGwAH+sMDh9OfLrb/pInXMFrMnTWMP6kBIsNTTnO9oMFlb/Nl07DGMl1eulAq50sq4L2MWySmXbw
XPYQC5++REUbAH4P9w7+57TcULhr38YZ1y74rp/cWnfbXg6GTvIUIo9UCy3MDlYmQVa9x4wbRCqA
xGw/UyTmu65RL00Vn1zuztkatSA9hGuRFkHfcn7TMcAgPqUv0D/a/4DFSgqhzpOQoJX4l4ubrts8
EFor8AICcvjURrj4dAQS3IpHTMAJQHsq7VtbkH2CHI2iZwxcEcI0T3KGWuFxYnTaqf2eDsTlhKK9
2iweARDMF4eFq3jouz2+3ybYVK4rNDgNVXyy1e2Ylt9LJiJLGU5pnyLVod27IIKsGIFeYzk9YnlE
XBfqEmJYNLeVTPpZkylEZlaqfr/nFrKBwPaAMFSbGYQ2ByUG4NmkI4OqNyuwCgapcAFRCnbopmMy
tQ/0mCgA5FW6yHic8/zJHvDgQeR2Wa5L25hkwmOZCnhXyhpm24EH6ebzeyXKWkbqtn7CujR5chvs
Yjl8e7OptvZ84+/7T0wk9XOWvbguerr4w8eaoL2f9Y8ungEBuX2m0Rl7zDo6u06WndSkzn07IMdu
2RdjmYV572FHbhOE6HEwj7DFSY9MmQ0JF727BwIWjwASHpl2MXl5eU5XdAEg1M7J/XZr/oyN1snd
TY+n4XDnpxq8TphEJ3P5ChXPxd8F1SKQ7qm78URERcJLDxupaDOYYONQWzX/RWkmLjGMbNzvlDcl
NbVpU663EBw74e6q6zAmghKBkSZVlF9V+eIHgDQA7Big/QoUK+Ly8RaQ8TTo28svaJuRd/Lz+tpV
wjMNEhdJbrZvp38nI38QOrHsCNjcbT9OQ8FqS0m5aDiMzUBr1q5oSUbFQtUygWu1lnV05YJY9H0b
k8cJJQeuMAKO6RPsY/NnX0lwZaVKDOM3OdGO7yNFAxt3ceaHI6p6G3ptalGO4mlhKmR6V8L17Ed1
jrXOheMZ0G5PISgglNtdyvL4lns2EwhY4oAdlM9xyRWsoS77eeOYrDZZVgErXeR/AtAv4WrOUETo
zJ3WvSzzzRWV9hsrfPZ8AsXYrkpkSZoE0MtemqwQJ/Q1LRmghxGfFOVnmpT0eUSetfR+TqHHuPqN
24XaleUlZuBd+cRton22YLLI66z4tvhHq8r5jhzzelDBwGoxVHb7WbP4XRE4J0vSIQbA+ghDygh8
cxBo82mAhZD/jwZ0xKQVLLZO3AgQ4kuQzNkqnDxmaJDlTx3i4ojTMycjwTEpxbOuRXdR79Y8iOAm
RX0LRMnrQrK7lJq+c7xyW1ICpq/16yFwtFqErHKiBEkaah1xvs9OD+iqOYiugMN5WGnsJ0Smg6LG
EEnPkRHvqHv3dS93eLfbS8BXWAAZWsVGyAw6VcGXJYj1N5KzA9RNcgQCZjdDv58jwmOKmsNv9zGh
5CwUq/jCO4xfP3JrObTXhj/Om7IyLq+RErcqeHl2eZaFc+ewGQ7iVCeX9/VeV2QQ9a6zeUvFcwBl
wG9UJeY54Ss+C87NBE0XKDzz3StuS5sgL1e/8FnpACqvqAmDHmHkkP4QdYdnySSbwJ5ZiYCbZijI
nNy3aYDNm+Ym23JOmKagpCxclklllcva2v1jR3sgiQCgBCKOuBKidxUIdatmJkKB9r0X+MNZiiqo
d5adWLh3Fkz7NAJnywoG8UQzpKTmx2YtGUxbfWzOtjXD+ABWsX0mMsV30OC6RL9dbQTlZNY1OJ52
lee5abuJ6ZrV1PgUfdtzIeD9+R4z5vYi1IneHla5HY9UU5DaqdJS33k8RBq4HMjysEENKUY5MMr0
wzpnJ4LNkRxEemmtWvvIyaG3qCgU+U+0KfmyBPEa92+x+fe90nz4JbQFMLL05xrX3JwpaW6qbJ64
4ZM9bw9oHYTUymJ1QojHpzaTlLBJCDntv/+yHGET9ilM8kaWZnwivnqH+j35b1lFwcJf4s5jaBRD
IQvt1Jy5Zk9SMA0doPB4Ruc9etwYDi27LLCdeMXcPpKbk4SDxuYibj1UPrX/YPuEuNN8XjYSU/Zv
n4FTjJWZBM8o36uf5o3OOqSiRxaWkK5ANenOS2XtFOk0l9iKED0Qt3VGavbdwCvjAYwGUuCiPXwH
U1skKS5jX/N4KydhQ8HXr0sNR/pcGXnnv5hjh22PTyKWqrJBVYyUcIcC8FCq3meIQI9iqo+b3HcL
6WSJsAzKYMJjhwvj884g4RNA8OcNounPU/fnVYzVgg2qfo+eEp/gbSa0NVGVhliXvYcWcf48vSiD
9t/TjGSIMWtzv/0XK6OLx+/AUqL9GnLS9JBP8MImqvNdrxTsASSuojP+eAR0AW83OqBfXjgTKb0n
9ILKjfOdPgBy5FDBTZCBEzBO9eeFFlDYoS2I06sLSFO7cG+kZTaJ6Y7vRZCGeCKMm2MXGQC5HEs2
W7QiTMKl8Ic8Hcf1q3pnIF2GYZwPt7QcK/2JJc+EUTcSCDtdo7BVwFGnSEXYhZ9ODxfj0vQ2Ips5
4IO0wPr28cYFMtPWHZQk/hSSw5LTDYmR5/BBaXVksY68qWj3HZcGFettnZMMPNmFycxdFXLBIcWI
VvVHwQJ+vQkG4FhdLDucIchzwenJONiMSLZQoABu0Gs5yYuVnkZhrVVG+zVAhAFQ6TfDYZ9PmJV1
Qz4HBXZZBL/0YGGYjK/sswlt2o7GVTS2IkTIC2JTy/pWze9cdlcSFrITfqXkP3ETzzYcj7rioTh5
3ov0WhUL2ILyLEzGm5IsTxTv7oLwrgYTewKvk3l/251ViBr2H1NsxyQSMP2yywzGrlFEf4NAStuK
EYypshniTL5uVZS6tSLz+Ng7B8iuPw+uFrWYnW1fcMLAMoH9rjmVnD1NQBNlFNdqCfY8aJlYp0sT
s+iFziS1okTNgPEVQh+P+hqtGzmuYMBxkXdQU1wAcHagGx98gPmnluDUKARrKVVYgxkqXi91QR8S
ZVKBtklhMVFzYXMt5AQS2tPKLz7UDYSeyPBVE4zgcOsy5CGjprRPjQYURqi1Rzp+NdgOR7xgWefU
LoN6kDoWxq/YMwLtcwpDZWpiRrdmnm8zSd00Sjz53NKiZo2r5ayhSw28tcKtg44czr3+6IvFhlxZ
PqN4B4wFfCFExd7HNjmtn6KPdgj+RzOPivBf7gGBLPhVo4zidkDrDjNuTx2/tDOCd3r9cUVDk6CB
cVgdVa/J/FNY7frRavh5oD5zjKiSX19xzqQvduhSbW6/bqyogw069aqAsiWqAdpsvI/bj/kBd6La
0TwSty0bwt0ruZYWCMJHZujOJjftpNLnatIsec6CK7aC9PjJHhNbxRIAHEzOJZFnbuj9KlgN3i6X
4U8iym3q1pkQwp3YRxND2m+TrpdxfYpg9Zss5cvyLLTDi8jhODo6ieohDMs+QY1vlasGzEz/5m37
z3SzrMOXGVgLJMTY89B2uW1RhfZKYWOIdXGiuxS1bHOBLIBxh0Z3LOLNF/bxMNA96Mm2T/Knpz4V
+bDN+3whEAt8Zf2QBQimBNvLjVzkX8wPgnS9yrgQn4Pe4o68Pislo4IcMhS9/Fuh+A8xjHpO8SxD
ytmMRNeVH4qA5RAIa9BsPdnIjwnqylCftNlQsdQX33yFrx1a4iZgVJ7Hi3PK7+zyOlg+/26RYF5k
qOt5Frvni/OCEgthQP+whaxDj1TZ2REQbMT6Shr7gFZ09KYXq5Yri7zNkL7VOhkMr6jxRajqpSz+
BdTmEndDfHttPX44edauBI6Nb1blz7z3Rd77d/8FE8by3Elkt2yFWauVqrhrLTHP8G0PZh6+fIUb
VeMldayfLoW9XrsVKPI0FtgR25yp6VwjFM0CnhEsoOL6jQr73HuNjgEU0Eeg9XEymcbAWRfJDhKf
NgnfZnMMEqH8ITX/p1MAm95u12qK++6qScqtFok6H6H5Wz0h1mfq3XvobTH+EnZSP5YY26HWEzlP
Sw8/ENkR+m91V99pG2aGedSJvy3LxTqDPJJXWbHwNUw7cAIwu/X6Z2vPKeivFLU9gyXSJqRWqOxc
tRQDBkerF+bHqzZlEmCjwgwTFctDTtZ22PmbQtktI7Q3fsuLvjUsNQTDMiNv/juiUT7ymT5BPBny
4ixy2rroONdFouHoVYLXdXecEhlkbhoImPwLA8X55+/bamxoL8g/rWai55FJDirVaV6eUqTFjFAM
eKLuG+i3qkjN/Lb3Ox4FHGrawGhmE5ig1s2+wAT1LzFCYmtBIkwwXPdzY5qIEWuO6V5wKvNW4dc9
U8wX8UxCcPhqW5m+5UM2B6piHWiculymjr7WSfIt0BTOKFnG9T8NPhpoJxAzxvU36qHq5kYElE7t
xxzEGctbgYZzejtwHwoxszBTe4cQ1WS+WoEMqyPAnT2iykUkNQBYZLWSzULN4vE4muUp+qmrL07m
OoBbleRPfQNsZ+3PNiNdklsHXddnad5eixoxaIqYSKslYi9EPwuV+/H+UIIqQ+PIbyUDt8Ws/CV/
Zu6FG/PALiVDa/wBtGBzrfkythniWzxCg446wHmHqheXj33u+0Lh9meOUwk4bwM6iu2Q3gZZDFhG
gcvjABXbOX7I6MVGfJ4Vows2Lti3qHITQMvuJZyc1AtS3BiZnrsOlJrseLA6CZjZqOviSCKkCTyH
2a+jmW6jM5kIKamZ40cOkfVtDVb47nMMwZVVvjSlH4pnn+Uu2EhqoB9MHevQNF59U0u5zTGK5up+
sQrAgkZ44dF4IVqhdf0w2kIMl+9Yfi0ttyZODLOPNRRwI/zv+zZzHkglzELCmV/vc8kDs0a4N99N
XZpP1IFTImhd7R5EMEjf7roEMBfCukK2ZIg1vV77LGGTWYvacCQT/gqzKo6TrXyAiovWwM5TW/yM
6pFm1X5ky7Fbqi+55zLX2arLx8aEg26y+rmX6bK6GVtj6i9kkODPZ4j0X7KncjngdM7cvsyVXAex
5ftmyGpLFhBZ7zPAxqmsP3aquz6L8u9JTo09FMvBz7u+pSKTq+qSsb5f+XRVnJf3LXrcYhP9A7AB
ji9IHQdJ6OBwSx+LtdTlyJxr2aK7N+YRcixHLF+gHyNHTmaRT5f5NBK06da0brdz7PM7EcP/Y4ax
n8U1hmMXr4vZ2NcOX5MZlHU0OmTpM92cJlade1snqB40NLxK9aVUZugUloUsRZXTgTba2SZdYSXc
g3HILCYcT/I2mGxS7OYjFwhhMYmNDM/bAZ0pOZFQojdYtfbYbSeegFvQuVbLQAhJvfFdoqYnzFz1
5xt0edZerhZ2MLnEAMRM/UcvJX4En6OH7hpPGm29nhhE5ohyAgZSXSHOJA1+rxxcUnfgnoe6g8uo
CUBAeTHT8+AWgDzVuM4OdoNuo1VIePukvVetXXwiSwSvNeLa4Fyxv8MVIoN3wW5Y891QdxbLVIUz
q67S1KFp7lwr72ZhteaPq8RiQHyslQyEQdRT/aK8Ygzhe6x2Fei88LkmVPEoYpbHfqsSblCqi/pS
u70ZYlDBcLrnlw555HuobDtCafTEa/0PpX/rpPm8Sxl+9kSEKQOh+FMmfqmm4POrqfOWVMTf2Sni
lzj9sVVlDCOXFuAHYdGxvXIRs5b+NYd1ieZpv9vUFO4N65ROuTDnKEQCuovmALOBOtuD/z5jScPn
9X4K0OzI6I3RTS5eAD74c6II1SVytUht9Zywn1GNtABYaM6KFdaAAezRO++0CgC+c0hBXIrJpNNQ
I5iXB2y/VDj1irzv+xNL+vUxaB4YnZU8W2xcmbDw45y4H3C+aNCeS1lVXggBjUrI2qaU/Na3JW6H
w+uWltxIRVjCL1NGRWPAwtpTE5m6Lm0KuphE1crJjXWhyZgLjXctwXatdhrJ/Z439wuZ9TBU/eIe
H5o3EES2rUqDVv0x0VuNZU9KURtDZDY92jQqVPlZMRUAC20FpzE0aCntt+4slLs9AyzDyGiGjxIZ
fnwO9q0sAUEFYPQ6W9FKS1SAn1IJmEb2pZ9RTl33/5p88b2+EPIcOLRGOly7kZJE7lyG46ndLbL2
hixNdu0tekD1Plr0ERrDiArVhf23TwjsyMcZLKULUsBXHzdSAdatPhppTf/EGoZ/lPjNY8Wj/Zrj
c/K90y0kFb+WH2mnV51YGu7XiGpGaunMXB+b8AbWzESZ+pbLZZQo4Hp4FwoG78SUGoFSPclpEOG+
g3hQ1o/v+5stAS2plIpyX2o7lshM+c59cFjDo9NbYoBgwBDz4y0ldahgsor9pjkprGEICbjJ5AuT
IrVj/0cUaANIUsfJJEodoKsBw24GYdkWccDi4G3LL/pvpIZ/5QFn7sBrWGld6pXJFq0n4eK9MHj+
Qemhm609rvoJXpOhvvwi5vX5Lu9KZtewzXvXD8GT5jliCLeEowq0GFc9NdM9Pxy4L+sYQ9yIlg5p
Fyu+zI2AsJSWAxnTpMsq6kWupRWi7ESzSF99XIiuNUUD5+w4b/Qh+Ekxa/5lFunHNydcK8p7uouF
k6Jue15+UW/2KWKtktRYTFFUab6HQQfBpqDX0y6+Wx9wk8NBFbyVGgvczl1YN4qkGnTkPr/wv/AL
E6NkAxoqt5XKHzqTcjqTkKlXhCVzGVz4XrFlsMGJOcIMgtBIKEEo7bXENwUi8hrAwj7lSIWQ9uVH
NfaJi9HTNr+i1lul1mgZ7q55joEdsIzS4eonfFCGVsubgQMj8uK18XEUG8Rd35z3W+nyd0u/dUnI
tslB8DfNuQWY8ZWNU18kZcvVja8gcrg3q1jWeZCXeS6XsZf5a5SaYT3JhVw7dg+lVprYTbWYt7ff
CA97Ku7C38t7SaEjtMHMyXtG6xhrPPygQYBDp/ypsYhmv0jYJGDADQqKWpCsozgKkU16Dk9ycg0q
y2j+do75Gt5GuI6tDYywDliIG8oq7koZVCR+D4QjqdHq+hjiyis2Op+56JQqT9ezL+9FRoR1m8ra
FcV58376kGzasPX6M3aofwixYOVjhXVdrJxy9/HtozjcAPiCx9O8bDjd8jQrW9cUBXjYTvgtRft+
zVxCYGjxlL8vUR0g+EKZbSJn6yrs7sr34RzJxxvR5y+zDZNym48TMU67m27dY90vC9+sZJCa3naf
dDj8aPx9sJMTazQjf4vKyU2uvSOBOB2xqGKGglDdM5TzVC96VKNWOFbIrghpGwlb1mFuuHQXRro+
fLcu1TXtXfyI2Cuj71wJaoOVQN5asUrk5pLoaUkeGRCTsz86A3edAqaYY0StXr+wWB6gIOwgSfeR
7dA0RTJUMglfT1OTXGUQxi/k6x2IEEF/EPP+DxAhtGkoYPjOP+aTkeJ0SnJe1oDNxbQ3bOohE/9i
SM2bjf9O567VpfOue3yPAHUnYOkMD6zgd4a+yAkbIgWqy45bhA7F21b4VZPUIfT2bW0ZlOmzB/x/
x63RW0aD6Ub9zFh2/AFFpQS61rqh7FExGSQU7Zo54MXTmouTh/klTslAVTXBu9hx8erCDvj93tmG
DhOqFx4ZS5fINdh1SwY1dunnKyBZoEaQxbbf8DWajyWOvlxb1ymHVAhxDa46dt2EdLHPeJN4uoWu
MkDa68cliM6REdYstDv4HWWrOfBU+hCQz0ZFTt7RZmOMkwFrZOWzOwNnWW84z0V6VK8HaxUVnWTQ
bMeMRqctOZct3DEXSXJ0hJfPPryYsjhGxXsPtRfOYbvBgJaw/ecgSMmGd2I1HfZAGOfrKzQeSOca
OgHeoNqc+xgoe420va1RhFmyv3P9arvRNIpr1lBFz0sy5hfORBsmrZ4tjEyysxr2jFuGlec0VyEs
LQvcR0Qf6EMKDMT1lityAROMJO4xn+2OkVBbqfL+uDnfOI+A8t34L6yix41TQZoCdBVCalK2R+az
JBl7J6JS2NnFoBICGTGGH9bRhmULdwjbii+5hO1GxIWi0gK9ZK8LjMx1gxSwkb9pZAoUBvrWcFKo
X4Bb+TZHhxSxRjW6SfZgfZchru4uuXWLOq/qsBfTzaT9solOmrJbtWHGGW4c0W1embRQQjMC1TNW
K1ijG1m5tsFLtu+FX3HFhUFq5axmqeHtLg02nC2XT2yria/YOtLyC4mrlhInPoQ1e43aelZGiNNF
3+nyY9BKMaMWqGyHxUkZvpQQSaFuiv6xklfc+R5zqQ2iDIIAC7WwtDMploJILyB+C6sVoqbcm1MI
WER33HZbp5MqYgOWfMQfhy2ymF6NWlGw4Y9CU64SWKxjnMBAK4xP0bMOEHKXq5/96y+PuT9wHIZC
Mmt7fUO5W0Bm89Pn6cpqdj7G5OaApUs4S2W+YXs6VR5OK6Vrb7r1P081RhTGG4pjx7CP3RlDibTA
TnP/cVA6Ec96qzCcsRhYMsePO4jlb4XdGzGd0zQ/Pnic7s5q19K/T0l8ahjmize9BH7Km+FKaD4M
6ePe9n7IEDXTXIALr3WYYWUVwpG/UfbvTpnfZIUn/0PO0iCOX3O4xxkNcInAgQVHmnjJSKXv/OM+
5q/wE2/htFoToKOOPt2wqMcABoUWsl0oUd3hq1TNNu9kAFmRc68UdOjoRX0cu0OYqFwMhIAea8R/
EvxAkLNJnOs6gKQ36fDwCvULGxZIZg8eKfDPqJDz/Rkhvf104w98mmGN4Ynz619enGJVHPptFkv5
+WE22l7NL+eXWlS+bzdGFSaj/7e7pwf2AC7wUVfHy77VyRHok7skLs8AY63mQtfAVozvbPVB/lk5
qXXgTrndKvJja7SdO/Z3UtOzBTuTNNi3Zc/s0UzSkQYHrQOULGIO4Kkddt8smd5baiJfIx2TFuge
nZ8ejYBQfVAeb1HhvTxsPFpOHyXDZOpH/qImlBmA8Atyp/F5zTX8sWy5VoDWFklexCMGEfIwMJZX
fNhgq2CakKYm/Dol2zpKjFlCfFF6EIGFU8CRt87TK6tCBOTbHfYIHofho2KkCv7cjUM0xAxd5Ekj
o/dkWMmhddyXQWl5Y1l/xxDLdYXmU1NrIUygOy3jupKuwSnQb0U4HkxMqLXWHJhIGPElyy8Z1N0k
755/gZ4+ZREF+FA7oitYpXsz9K797p/TrzZ7Xbgqqj63KTKZVtIgsSoTeMQoAarWcoFsLSAWXliS
dL16JWbxlOO9ZAa39oCHCtE3egbl1E6MkIZdoy0+J7V7jVPSMqKM3y0aqZY/ZIpxkLHIEIUEAue3
iJXT7WzVGlERAvDCJCdMBseOjJARZTCBAiTC3wP2ZUIU1QD2AdY3zPlLMgR3/jX0U3z8C6HRw0jY
Izoh3uMzgm1DIjhtiN98TfMnQEGKkUd6Y3Dx4d+Ewgo6rT8USH5JEFAxNFJIRdxiT/+K7K0YG1/i
OTyXXHvdfCNaeBG9Tex0kLs+IP/v1hSlaORoU2PVb42hpEVN2bBAQwpDPvLNBLSm0EmTqBegpaHO
rWXwk+wWPdgduA3V18VFcFSFQTo8bB8L2VAnNuQIwZyoFX1eC0fRkuEpmBtzicXCPe5+NX3Lb3Cs
nJl307u4dOzRTin8UWATO1CAznvnim/5Fii1AogqblQ2x3rAq0/B+R2bum5H4uHXUJihHHjG0Tt9
uiKDJf+2Dd1jvcmmYdH6Ff2qmwfNbCD9FSHJjNL8RSuca98y1ZV7Koht198f5yWskSRzCcAIiBAq
3HGvc1pxU/vxTqxd9RWQrDkO21Lfz0B39stxk0H9t3hSrQm98IDrsMMK46AAUsndgxWNlkmvF3BS
6/Epysvs8yHe/RkjX9NNqV9yAYeXM/hSdEtdP1ZK9kT1O2a0g/3A9qL9AUiy5b/Y5JwjYfxGJg9v
2EUuspPHMLxhEu+ZVT6+qG1jl52RvBtMCoFvMtrCg8lcBcewR7MHwS0J28MpClahnd4gFrunpixb
AQFrZknlIfDaYdU7KmghyQGUhlwGIkxeBCRSqU9yQMrWWx4CWsrLCni9zgxnFOutWpqr8gnZkNxV
4tViXFz0xwjGZBBXuUryrM1papVysfKns6N2o9reH55QHQWGyFVSwvzsQBJVUiiEYU8io+eQ3Gxo
iqMWAgpMWILO8NjX8V7D5PH+b9LCt1IrXdLZBX6TGgAS75BlyCwzSqaz3qZ8/RhiqKNZuUZFzQTw
eO3valYgmulR4Pu/+5LFCI2WMVXK5Hr6yiS2Z4RChw6k+pq4Yj/ejSXkdQyWtsU7V6BB3TnT4Uju
9NAdM9MVxn1iW0f0a1jAyl5tU5k5cgl+QGjP1GyxchEAo5/AW/XFd6dO/KQDtb6USGvkmi6qkWEm
gFU4dZmxeOZoPIRv367fMBggzGiOjAHaA671+999ZYDYQUuoZ8sqkI2zSqzboSQqgyv2qJctw2lS
Xrl11OUo1uHJ0RiendCCjHe0mdLC6gGbbJ+OGPFxz1A00MfuQeeLERrzyEHnVnBemKZPsOR/mOAH
8HNK0npaA+Ii7uq777OtjKviNAKbs1mTCNEEhAxLbaDckzYlFY6U72NwwPS9QkeNUiMeAJ09MKoR
zvaYrt/3k4FlkqW/+3th0akQRBr6sgmo6PG3FOXJxlbsQGkg/8EmVccOYG57fAiUrr4HdCGrha9Q
r/YTxnBGNaev4wlG95lY9p9BZk/B84LufOM7D/WZ/lUh77O1cAGA2OWGaHy6RPZevWENaALAATBb
TPwbqTqUuruNSfhRKe2AbRBWNOgJk3uspykyEo23LQt969GU/h8hGBQfKpzup+Q1P1t5Kp3VFXuG
TW1fTCrKBaYSOnpL0F0PIFydbst0XL8UK7MssObmCL+ubQ8Q/t/L+UYS5a3FLoY/htyDDpNFZPuU
jLdZO1syV2xvQlokFT6ttl6lJm8wcDwXyB5CpGBGjBHh9YduN9xvkggYTV0pZnpr7B297ZBDUcn9
iC5XBQPG7qU2geMxAoSihx4dSCl+Tx8QaaadX2VFjp6NYzKwUHXMZlbHSAHVCkQzLVFForpIbLrT
MzHqdx4DVsBN17pZ7F811RpQpaP2gaVSuuwpEWFsEmNEw1SLohAHOwaOrS82GgMT6Ah8ubaSzqrS
4ZvWFR5WfjbasVVPCTUyuOOSudzmA4uophGY/ufQV3AB8p2o9BrNaY2440zqGA8n9KNnkWC03eFR
3GDDb+yYL3mOeaskPRT0BkatRYxQXNzxqG70ptWaW68Fmoa/5KZoq9V5iPLp15q57jG/jLFlVGWg
oWj4Wg/9Z1mybm0YjGK2+xWqZzFBEmyTZXZp8T3eJQQ8P3q90QVK+mkHvP8l4pCKzPEJd+do16Yr
hjVRYYwsdG8Kvjqhk07oLyOemWmTTSnQJIcST+nCTixBbHE+rKo+hDrtGElE4sVApaayqAromduz
iVQWt/GxAHSvV0nbAD8xOAbT14BiaIFkT1I3kxZA/Ynmv/wZsw+XF9JN9Q+3meTyHPRO1XRoIAfB
frGBOCe/CLkHq5ISiyE1nH1cw6glNX38IEozEfMKPoSZJp28zgT902Rkq1RxKHC4fA9fpaUt4f5o
4MfYFQPRjgdBoqTfKGqzL8RgzR//mVomjQxz/PMBugH8pnG8h97GmWxBhYnRDLeaYXYwFP6w2swk
1cYYGielBeYcDNb/0Us2mx5/FSdtCUhyK3DBtGR2jh0GZ0WxoiKzb6KGkcykn/SiuIiIzxL1X6fg
ilB/Uiianz5CAml2TsNN29sdDZuOQypUhABvlk5xuFHFuzmSr5mTT9GTIxdY7RoW4uHDMvUdN6b5
yOKMQXTmEkzVbeMVj9t44wANIAAHnM94UJwv3k6RWeN4KBzX3kvC4AaSvXghKrXuoczIur95MmIc
iobxEWE3GG4dgAtBjSmpW9krkwdcwAYIkQh4E0oLP244IrkK5W7ri/yTFOzdWweLh+jXHrqhfYGG
aK+oUsuYS5EKwW6ykOSV1iKPpORuKleiSS3B3AuhsEnsmDfaAw0oqjslxUI9bcJTsd1n7/d9oOPs
jiuu2ZO90MPliN4CAORPJ1LctBCJ8fHPthSsNNH3H9DcnqJ0tpqGzFhZ0nVlEO6A1+laGdTsKYeE
MLu/hXiTxjJoHETlctDNrCjZzNNj/B23PHpZzTLNJCVA3WYb+D1RF257o5U9qQO7lyKC/8zBZD1E
PGgKd417DxYARJFl1kJ9oy4EfVCSP8/PIFTvqTPJQAzziarcygG1gfaO7/4w5tiNfm/IgFEB6TPF
D4c55WIgteVBOHKilJTtZeb47R2jllMMLMCFdnVIB6LeFlr70Gl/JUdqvY7kx8NKd0m8iGVomUh9
/riELTQqx4da9PeXcDz6ew7VrL5Xa0GV/gzGiClLhpE1zBUl4sz+2enYZVzoQciC+YNzg41rbRy4
FdS9QMikuCj+Ckhnp3RnGADPhlSeJb1QO8QGd/atDVss/A3c+e2zmplHutPM1yPnChuVeG2CfUzM
SMK8ixfCvhnSUYVbcs+ymiD7titR/wWjU+VS4eUCXnFSlavD6epIHC2wmf2OU0yjkIKkWvZ9xtFy
GvMucDw8QiExUeQ7y7eVYt3lJ6e0wqzGMi3M3UiRoidwCLDWRHMWFqOO3Z48UkTwFAg36b/M7iOC
jCkLoVVOoEv7/5Ie5XOKvAmXJBV63TKNHM4W1YoDu5zYAlRPnNkxZxRR5paWHUT3DpGRTBc33oB6
xnInSiTM387ZkE1whc71nInW+pzUIN5XIOROZBZ+T/vIzBr/fQ9HOjh+7qmzgf7ELft5J2JJ+Yjp
iLsUo5lY5j/XNTg2YsaYrVh4YHj5CS5ao0lBuqD3u0a2WpM1cdsSJ4GzmT9i1bXRmZfj4aqHySBM
A7FIIPOTUIcoIIgxPA8hdIpmXpOM2Rnvo02EJZ9mGI8opMxm3ZQZe9A46qsB+ZT/bFpM1+Fqei0b
+F4hSSurMuqm75rH6CnWrNRlcYYBJ8eT5B7ARgqEXexX7gxYHfcvQACwJlIwcsIedjrtX29zNqiG
Ru8rCjjCshEk7Z6ICwDJEfgTqkQdPHiBcJzdtVUY9URJXDEmlILutpg7Qq7YjLR6gUZ2uj8VljAq
GeKuxNPQEzmP73eJ1yXZqfi5dLALatp4OW/4zc4IZq6k+7KjXLD+zVpbamVEO+49NtducBvITaOB
UawNIrGIQvmONeu0f+L6npuzgxxQ3u2Mzu7/q6Uxn/+DGz5fyEI+po5NZRq0jVE4Q09yqLul7WlR
AR6B2isQLhpg7Yqjcw7jEU+0BGA+oz68rrjEMqIdQ5r12o9AdN1lZyf8pjy7NG7s0OG1blBN54YW
7mCEXl4q7FgqSfjOcOp2aTVj1SanyfXbOpJ80x9Tb4/t5uL0Ab1PCT0T+kFp2W6nb8DrEAx+bntS
SEEN9T1tI2IIXxqX8I6uRoEhwpmSnqAALX0TorGyVegCIXctcNp7duq+8MDzXKsVpHEuRHcwlIpu
RT7pbyikPnY63RxZoqbgJXzuZEAZ4zUO8kjuv2qnUfSY54762ksQCWlJDG+xexDjbR0KdwLatW/Q
mZ6c7mRdR18M1k9DGFTN6yqKYo1QzNuXmcuMh6qnwPPC6rADBjRqKv5+yjRgjAYLLjZk8BMCmGB9
o++F1YJTk6vXAcv3Pu2yiox9lU8MWRUaNjrTmzaSsbnsyezJ9BS1iFMBcgTiJq6Vg/CExWLu+9ld
ILYKMrrsAlOYm7snQsa6Tb/bP/2ouAUwaYYFuB/Ua0jUIp7y2xHeVRAoSyCtjt82j07O3/su70uN
itrkGdYh0HwcUcLXoLDk7KnWRTcK8nUbC3QHoYZAxunr9RU2OkzR8stmlijqyX6Lk0GjL5fqi7DV
gLvgTj8vOwlj55cmOtVhnl0VgB5RIRppKG6EkhtmPEfSOfvsjuKLMAivJlENSf8u6gzKQO2UILhc
Mjv4+tawYSp4vdtoulKErEVq+/8dguIVLMldHHAiUe7/0yP4OGd6tOhRqspE4v0VqH//H68qxqNW
XuhOGejfOlL6kmjKzDyJKrphXDVaJ3wF9VVUvw7LcipgeSXY/ZCPCp+Q5TQvyGeMSuIdCMwAPgjV
QVnqNfBjHr7hHtjIJy7muuGyBIy++82la3nyqvC/V5LtL3kzsQtD6FsSsMu8yXqWqDio+YYoQ2YX
x26eWJwG2dffRaMw2/fYxLtmChF8tbVlw7WHre/BPwLAIuvKyQ11ZGB7p2kWHLcBFkhF61URVz60
dFBSJmjHyD6KZ/Ll03P0UFLvvR/UNqp/IjFb0JQGNhfCjyaHSvwpnOMxvc+GKHCSELrj01YQXzU0
SJjqqACi3H96SKgxVapeaEsKhkB8u6HKrV0rQA5GcjFsWGf5wvT4oUVHq2j4ggOG5qSLDE44Idkd
rNxhne+oRnLhCRTN10azVHAujAhj3NYLYqXIpaC/J0Yh1RY2qLMWb7OmOh7+SacUtRk7OmFFA/H3
dnOydoInYd9YocImXctIO6/RGB0y9i0bHYCXGQG/DT6Sl4kCp1ZmXr2kFk2XGEHlYeQYmFnCeSPy
RAU2XMK7tz9tyGAa4NDd/r1us1CXl7V9YMs/YQSH51uZqGgGTzN5kgHMIdzJ8927enPkTLFjg9Ga
utaqFC0HYPa75UcDl6iyqe96iAAuiynEshWy1xnmlRoonR7SPJc0xLbb3Y/pXXY4aNxTkq7aXny1
Dlw/8ZL34FqH5Pbi/IGkKzs3iygHkTWxGz9BpbA2vWpgMgbe60L5qJNlqM66rQU+68K3EUfzwgkP
ntf9SaVVvGaPkMkDzHLfSMCXjBmSb9lQj4QO5AERfnvPellaX7Vzl8RPVrySWyyLrWmgBr6psDEb
xK5Q3eOTKa9ousP7Cz+SLjmIfDHFLudd3hyMfVSTe9+rtE/QbpEQ9mXRYbopeyOV9K3cvXhHiFzh
OsBROdehQuuYtjv6gZyd/LJ5Zfl6PXe7zmWmQXx/gKHzclG9QO8sm4vVlwW+SunMUavYSe2uZFjg
u6ptn3ojUtodHNxtNfX4yEbW2nxsvpDZE2098vnVEacar/O5T8f4TB9xqOVGrpYP6CvXJctWOSOw
yfEdjcFywoZmvB7G1XaLoiujK0tVV9EQ7N4DCIDdEFPtzOo25368Gstuxm2RskOWDeboOF75doVE
6kWKar6Ey2ZNZsiDm06d5phmnypWNLFpdk4T3VQI5+9Nk8j6gJSJxSS3DVKNJiskYV/Gjp1twvGK
Zu/cJn9FbvZvqGmsC1TmS1XfSF30XXsjBtczwjRSQYfkobXOkNh2kQuGgkOxBksgeOwYqjebmwfE
8l3cKgSKI8Iu1vdv6+jlkYBh/XDTtXUVKrr5V9fnwGa0x+mrgHYHQmohoUD1sRFctf5BvDNhLCYo
e95qHLpQ0ZBq2N0pGQieeBsqfbO+C7L4fuMkXRjhhPShgpnzveSCqSP+dFgs2CELTnrapGxCsz8i
UVoP0BmoWob4d+1DhQYSiLoJRTotyolJNqgBsPWnY/V9qiUWKJySdMTBGQ/7jTd/fhRuCitsCCL+
3xAVsACAYVYf4QcyoQCQQ0Vf3EM0YU/ZdJd1AVobnib3cT0lcEr51+hcShSBja2XlXnfD6DPAqwz
3aBMzq4vASw7TFxzIGiFAPFIXLDvCfW1mFY56Tak3jn5HV49/smbYvF1LLzcqsoEuLpv1HHZmhEr
h8WJ/ALV6Cku9Vkrwa1EGvOfIpcRnx94vf2GjXcsL2TDenYM+/GxMP8g0x3aFiQj8aZvGT2456sA
49pPK3IPEuut7xP5gCWn6pQ8mxFDuPneMzCRQa1BROtJhHSCn3TvdInUuxpyuZ/TgshWoZj/yCv8
lFt+8ZwfD0jO8er2BR5NrX8CEAxN9aYc4NB97DkzJswtyo/mSmilUVYDS7ZdD1HUebGotHKC2trm
1LZL//oppwgp5pTdRFZVGznWnd6ykcBu+eqKQOQ9CgPb/3YMUhBhvqZ52mQAbs0mTkn/1QsFA3BR
aIgdy7/r2iVDOmadiYudJ77eR1JahRbDkjTLlUhA78TZnjiKM43CRgH0zzZjEsfQPmKfYNdhvw0V
76gP6glFM/kjZtVRxxyqHFUuJYMtoiEERGgzXKWypaFXJdxOhEnznSwhT8+Q22rltGAZ/Pj4oWaz
7jIMKVMA0CyddrztlopN/NgxiC+yBSIkPrUfZ+bAZJXdxsEBKUqAWiIaa8zfGE8lD+lIDhD1QBg4
YcwezTPmwiRQm1usT5gpCHe9hQziG3lbHax+npivBuGxIJLIrjdyB+/WewZ+V/BIJhbXjfU+rkaX
09EkaY0avsmJ26xpzOcZoBfdH4z7GEsYuSu2tuIktDPqtldxBp942yxbrLoYwF4OHWgmabkaoH+/
+mhsbqPGAWhRlXJpMwhRtErsp9gGdmK7+5vLMnuNftbXVEIEdL08cKDOmGAcTtHab7WMi9Oypuyk
mHD2LqXKQQRzyb79uG8TZzjses08EMzwmDYJUlGB/aFAZ1rMcRjJqMkuXNj4vu3yizIi5HnOH9HM
JcNGAUlizeWXslRIRRcKVyH809JpTpxS4pnakXmbtdbKZK3PCMxmRqrRNTuXr75RfE4idsQYb3Iy
+nLbLEvgHHJBb5mjHvgZJVguDQgslDXU8QakyboCoGG57AP/3BdKtvVSKiL1IzUMqfCB91Ur9Kf7
pVChE2Q4d0tdAaCAYlB88BbiVCwOt3qZwdm4lEuqgNgVJ1horKBKAYTHEmyQ9H6se0VJR4VZxPQ9
YKrzlLIVchMfmAhhUrqChRudbG8ufCOBsV/siZVkkFnpr/lvj22qnZFEJLfjDnWVBCxk4DRjpdiP
wR1GD0C/Tw+E6C2JIOO6nlKQl7opvEPV5bgYpfDPYK1iL634Saiebq0S+x83BVC2xxqaLwKvSKFY
JSaeuj2BUoSN0MCKgkFABr4a/DqFLRTE03N+ODuvezTtu30TrskQ3gK9LO79TO45uHsPb4IERadb
EWUOl7PB7pQweUQrnUzYNGj3PcLtwmBVASrUERCZx+LtAz3ZgwMY7h6V4htuh1km1xZM4DcL4gc3
upplmLq2GQLR2s0AblIFxoAyFNUS7l5SSeuKm3RJqgopltJhLu2kUxD0dFJ0uVTmdRk+TC38T5nK
MJzRx7sGx+VtFrN1Aut7XRZO1/2ycfrR7KuDYZL95qWuNh9Pyq4I9dfew102ArU+VQQCUqvlodod
JaSda4DcaCcrEEZi0Tk4WE7mm9zKxL7aAY+ZItXCvxsrf5BkNHRWrGw1xAv0uWGcwPPv2n0z6q6c
TN+nNjJ/415u+kBVzhqYhOmwF4+JBo35k6W3fwyGl/MpKxp81OQXQuNAaJ1dQ19jbWDbqQqzYSfv
xsCNqkGceii3y6x81EM5xUv/0IQsvzURvifhvJU6h+No4zY7/rWEVJvwK+IrGe+5SMA2qgTV8jM/
G736Bc+kFuS/be+/y/bowYeQ7zEBTvYy4eHZUiu2WRXW7RVlguH0drSIcOlfIknv5K4/i6F+1MhU
65JIIPVjlaVxjbuhhVS7CW7Pfo4dXYXpTfbd5xl7wbxTT4rQt1bTmcWVk0G9Rq1I9G7Rr3GE0HII
+Yxq4ev9qZ8X9YcLj8GXsPiD4a7S2tPGSg5afQz45iIZCcbz//757m0stbRtaq2DTwZm/c3xQdsV
XBeflc8DgCnMQ6e4WfR75iieIpxwcqDXoXCr4e4gzDE0+iwTip8RnrfjD6AJQmu42nJ6Kqh9/CpE
SxDJp3zbuAey2l1MxzF7XC2P5I6X4r4lNy5VmKG1xb+PAh57fQQe+Bzvp+CflEgCB575zHq7A9Fp
gh8P+PohVwXkUm64GW0dVaD/Cok57XXR3JHL235beReZjKN/mL9bkOjrmCPu0qZ62QQeEGdtXtD2
89yESTxq28bty/kMlY9xhlgB3eiIWekvmS5KhzkuZpv/vcGRPKcfddyM8M7/DAror6spCR9S51ZI
f+lnSyJW0IzLUw+mqGXfL68U48jwD+06zn9nvylWOP8oEvg4cinKQlMmcmggrS/x4N9kZthO3uVV
nplcuFjFX0EI3PbSmYGYr3YImjhCvqSrYAiQfivcmw6ObtfChviiQMoplqKu2pI7ZeeDKzGwTUV3
/p7MztYDGGl/1rxk5XrMz9lLwyIDF8x2EAPs+kPO4TmT5GHJTY68pRmEWV9vjSVRLIvij5Y7UyGi
CP8b/UHW9YeLdui2ryzKXHUgXg+/67mujlaEGw3ZTGjTs9fqk1tsyMKehcAWbc+KYZmTQRubf5ET
NO1FvLLoqSzJgJkq+TYx88Dd8EgZm5usPE6FyvuU0Vy0Xf6+JerakQ+12dpY9sdcFTLyasY1SsBF
Fh051ErwlNwLAaNF2R4b3GEKiSFiXHHsikqP5lgJ/7Q14eFvBlBI1UkS8D8o2r234oT01m/Gt1+5
u8ShBFS1nucb7b+NRcIsrCylLInY/uGALG/u8heQdN5jVwaqttqe7POaAjnxJmFygLW8NGwVXpHb
oSz4r8HcI5K5KxylugDHKl6KHr6m8o+LmcIO5KZ5rIbAHpT2AsuNphTuX9No1ApxJU7IEMH6CDzG
wJXjt/mJhnL0OuGfItjp65PSqx75G8RCI1PgrwSKCwBg/l+eA97813Yajq3vaHWjobXr/hSdYgnF
awxrmxr8HsIPXKIreMdsk67dxESe0YrG1LPaydZszlSvMBOVRqUemXQm9d8J1+jWCiYCMmWMgrXp
iPp5h6k9evExvIeeADNqd7JDdtg66Q9hKbfSa8Wo/gOGvghVOFVChEj35tEg5yr53Ne3fSHlXdq4
JIEBZqx0zqhRxQsdTuK3ExTmrCKsvvzcWhZO7+ETjG59p+OqIbLO8DjFSCKV0syAmfE2N3pAbdXd
ISa0v4RJw3Y/Hg4838hXUwr1dbeRiQUdOBf1yq3q4bb14j148MMyqL9aOisR2vwW7jQ6JveqqMrV
GMLGga/dXmHYYlS4vyd3RtRQsoTcMtQpn7DIcG+pukB95gVc1i4zwXwZbSEjOCQD0wCLEpnVWs+b
vzKyuOe9XimmqorBIjPQf+jtjj4YGxtb58al2DpQMySi99Yq+uRW66dIIwjDEDlun8shGs2HHBlz
E+JS9y+MmHh7B2SSRegpc7lKpvQTBb3LJ8EFAOLyYP4oXrlCT1XizFXoi3NclsBFZ2uLjzflCM6m
m6ZeTV2ldS+lMkM2cTxlAA+kN0kyADLqd/zhgC0Kj/4Rw/38NTcpMDecLdf3SBGLnYJxUakYWq+j
/wBlRzOkGLULj/GUQSZMwYxxLd5SBz7VXoCdX2mOCMPtHYoRZr7UWs0AgSWVAtkgjlrd4DTCg6BP
bG5Q5PYOqg5G/wS6fUO+Y9B9+2tU5TdbQhVlOx4fCFyBKWr9izW0oFBmnxnrYn/Rp46KlKZ9ZREY
YRzwbuWw27L8gKkjwy9EFQs1FlpyLHVXOefeddITRPXbkrfm+2WB+8y3HE0rPgWhg3cHo6mouHTe
OYSTN1riIax33XJUxvuZw9kSklnI7+MfH1P2DhEa+K/z66cW7SZcLRmRdGvA4kWfmnV5xuSP5Z3Q
QfZGsy6MRE2zr3rNbW1Thr3DH/e34pDYxhnJWJz25R49Yb7WPqZIeDLU1nAnLo6fhvg9vHhVQfFi
GKYBm2NUA9Xh5ImD8DKXSrSOOAGVnYX10okcgLKO2NDhUJchAJ9q0OqJhFzxNBf6XlwBKfkkK/t+
wrGaaXU6sgPnJmh1ET3SZrRycOLZ5h8nYfAp+XqMMNaT43B95C8NKojDE/2B/tucO2/GExhTleTR
OJEvWWfddp9a2GOTP8qCqUj/XodEQYsmumzXK/3hijJ9HUlo4ow8sx3JA9CAuDlfB1WrA3K28uA/
ac/yrgXYgyhXk8Eg625kPJE5ua77VL2PnEOc8zNdadfiYpp0DdD/2MtKOWAMHweTZnfZnrJ4OfUN
7EmKC0I69NMfWRG3aZogVN1VPvoASfUf4+5HKPkz8EE+9uNmV5huRh5d0oufxz3jnsw+cAoeyJ/y
oWDOX79nDPQIJiVwltU04TAM8sYaRHA0W22vVImwxj58ba8rvqAdCp9y6aL363XQyE2RgVUkwGAj
VOtPnAQdUDFs0S8wRqADY0m6CCdjg0tNbDOzkpK+F+j3j2VHG4DptVII00VUYLu87MPg5tTBP1Mi
bAwBkmoQShrxv0snTOcDiim6wGsWroa89nvLTxew6LNP4RsBZOutFdkYmID/0CUsJ44eUU91W1Lm
DGYR2i1K8ueeehRQRtfN3x6bmozFGks7WpQJ6S1jvCAX1JPyWfLLOfpBvU6OTOjvANTguP7ogBXJ
J7IOr/zaeLKwltmt2okarAdeeQ6MC0oNFRIB2709WMPSp+s+c3X51N/rVU0v23kZsyRViCl2P6Av
IPj/XPriBRHUYvOwVBXryqMCyyVLdJ9+Vce/r3Ibu+DsMqObADpNmjlYSOS+D847l8OSP7quYrzA
A4pfNSg4aMsxPXqK1b9rqLUrVNU9QviJyqoig7mI1VtPFy5Z14YhDG+dsO8t1D3jLmguqX1ejbof
G3K70TDq7PCgCqSQQovLUp4x4B4kPVQ+OOHGLxqVY6Skd/sKS5RUtK+oeHELV+qlubP2FybFM5HF
+SjiUng5vVDqNgYVSK1yL7YYDgf6prYcMgYArKBYdSsETiTfFbUcz7F3VX1rkT0AqK7ERbdHiNh+
DMXHUWaQmjryl31TekbnuYB7+cRk4KZReR+3pOSxXYvc/rH08WvoyJZaH8uktHkBw4IubEnwAkyD
WbV49u1T3Q9ZEcrEIOIQehCXo2R02dE8CvZxdgzw9WHwsotkn4G1Taj4WbdMi7Bmoj4JLzxX9At8
La4CJWjEPBCfDc2VPT1y/FpImU0m+a5s6cFuhziNsey2aIRz9S2Okp5MmcLs0xtRftbX1c63EekT
E+GGMVnNV5GtDK9NxpzOAVOGWzKDMszG1ljNMESnhcapwT11Wg0mk/LaUee0I5/Qos1sMz0utD7Z
3aFZ39EP1yXvXhx9dpoYok7avTSzy+FSzy5jtUT5SoiJTmUqjSD1KTLDqEAeXhobT1NpozjVj+qK
qr6uwoN+FdZ+dZISdoBIwwC7lIp5n51czUCc4qMCSr+OuNYPcHdW57WQM+weVG/98O0jeFg/gzUt
YEm4wANyC7AhYw9zWqmtM8gcV95kjc1L1y2Nh5EwhG4OQowxjjIQmHX2hSqtHGjtQWtZzOX1bhCW
4bug+MDLuyZaI8xPeN1IH/mSAdV/1fcllboYdC1agkYMnvHeZoIbqaFcZCsCi3//CyKRIA5qT9GK
fataAUALfZtnc3YOvZB+XY4lgNRLhjUE/V1leeOELFpCC0EnXw/tiq158Hj1YWhlxs6EbEhxESSZ
EVlJc/BUJbret8iXByA5mbbTOkOGA/TaYClaSuS90oztYy/2q0qjsE2OkPPgt0WczqgwCLp9HgiX
sLJ7OR8xF0h3aK2BUjVVN1i8VGVUlYoynKaXt3a0RjTWSTPQyylTWJ+6GYzAIhKbjJpwff7RrjE+
ut6bQpw+fVNj/YLd7mwGUNXFo5T3KzXOYnUl+1vP+d7sz/Pg+W82dw0Xn51pIXwpSbhTtMlXCYye
FjdwP9OkHoalWXHs9ebmzKrsVXbAWrtUE1HHUpd1I/fJeaLEyCw8Ui8e+mYk8k3BN3AQiEAOzukc
me46Iq1Fjz30LaJkLvOD1y/iuWVWRvdXLwZCuMWWFa4K81hQUXbzR/3aJx8gmkrQs4IgjaJ9UU0O
Y8/hOt2A2no1dTj5qYA1vJ7VE0/t7qfmXDRw1Nbvq7Epd7PYhXdeg4Lm1A/ShmJGhrusG8ejADQS
EXRnpiojdbVshl6QKkt0446oqgXS9ByJknKtUO785N1DImBI8R3XsxKbbtxcX+cyReSge289eQ24
2UiUo89Vj6v8XiJBcsIShiOolh8CciE/5SAJQ8BSPfgW5Km1iiWmK1NlHPaWffq/EQQi5LpDwYpL
Q7BdiwpZuJVlvBrF0L9gOuoDnDUFk9enAriEzAdZronxkdnukR4Hje4Vp7xvKMXriLGfAQQpfPfW
1v/3lJRRVGQ8v/qRgd47co8hsNIrJzLIiM/fRIsQ90iNBNDKcYNzorENk2Oqah7/FShXU//M5P7P
oVEGyXI7m5fNypjQ5vr2xTh0CWsa2nwFJ6aVBEgfO15EFVKLILpe1mY5Kcl+nQ5hfZdhXIl/T4O0
GC0XY8KO/2VyC47PXic2DZjNMwuRjNDV2tAgJdNPFteMv3l8D20IKwVj/KQHV1EwZr+/420aOmf6
YGR97+Ep5+2uKIoymtRCSl5lxWKREkHUc1LJvwd6Oh35q4a2HXoxNYNjnh9qhakl3dhfGLXnRHu7
OCbYzzIb9W3mEAr040XnfCoUiuBsoen2rkIWaeXov4cszX2gpMh7ta4z8qLWfK9+qHWEvbaFV2Bd
+dajPAHtutGv91R/vTGAy0BkQaEwwG/NJTPNbu7izxaUoTyDGQUSW40aK4w43TCvLRAh8st90Qvp
rsjCBF2/U8fou6JC01qwXOT2NS6eQJVcsUybUx3Yg2f1jWzzESCmdI1SEUjsxOy8blZXXKlN0T1T
/9aKjehGo5N60rY1TwfqaD9LBDse2p7Npi/1ZPBRT4Ij57uZnz42o3TBbRiyq1sYN9rPjA+w7xd7
QD7FlMWkoJ7hbEREbYaxNRGK/RyyPb5Gzg4nUdYb5Se2vXltTG8kj1Km/TNNQWHQNZg87PlP26y+
WplLvvXaNR1oF/yy6Nl2EQuDh/wNADDVkhlLUTDE9fetyVTBSZdt5Be9N1X7NDpmsEEYfw9iDrEQ
JvtNZoeMXJR2xoW/MxkTh754pED0SHubUz55Fp65NPPYpbdnGxjUpqkUXKazL6rsEDyZsy7mbvVW
dU5C/7iWkFwOpdL5lHLoZAg3GPMMPToHrOJZuy2i1STi+OGfGX9qFmqyEk70PSI44+Ho7vEBNhds
gDnimURaLdA46RWWdAh9hSPqIVmnv7lnsxIZBFZaJuPg6hLApHYiRI/qvmE75u1lnoUUo5NrupcF
AxbMwwGHXP8cQFi8a2v+GzG25hCv0fxQuzRArMO6I7Bntw9rTniNyZ8zBg1B2hvSYZiWzdl/fsrN
ytdnRx9nI1p+wXZlDsVvRhTPJZktaD7vcAfPRXVX6NXt99MziRBuH4gBvDc/wKj6ZqqoNnZina6/
iRTdLGRwnPKbgRhtxp5bAS0lmJHVXePJOKIL2qg7n5Kn9S5IFvAU8eQpiJuAEtAUHgBVEP1dFhNu
qNKK9QLweErNOCMPdPGopOQGGyz1c7VAIECU2Qko4DiLpokL+w0BMIpaiggFEjIYcifZ7VSHWawc
IN8P4Zfr4z6Zxa9yPurJIXXz+ztv9VjDDynywZ6PTLxUD4qXDFyKdfD1NUkc3zChIMdNMmRRKpDE
os0i5OlyQaAHDs3zbMAxPibFADsIsDmkgnDSlkMnbXJ0Bmhn3I5tVGORla9s4rAd0S2+ERgEGHoY
bppbTTC0p4CXtACBPvJ+OLVBKFk9iStJWNQrx4q6Ugehzw8lsQ5DeMowy/ofy4ZcPyY87ZAsvEAE
YAW/fSBCfi4Iw/vi6Qn6LaNbhT/PIMU4AyHhpOjRlqbNXj7Dc23Tentbj6xS1QJKGC8HdPlBvp5N
CiqZoNxVI/+TVUvSFdsBHx4vV5Iv97apv5kcyNeZdkndJeDi4KDczzCHq0BKgC/g1S0hH02IfaS5
Vpnlk0qGnSOakPzyPVpG6jz/ZrnHwGu2vL43nlPrnyVzDOe87D1daF5wjL+B2n1xIpB7G0Bf63nK
dNaRVEkZ0a+DBAdarIGqu8o1bUerWgZR6+RxbaGR10Fgd0v/x5x6ViMGbhYXfiikxJ5enGpfI/1c
7sAJpI2Ty8GntN1HeN8jFXMc+QJ2PTXyHLELqoAHC2RoKt9UtPSKWgqsfLKSQUsdSAid7ZeAZWG3
wxYkR/I7W92j2Ee5CCDxeqNEMMVRW8q3YK9jasBm/95bjmHytTty7NM/1w3lcGPUuDglwGgJRe+2
2gjAh5Lhv6s3y1G31/qFtivKf5KLFRqWvl2lW6PTyeh/tXMHBpB2SVvgdBtp8Ib7MnEwpKf8g2/q
69zH55YACqykg1i8RC9AtHBjtEpzo+sDb/UiX19dGk+gmPfnsKTlzPArBAe1h5auGD5TEblb68WB
8XjMegUmOjnFFI2KG3XSRlKNjmFyxcgpXmq0dr6T52IP+aR/cxHkDZDx//uokYEWpDOmJ4Te9ytz
cdXbVMaR+OzqFn+1m2w4Vpp1nrD0zfunWE4LOD63CmYh93AKD6hb0QC3DOHVXJ20mMPfAjxVmkl3
99k+xTfcWOf8choMSpKchCKpIvzI6O/pW7FJNtYf/5OemQaqpK7XSL5AL+ha7qaTf1q456VmRX55
1yePW2HerPsva9cpV2AyDsYQz/sPFOgimRLfFDiDAjWAYjN139ak8QF0Yl5AMi9M7lVMUaZgWV44
c7sgw1oejCWgie9TbpLWkc0g2U57jj1iGrpJc2ycnoO8CyanGOWHhvp0rLwJWhwWvnFmY6lQjsBF
TOe//xx20wFoDv2o+zqybUdVWjgJlu7A3SQd6aa+LVA4yWJk74XcGP0h8BkDKrA/+zVz27jcgzAD
h7khj2ra/OH4h/wFTpUwPkTLDG2k/MDl5WGsArU8r7QNXu9YAfcN/1G+eCpRpwL5ZDL/LKctb+0O
DUtQH13PFx0nnMTRY37uIEyb58bnFK80Q3KmO1UTJ5dnPKTP3rL0/zatHmmfzCdaGQRdSTPexUzk
Ju5TfD0Aj4UZqz1SbVpCwJ2XxlC5s6W69jzZg45az7RmUudOpFDhxRbRWH4kBP8S/JTEvXTqR9Ny
HpNh/hEBqod0xxayVjsDg6xWsWpUuH2y3KEhhTi11tlYbH05QexbX9IQ6SBXdY3IjPkyOWUYgH3f
vkA2i3pSwnD5TM4uz8kflzlW6i6cIrsuu22PfUakCTshtaeBhpWXOYZv/enVwktT/ljypVUTYuoD
CMZjE0SCN3ZXycFqxyLLKvHtH0aaIV02yPG0Dk8lg2ieGSExlnUHTjAeuHssCs60u1U5sf6QljUn
Eui+t9rpChOBT5Fju3LSetlEHG7yqfRgIFn2fZx6XFxPTDN5+ImKzbs+ihi1v+5QIrXoiiL2XGon
Ndx/YHqxd+9VmOeFpmWWWMALECn5pcet7wMV3I0y8pPzQbsynp0GGvYAiPcFPsBkOhdEmjRHypcS
YwUXISUSHlqWicB1L2AS9OIgTLTtkcnIgoe25nF6akbeQRLuAnbQ3BM3B96fFXIFiJW457TrkTUH
Kso54J7d0mZIqim9C1tAuKH6zsYJg9jBsPse89Z90YCbghusKWNOW54XAEhJLC0mfZCoNxz/ieaA
e4Sl2YfoY7vpoJNV4ZZkejM23aunFKwvfZcux+RtuF37Z9wrOZHLAmrIJ7Ae4VSTuhdD0joSfKDY
vzCRRHnugeh9YYuZDRcY837NWc1sygzaWGRCvnTkAbbCvUi8u+jcdaRRJZfZ1yNQgdOGv9naL+4Z
rjYTN2NOUznZUVvChF/nPncarv8kKHCMukStDJ4bqBhnDFyfKWkr7pZ5WN1NIoqjq93IH98xBZiw
zA5nikfeTGcLJ/E6uQiDRVAj1gef4pfIKsFo5+5/Zo8WzaJji2TLGcO593BVxI8SW5bQ+vYsZegA
/oLKfKFZHSOVBRm606cfSssAsGQ8sQuZc+LC+yH+St40/MlEb3/gAp1XBdMYRBvi9qERzTkmnj5y
mT+4ndjdCONvmFPfbBmNYfSx3ghWBdHU9qBtC4M0pe9VPdyPyLeGt3Fkr3xuHyk73UiGCa+pMS+U
Qh9Knn68xYzXH58CtLOukhMAMt5g7krRCax4miOn77NNGHwC2FQqnVhCN+z0mLDJJhATTmTwjGIy
glIPEs0sxnC8Ey6eqzuCGwKmf8nMooxxLd4lGj5zVYTh8YIZ3lY2KhcPKjqdnn5+AgbDUb+LwWp1
760osiTZRkeNI7mkGr6Gx8AOGl7FYCVKhosBDaKN+R118M8iD/R6Vo4VMH3QgNOC8OB4iwU1z/R6
hjyB/hjyIPLZ2yISTwXOYJ2iusWCcg6tz/TuN1KzvyxeZXxGeO0vqHTijjEnZqpxmxxiAljpaTQQ
UEe+ZT3RIitaLCQ6ASwjRYeoEYolPbhs2CuQpNK1SIofICcvXfweg+tJ75WK6oIsb0AVoKwhgEFi
NjVELbu0Vz5UJRB0fJx3uU79XgG6CtZKF8j7Hy0OYgc1lger3PzykvwKQqHTLbItTKoto5X5zdYh
rYWp7zx2uPd7YjP8RTMan35SGtgL4VXy3D5MsGp6eeEFP08rEgNnRDYLjssQE2blxGFosGBSv6DV
J9Gud5s+Vlx3XY1WicBVFd+PXQ5jQVEwrtVEeHX6kIXaLexKQZJfcwFYmuQ+Srikx9C31hhMdale
nTCxGlGtwYRZJfQSo0Y7LoUyVLq3+XK4Euq7RRQ90B8vAbaHnhtTX5wLESrkmh69QLJqvceiqD/V
uE+AiVC3rigsmaXq3wE5tXKtcpOj1zuIUNCIG1kmp9E20HT3WEMx22qDTWdqTNos01uKhfFeLpS0
tKRvUVeKmzmL55aeEiNJzsloIVYWpvGrwFgJBz+zgpU13Upq0saJadhPV35VrShMIUkYwT6Y+Dtk
OtWbDvHapvBsHE5mNA60kzTQSScrWXPTWN4d6Uz0TSUa7DAu5uwKxPQJ7/G8WvtF1TQ4KE3WijXh
iNJMXimhzr4FqXksvyBdXEYlQl0NCcRU/CODCQtvY1APQrgKDzfbImrB1Y12N4WokUpBNrsPYtJf
6n4YDPG3mqLEKWRApdCv1/dTlP9kECDAQUpuztFAasag4tQAbozvGhw5QM/DygbFSPIUKGOYzXjS
Kz21xgPRIJ6vhr2pHU7wqVO5ZFuv9v5cMTBiOADAPcRq1nFcBhIHQGVj6I1XbOF+3LDon62ujVx+
EsN8CyP3wM3XS/PgIjbXSaa3NsHS8Rkfp+rq9uw/p4qk7YCWYX8VXmizaUueeyfh01rNXdLP2brX
mFAn0qlqfHhA/WYhcAMQVpSvv32uTtGV8nzNfgDoRg7Szj/+wyDwNnjams5psp8/3Df5ULPcHfxC
L2teHCUFnyBTPaUsvgIo2zLbAmO8edONKnqq2ywMEnqCMpw5A/HSPKsLOKD9l3b7ST4BWuvnsft+
A5W+QJ67AbAjfgf/+xokSpPMI19sRNgbIC9vvD/fg00OX/Vn0AUIwug2e/DOpPjuvkWs2GzbmnfU
GbHFdOqE2Dj0TWPAnk+5CzGjPe/sFZI0x/143CU1aKOjB7TSXX03+pqB378BV7hwQWU6i9FEdzJi
mbC5TSbDGhgAYYRzfkk8blNbMngSSG8RjnlUoK0Ep/Jq7urANEMyDBsrjQxHYBqrJRpn83rWVYnR
QKJm6W56dZlc5CCWEOonc7IrI+fktlOIe+hmKr2lfN4RzdP38SZSHBT/MpzI46Ogx+WHZooAH8DV
30cYPHhYa+GfZ2PUW9UlZumCj9LFQQ4uPAQhsjvzcAu7XyW9LIzjiMnctGK57uv3IsAVC8iuwMyw
Hrx2PXdD55+TZL6Vgvsp8cIMrgVmVzpHh09UIvfKeBSD/FShTPjT49Y4sKKtBp20NL8kGcnbxnmU
ohdqZt2prfY7mj821uQmW/KifxC6aO3BVWS0KKsS6aTClF+2NVyMQY0tUb90UAT1hX5BLNMBjDeQ
WWrfv+kZVpi8p31a0CQ1WUiD3LsNvJnx/ao1oLb/VXhPDqlNSXt9XD5eSFt/ifT1botWGG9ZxaNh
MIUEJgNvva1Y8Dwl0sz7QVeWJeYcZdblk/238szAmdvzPH9JFKquErT0mLyGua9yTJ4jqgvhs5Z0
G5/eFrBgJXtqJZjPJuzIOu+XX+/NeP7A0EPnlk9a7LXYNmgbyEE/rrcuMCzGs+mKsrn2XvtlFgfH
FiDfGmWwub++09MLYmTyQcHrmy1pZhhN1TMcMDMJgqmxmvji5Q16YS6WLO+dBZVsKq4ebZroW6Ly
QjpQyxrzlkeIDQnVND8kXHPpn5lBCgf+Wuj08WOvUPcZZq3uXuKNUdrinOVKBNeQ3WaiMN/qwDrp
C5EutxqfUqbQ0mu85/2wF6pnDM7s0+nGsq2L2MOkqnBnGUDMlMX/p/cHFB/TNhixNoJe8BZPMkgY
3GorXwFgxzjml0fUert52IpfauLZsitOZfZTnXLw5tMUGx7PF9FbVhM/FzzTwsvRZHBfuGaYMNV0
d307VWk2pJhdzN/ddBODCxCIZeDVJmOTsXxj9yB/hwFpo1V0/v/J2Gy3iFFhCJPEsQyvP4/A03wY
6HtI1K5aQzEGPRzRXMqwqFt5rxHrGXSvfed3PVLf3EL0127QKVLd8tqMWE88bgx8+pfSBN9Zqkqp
uDeoeTRuef8WBreekei0F87C4jyJKs7JxcIbOZolEO/s5HD1umgsvia9eBnHpaUzWyRaK8QxPe35
/buQVlGg3EfqkbWNGlBwSZv9dV9r8nAZQX8SjwjNYcY1Y1UYe4wXDmj9a/iqN7bRJdPqeUHlFCPX
29NUVkfTJ53jwQVbPbEWOIsxZbGiAQ6Y4J0Vb7gtPuhbX7ohDvEDUosqEQy/BUHaqw7xui4aNK5c
9f4AIRtHGe6IC42wLZMy6gGQ8YGbIN+yYc3UDsDGf/DyH7w9He3+mEdR35vOv09IfdZ2Qsdce9lQ
9fobZkNhTcrfDR0L7MS3as/rZ8E9F7Hp3scQ1pun1VoljI0H9mrqzU4Fp9UuxtCHpe6Rd96++/bk
Ij+O93yNLPREs/73bH8EYUXdhHURMxFD1Ly4uWkBn4kV2i8PEiQ5vtW0i4jzFz8SkEUfs375zDvt
8kkWU9ZKU2lkn1vdSr6Q+YCsqBGljSETd/I97/ITLAXcNkl7rXmblNucmxjbO/tiUtvEvheWfo53
0hosjyxfKSexWTL0vikgnQm/nhu9uesbgi6Ix+4iIPHznKBaZ0JNGO3eOFLWnSOI/Lwrhf9pVo5R
PPulekYF/CuoQrapG5lQsH5xn+K3vyAb+xiEwwy/d24/YPYkUkVdg1RC4DycpXnFIqhVFi4hbjuy
kJIMfm7CIJex2S44MR5kVa9z0d6hKO8pNwyLMVe62fvh500b65TMvkifOwHAzMInuraTb1Qu9Bta
Fo4grkMhfzNWAWVw0uL/8iCj/8S3O7NEFvOnyEeWvE3Wkmw9y+/WwiHWW6mBwmfmBlUmydvwQyK8
2yZphArB/sYY8Fy41NS7j7Ndm6PCQN29nGkbs0O7Gksyi6FssfM0weDkVvPESxkf10brd97/yn8w
BRY/Stuto/q7fOO4tPKOXCHjS30j9V3LNsJHFhVRFneiWeTRDHkolzUoUOvhce20ET6PdA1Rvh0b
ppWA9aHk5xAtxnuU52/rYdg/zENafQURYidmRICao87dA6d8m90WabdnV3YfN+RkUjBk08gbOvHg
MvOwnQf1usTsnBp3j4LJpjjxJrKPaKweKxiWO9XyMBnFBfLErmH1z58bRGxBQ61Erl//Dd4rgd4P
lVxRZzIdjhOo0mujAQtPZ8clBDNCAj6lXf5gMFYNGGmI7tn9hBGaMOtdBh4KurfSzE6FoqEbxeDc
xAkmy4umsQx9KfL+2bKdITiZG1teTom+Z+xb9IuT3hwKVIQhjOJ+FhnDghVWhv4R1iMrw/jqMN4R
aGs96Wk3+mrv9/J3uwkLAWFQooU6lCLq2RubtjYcVk0OPhohupGY6WSc4nCio8WBEYqM20TAc36/
WeMxRn1WYVCvjrknNJvSpgMtHrwZ2GVYDDb7b/CVd06TgAMoH8f74R2vOFjWyGQVWhEOuViPdmtd
S3Q11G144xajOIN2/e7Mpzh/PsFJwaso3E+0nxPwGesMiSrZNRp9XT3Ar5fuYeNJ9denmK6DMrGG
as3WM6UUkUy3frPwmX2NSflWcbq6MOoZDcbTa7E/asGO9N61OckVYYhd97/9ZUr1lcEJExDGVVJv
yhAwkeafA43G6t1SdwezCQ3xaY5GYMi+321o3AOhaUslzgeGiUe+XIJk1elTdbjdNVLTt5VbZp0l
7AffMATR9oRxHNwZFXIKzbhPCvTjAdjq7dDf77sdr+Rf2nMAQeITThbbPzjw9LX9kK2o9ALFVH/6
C2biKZYuS/+2sBqoCK/w+2fI115dyFOxppRWRUMBVcCc15+F46uZDtMmoJPoKINm3Ys6qM8aPgXO
tZcTe1s66fjJxZ6fawzUPIPhqzF+tNDBmr/WcLo8NnWj5BYTE6k+SOAunYfnsWCdwkjyGnnprlss
niHmecQZ3inwiyeU51iT3uB5Ep1v927Q3AYs5Ko53RcGFLqpDGrwLjk/fab0wEfQhO5euS6DF8Lp
38jRbekL3tzkI7A3xly2MnLA3Yqv1ETXsucC05Bm1KTKgloWftTGKRJAbkLKM1jpiCPg6olWlBRq
bjTH6R5YTwIeEAyi+SltkMLO6gpDVmfb95QdD1SX0pPD6t5IupwBZ3Y4f7PVYb1kO+d7c8Z4NBAx
VlhGC/Lfo7Ne5MsQRDuYOzfeUxAIWh3AfQth0jSwJMS2cSUpwpvA2nnUIj79aIZIMLXtmFmPQLUM
na4rsjwlZdPJ7Xi16HkeW40oOYAUn5d/cG8vuPRbBJOOWpfSBALxusUpHthmhs3TDGIvjfqKMH78
X7NrNFcFpqspJd++611UyCwnqqcAUsCiVHY5PmVv0d/R4Cn43jZTneH1sTX+PbeFWdIeiYIkaF8G
gq234IZcQb+VXwoAubZ0qGpIgbVydfyMJ/no8EaNxcuAAznrwraodwCd8DC7CnjPPgrJa2YhTwq8
0GwPkOIUcSxXpVcTQFl20O9aWg2XJg8XEFnysBifP1nY171DJ+uq8AtxZ3s6NYP4I/IZ7gaj8ua6
tO92pYtIWpI6ihqR367OloMYDmU4Lm7gDt6q6LXvXK/f4A5oKdUzt7LeyzBQFhsErxT14Kh/Pv1P
wTCrJhorZO14g4g1uOWZb6Of37PT42wcWU7Ijcqmhi/za0uwrmctMotzpMdb+il60DODaIeRgxll
JcY0s5BGl3I/7Kpvgsh1wuRREWeX0zhUhlMe1H/dz4o/RSse3Z+LKk/LsxtEukPWGSn0Wg8gb3iy
7S/9YZIM5OJZaZ/sDQfcJC1CEbEuSC0c5ivhppjComeg+FuGMUQhyg7WAsabj2qEmrcUGJq5dXNh
sNFoxZWDCV7ExwMjQ7hCtGexhIsQEp29LohuVcFbZ1Hdt6y5Ctbj0iJJbazvWzQ7FHKXsJsIPopl
KR1HXAFU6IJJBVm3nLmMevsym79xy7vJa4AtRq5hwhhUZGw7CSJRf6lqLM7GhQiWVTbkdy672kpO
TK4eyb/NWWVt+0HjiBwlQE8enLAtCrUOkqxYOON0CfYuJTiTNrhjjNU/JWF4YHZo4ugUyKLDQqpj
+eBFoWUCTmvgQBLi/JaCb8CNjS2VCFHFTHByXT71QWa/pnJe1L4Da5DRkX9WmFvnXeyYZT73JUDO
i7Io4134/QUnyRLRdZx8hLt2gchLLV8AVI6d/nt/uvjl7b9g1ZD2uoBuOktululv2edRu1w4UNuk
9QL+W3HtRL1fQtM/KATsVTrLOBHYVV28exBT6a0alOEf3Mkt0YR9SosIzKw06MOgeRmNf+HUmXFg
dv1ZAt+Rot6eene5/Mz8Ia7d7hchAh/4qnzNf+RAXptWzmzigScgH0+cW/2s+rEFklAc4oBY7PVH
P2F579Fu+uDGqP0TrguwyN1enexu+K1H8ODpeNU+NW9bG5sn2xDx3qaF0DJl8dTi/YlUeEm5c3lG
Cpy8dimbpa2RA1wQZ8hNcVRBEA/voS97IxM+s+sBqQK7IHTNogRKSsLE9jfWER1YMMWZ5bw0yUte
Rpr198r81bBH+GkG4y5IDYAasWXlDv+E5qNqLQiAasBHGSUgX4E7J3ZNp+dmCFuPooxSFuMS8C6U
19XkPh0VXQCskbLiHR3WEpXpqfTl9d1G62QbQPe5e7DatBuQt0pkFcjalUtJtacAA7GljVmjMHFx
HVbQYmfUCxHuE3dLmQabnk/fSGQQuJD5me9/wns30XPJubGZeFRlgLwtyMJOCM9CyokHowLPhSst
Ogp9f9YukIZ15zdbtpOHK1b/NvBSJPxdovnsNI2J2tMu8hiT9QhHExkdnnZMe2MDJ3PkDv+MqbtI
f9MHVGQu1WI+HzSK1f7uxc/sMisXum/rvQWehoWPi864qxCeiQ7TxUmbVhelAzNX7YcZDAyDqnL8
cjxKBZkHyWSssOPB1l5Anvxfbpbdubv3yLbmLlOeCRk2KfkmoJao1ChIC8QM44eZ3C+qGkr5cZ5i
o8jxMoD8QNh0TGdRe/rail2vb1oIH5cyrjCi3AQaNR6sBLoHxGMwv8JDgW16Wf0XnkEzfJpmGwep
+JW81g9Lq1rsbMS6r3bqD3gpaDdT2pCwvgVFKWZ4VYX9A3WbojJmLrfvvD6V3Q1MHH9t9p9Y4UqB
qS8mmXt+uv60cwvHw+Hu7vQRkPVqET5RKq82xTVaF0AHjj1W74P3MfNd0w4njhSq9X5vtQ7YmN+n
YznLS8MxBDQqNQtnmQxjc3YDTImLAiRUXyrETamS1V4iESpN+Aw0CcrvHKMQwwBs7CDNhOX5CFsR
9mYMY/B2yOZN7M8hnLfWzn5eEDmtVnclgBdKxnaboPfnkCN7qFpDj+cjEs9npmNseRW3y2812h/h
WZ2FJvb22bBEPqxLTQyqtxLhlfHylNlJ229Zc95KRchgR2MS/px3PExhgYyP/FLdFuX1oBwdRAZf
rwrR2cUGr1vElTI08k6KhNhkwqXkKwobexHc0rgGK7pJFoHqVQTHumeunh1CRD4v9X/tc8MzNOcN
3UvgNzQGhyvbW8dR0EhQPJBhmYeDy+nCeMyHX0h26KAjcFiIOvaPxEAjngP1PVZxwT4M55xOFXmC
jbNOsE/+vnswOl1g3/czJVB0GCFUbRe4IWPKT1S3anl9mwFwS7VjIJTk+e0kY0hdCgxWJEgTdGcn
XG8EnhNR26DQ6uESbdqPyx9CjygS0O5xy3PjMwGE8UI/2GBsCGA9y1u3GFNzSqqqG41Qolppk8BL
lk6JMSdXj1b/SqMbJuDC7UXZOvU7QBw++NL/yus1c8LzgOMX7Ma+gYCE8slG53mURjaYujGHNnZc
TiguUKZbWIrFitqS4KC+hhpqlal/ivlwo+w5oipEf3UJvgmZnHa9JictaUErhF1wRD4zTd3Cssj+
L9V1Kpg0WOI3Dpine5YsKufW5L+XPZPMOtjY/F/y8ubse6NuzMd3HivJk6d2sw5Zs3oa+t/e++qu
HyxBHKWyZgdSsFWmHZQ0JwuMo551peIazvyu/iCdKxoe32J8TWHipo8zCNQ+s3mUA8X/4E0w4LIX
vtrvfrqUdgqCVgkwe2uLd1WuokjaHNEyWR4Iy0q3ygmK8Ei6HJvEGW0DlDzTAo3NNXjR1hTTPeh5
rV5ykWeckjBi+1wi+kpznBbRC1MstwMYh+kBj/grZujCj13fW9eD7Y0YCPi+uTphAPMVJYLZk6QT
QIEb0qKi5X/O2eYpvMHzK9LSAWYh0bmUu80PETVVh2JSENPbB8DBJ67nOq2+T2RlFchDnq1Bm/Bf
PrcKjzYbaXf29hDBve2MsCoyeRc0ijE4Ya1tWL96MQmuY3e9z9+cWVHePmZPIBaja8p1UI0IqsCQ
5l5pJUHbd/b5/nWnS7CjexpO99IQbyIkQvWtydTRuTggw00mXwRlQlVCvs3V9l2z0EzvFKN2To7a
lon1lFoZX8pLMSrSBxByE3fVvPszJB8K4XAUgIwuGCihYfdbofDMQvu1zMcSiayHq2MNv8HOEgdK
BT7zqVFXZ8EkiakrCLTbiGB8NhAYVEt5R44gb4Xzv59BuBTOBEJPoZgmkYoIzTsF1qiuJcq+XRK7
h2+kAeo+RjDoXD1mGp2hwm4dZp/mjgtqTrc1uwVHxUonEpjuplyYd2E6iR30Y6sTAL8nMzbGceUF
6fW3DqJ1jntT6/2qm4eO4mEs5KjTwe8ObkekAz1d80RObTwoMS+XIAgoLQTZBjApE9IbVJg+Zvv/
813TSfjIgoCmA2H210kmlBd8q4hE8VunF1B+NYCVp8Ay8yqfyJVzYlOEsKVYkAJ3fEBMtzvv6/5m
MPob2HTZLfaJqn3jrWvYZycwrAoyL+bG5Y3f05rxf3nrPkxC0yC6/62zDibdyIKB/GOnRDLDD+ag
mZyi2iIpN9bk/l2hpGJds2oRshC3b7ftcc2S85/OTgev7/ZcH6xbwJZ6TA1wRi/p8l1W70dIXrEo
Xub28jTJJJr+zuBFp4Plz/2JUI9XV6SrzHhe9RihxHPfW5/cMZGgnAGLd1NN8gKtBjJEN4amWpFd
16QxdVe9v0sf8XENiTI0S1kGUh6X7bcbDUyQ2/HBloeyVLdiGky3C+u3RIVrMiY/Yw8vKSt56oBo
eIJxkIh/BXdS99ikf6RRS5Vdb7Zn+2tQto2WwtPdpcb9jn87ZCTzpXbyJV6mvsWNC+fzrB1cf7W5
VhCO2NuKG+dEaFebEx/Vbp9Ncb/CGYRtKlYVOW1+1mHqemus1Xya0k6KxuA8PFmMdUUkjYqAZoFf
PP/p8pNkuiVE4KiXh0s086KYLdhiKC1I375pdbuXWZ3t+uOpUfWudocEi2UqC/qnfvwYXzjpvy5q
fqoMN1PKVZn7wAK4QAsyLwOqmOJLxsxqjUzkvmxrCYsrUNJtEBSlm3KCLnCPb/K8deiYiRciO3QE
Mz3ek61+AE2f/jWqQlG4LK/2y93jpAW1S0qkV8divSTFN92SYs+RoetXHDoGgCtlMDq5PmhqELKJ
0wgVhg5OuOwBCwwhOvkDHojLJQV1ijX8Fv+tMacK/1JkN5TZKklhUl4AurbDryfwPf+7eOrO/Gys
HIE6uKBn4T5DbzIZxT6aBNzxYFJLd6wPEhRTnRvqsMph1NMsgZ3HgmAbv2hS6cd5x+So/LuYzWFy
aZ1EI/qa7whkaDLNGeBUs3fC5z+7ee3CZ0JwYT3BQHCbnL2WCs0RQLlDWwkG09Fm5UHw+9A8ZUmP
J1P+JJ4Xa3RtM4IhfBbOpxtw1Re+NP0NpDh055MBtqrf8Gdj+Z0xbv1YZwdwSR+puv0mhwljyC9u
48cM0YezO7SiQzXHRJADDY+stjiGj9dlgxCzSMlqzKroDwa/EcBkOQizHD1Kyb+P7i+MWFeua0yF
5uDcWMf/sUz9tKi1d9gei9S0afSck1dSMRV/1YimwjTMpeC9MH2U/2JfWNHmcyZ6t3yTKWYG5BCT
FHWgl0sKeNDSl5Sdr6cbJbOkrKjc1ILYJeP4UgD4QsH9P+1oTdXgJnAO2oxeYSyMDEwnD3IMT7SV
1FUYFdsowbSvNXa0WxTa47JHjZ/n4YWN6XrEaI2GXAVfcQgGxXdPNF6qqwOu7en0AmQA95VIqh4g
ojnlLkyyYsGl2ToKIMhg7MLIZsTUcPb5i9x3bGzGaYaZYsljOC8qDJ0zZu+HD0CBKBacs2FGkxOG
/wJUwsDDn4WUs/j1xE943HaPoninFlSFzaSykyrEcBiQMTvFSTsRKlkpn+nUpOFAeGw9ehXOlti2
69SASC7YMfcTiSWLYQD13X2B1vEbGpxfKQ6GwUMH/BYlRk0sSVuLiAgUITuF4IwM/AfXEMG3aOrY
lJMo6tfUHOU5BmGjTn/l/6Vu1WBwFvfJdK16iTA8VXYHKF/uQszEW1Tq3RgJP95OYdH5C3tJSI8i
Npy0yOTf1swRWT2aXzdMV1/8KLnEaGBZ0rlcCVJxILkyznpc1hjvW7NPa0fCZu1hLz8vaO8+drme
LtfszxBW5xVJnp49OjrCxMSwJHAIDPMPgZUoxZ21sC2AullkQGi+SmV7KDT0JKH5BX3eLqpfb2MF
J76VAcfE62enIrxqBqcHAqHKFbwR6MEYAySB97+1QGjzLi52iRWKH4XI4G6rFIfmcuq5weP539O3
oZBBj888JHY2Q96/oYG0nAMG3MRONEnhSfGNMZPqo/fTw2TeEEORNuMr3PFRXEKYZLDCsHRQcd91
PngN96w+xOKaopuIYu7mjCX8i/vYPvuSnA9WpI3S0CsjTbAiAFeAFTxOj/i4CJGfOj1WdPuyC8/b
cEmnRRWO9raNPdETtzL5aPUWiLksYCM/wdLaLjP2otMkAR/spv5Hts1R/oXj1bnixUpZ6+mI9XHh
ZwRk3D3nFM1H0lPJ0OrIEUwsfpfFI3IAA97ncNAifFHIaddGA3ks7CsUBKPhDlNmkM1atJ4kjnzo
VoASsIlqyYWRrzvfHasXJ+mKn6mQnruLNBjTPrs5PzXS0+HZMjt/mxj3Zy1Pcbz5aDFhgMKbAIB7
ZkjVJ9ja9r2x7eouSe34jZu5svA038RANuuhhi7GRJLZrWYFvdf/38449zV+/G9hz7z1j7pZy5nZ
qdD/LzolIpmIy9m96+6NrQIUY7L6gmxUXMKUMNa9K9mYYBo89aewKSF1D+nYOk09k9eOGK6WUBCn
OXdh1/vSHP0tes+OavOCibTZeKmuqdqvP0VAfh74G+V3Kh/3rUAMAmt5bcMzoBlqEjkqQiuqbG4i
CVOi9wyqKaNqzp6nlq3iM52u1hI62H6+U46DOTxtvmem1xtFesoMd+dpcUpnzCt1hUeinoQlGc3B
2AcMHVlojrEcVoYnav2ppF+5GrtcUVDk4xVVfAIFyXXa2tTtfSZlGXhkLAXeSAFR/RabO02tnPpy
4FKsmAs6gcqDwoOdFMa+/72wCQIF2mmiPlrjB7nFje4EXhVHiZfQvAfJPFeGJEFjdyVrSczgZ8Gm
79V8cS4PD6MbKNvQEAXc2fma0WOJIdeFr/MDEEU6aMDBwZvIFk0tea0hdKtu3lqqr1pTBLkl0M7/
WCsIp6oEwwI/PCnVG+CSC7tv1qeAC54ee7LvKRT/OQIZBp9rt+ston44jWp4lVKo9vgs1IZrCuCc
HGnpHGP3GGBQ9oPGY3dWpPFuReKTnYF58YtKRnRN0GJySZC+qnHlydqJarbFzQwyWOjIo8ZQU5XT
hTee214dZMMSpFDyEInfDIEstFhGw6GJMa4jI7A910qgL7cIVyhfN6whsA/qe7QrdwlZPx4znguG
B9khloqMN65D4qd8PCLxAckNP942FGIgogA3EaBvDENf9ejLz68UqUyhRThPF6rBm9g+3apILIxz
4u6FRsMxqj94wpF5ICaXUggw74IYXQx4FKb13MH27g8WsoAgUF7/X3zEs2LPyP66hw6vks0Z/gYb
d0RzOijzl6JSbEZgeSDPcaHzO/xRwGt0OS+aplGhjIZ9FhrgjQpbTpGTs8hYxgv/G+oGEz6+QPhU
fcTHY9BhpEAYbmBjkg080ehA3mVLRg+Va3wQmrQinJELCJebAWPCNVN5cg6Z32rheCf9SxBQMIv1
THcV5PxKXKnYTDjbFmNxtYTLntGTpnudoveyHMJqmhtIrdoQcixFAiPVBNNkFDhV0728X7jJvMWq
I4gUIg3HLx4y3r3xOqqoQFiOp59pJMoN9XIw22b0GRGWMScQi5fHn+glVLx7//k5a159qXuqdYAp
HqQWfMpA5dkKTZHs0ww/UkWbMUcOzmlnJ1uyHqj1ujQF1fzwbjK3E0rpNTt6xmg88xu+6AjA/uQ6
pAyecT8IpeyCcjGAwqjEt62YNhesvAOhSqF0blmf63BGTC+VYsVZsTNwfoULgvsnPlEBxcF2rUty
zqhmnDN/YFvqDu7dftrYa6y6k61JPEL2hzz3IKgsWsw7vrwHqLWKbDI3HqUSXl2GvhNLtuA8EIot
1K5MRqrcGn5uAn1tWiycrw+HjYa8rqORYmagJTpl87R4cVIlKWj0tMb4Fr21SSdEX4u9qCbpazZa
6bUVbz6kIWk5zBvwyR8pwz4YgkoH8LzxVmnQTW8zE+PqK+CtdczWsGkXkk809SxyqF8MRm1bofYw
oIzbFjg2jaZYRplDzuI7dW7zQJcVPnOM1KgFH9FcBE4dHd5OjtgFDOP5GJOc5yXglf4Y4v8wuoL8
hXW2CQYgdEyA875RbW8GiEQE5e3DdkKz1UXvHfuGEUz6GFLkfiUIalw5wDTcO1ixEemT89AxNsEo
7QE43TL2cY3OeSwSxsq7xERFXVhTxke04u4wERlqsD6QUKyM87fcicikVfbBpSyCGCPo0zKwquP6
pPYgX859wbzYGn+GviYFPtrfvSQendrelyWADlhbe94tOQ2wH6MP8wa4v76G7FqmD1YQBlpSFsvq
w0pD3pbYhfxTCI18vBqb0eE3Y/z8OqjJFgPBpS9dmFrkRwICyliWIAT1TnMBIRq0s7HG/kKB0SM9
Lmwjq0Cs12K65BZCJ2GSgyqmJKCORYKdc60HdL69wn465GUlhSFzw4mLYMn7IFqDr16iuumgZGD+
HKQsMkICpKeT+R7a50kmUpekKms+i8ZeS6fJj5erqGOByMsdPvsUK4VGMGPG1B+6DbcwG4Sg+46R
7EJXqJW2emlxP9mGL8K6RKUTMNRiGALOhL+RIsNNi4LdlDKeGhF92QOyR5bvZXpLO561CtCdiE5/
MpLCnPcXvUB1z5Zcaqs/c9ZR/B+Zus7MOEgwyyYsSTQVEpZ0sOWxfFVZzp7/idkZEBFD0E9uetEo
Dqh+uvfw19G4d1lw3Iusix3fklheAGUqSA2wLKwB0SjXLnSA5OQg5AN6mJaWisu2TCFua84JdNkf
MvvQz9knV8rh1q3ZTlxho6O/yctjrVSeW3EzXGilVgQJGtCSMnLT0p/zRMhQVHfirsyvHLoDB51h
W4AuCmRG3pS7RuX29Nf/l8MBxdM0Tx7QtBLx+f0BQ48+xS35gjhsXJicTl8Oax3p2TXjW+OOWOsO
LAXHjq+XTzwqpPta5bUSvDLsRUpN63h0u0Gm8HIHrob8pVq5jF4b9ZRmm6wVQOnQ3oxY6Xg3lZET
V6axobNrb4rS+smFYhhkG+cjQVU3gFf1bqI0PVxkloC6VS2hV79F+moHxQWGZ5aIfO4a8I6S9Ygj
nAF4P2bRpklPe05WSy7A01ncFEgNfhwWGzlclqJasvJCmX3v+cSY2ISn6xiNOaj1mGfFqDjCubp0
Qu/zi3VBJm9uQvXqg0IuyZzUFBeDPtZ+2CCoJaltmM2feB9tAf0jI4Q4wvg0qcoOC/jh+bHHJ25J
A1aUb+c8c9co9ehLa6MR3UNADHNzMW1qssAg3SsNJKRZi5KSW4FFtxhATeTCjh1HyVveC1+OQAu9
MIuLdJrZ7OYU2IOGSMMIYS7aL6RgeCJq1u7mbnLdj7vHq+vdpSoos5VMmToDpJLJSr8B77zjfiI2
Ets8Aytzw9hV753E1MkQk9pbZ6o5Hcp9CMZZ2Twb5oC4EeOvUiotkusHfPdHyJ0izaNY1N56pJgi
FTcfAFWmBAKeLtBuc+2owA6wgufkdgixPtr6hEwhTdNk0I4jFwdbHds4rLCOuimv2alT4ARpk709
yWANaKzoFj7pJbPPWfwUPIDHJ9JDq1YYHoEJBAejmy/mXH1G+zcDCLD6rNJVCsza0mK4tJTe6VzY
Q1CUTsvRpyqZcy2oJyhwg7xrVGi02ppnI6UdD1HZyTsNnMKvtBaQ/p8xdssVZKGRw6Xk9Ynk2sIo
dYS1fnRjfXimXXgnbBRizfn2l7Oon2WQYvnde2v3b1POddE4cFth6COEYMnGNecbFBpsqWL0xWEx
K4xLJ0qtuzbUu6a6khoQx82sH2xXwXluNUL3ZBJgOi+4sDVoWD3BbAD3B2i4S9bi1Ts5PiQZK8R4
X9PECUWVnK+bnCrfu1pr3mttv5ADW9uw+L9IDt9zEFzYMvqAJaadzTDNOAfZ9J6Ep+lv44NqSogj
CaNhuvFrAGCcJx5DKDaYy7PHnr+8pbfGd4J3tbhkhR31F08bhS5Eb0NdRv/3EnHgFMmX+duZmoyW
7nzE43Tcicm1P0KjBMYMs0nCiP4xdAVEtnLmyCzvttlLHaoBo0zq+dO9pftDL/uGba32jVAO2bgc
AjiMPVjTmST5MQjMKtuH5pW8ElRDQ5v3YOj+fOUxozNB7WWB553Ijl4BMVIkopQ7CnlxHkgCpcEF
gbIOivYO6ZPJ0mTjyOlG10uFY8F4oQyrqwkvzp5B/apNocPxzFE0km41UK8VoLsGJqIUvMseFNzA
0dS6HuvEKbNL0HhhsJmVYv3aLb2FpLSAkhqNJjmIlGLK5Mrp1KeFILofwrKPQ3CbiZVcF7ckgEVR
kUmcY/WVvoZGgK2IU3vZn+6NcdyiPGGrL/9arltdg0bej3UEdCoAlKjEkORyZrD4aXKzEFnm6bEh
lcB3HWMatQVgD/aKlR6ngZBbFwX0VIes9h2RruWuHqVgs6Edhcmt3ZraJuAaDNsj3ZJABg4jdGSk
HHC613rXSCL/1tVxqZvUPLzLQ8erMYoSJESIKpIuUE4J5+2Rs0EQNz/YwXxCz7oDhLdcgzw2jA2v
thPqHEp6xpcILPmV1nMjnAW7DgZlZ9Dm+2qyl4BqFSD9m9Yoa42SU3eUnmJnrNpQ0BbzU8y9iUs7
EWiupMTvLblumdt2FepzEXQyZhW1L5vibi87v4oYc/qU41nj5F5svZomiKDVbx8b2TdDeg+MFUMT
VbVTX+Zeeoq4GIhQ9a3Iic/uiLmFbjBGMgaNwGxif1Qze//ZaCbcl0cT9z6l0bzPDtKTzSjSrekV
FlYgSJq6hbky/UgFy0XZPCCxHzmuYcdca7zCm8rYfu9jtmAEhxZiv8H3WgdjykG15r/hGw5e7sgZ
ki8nA7lVtErr2g5AxW3Mittq+Difzadk1TZ+bXFLLeYv1LVosOnmmNVXh3L4e2qiwsZJABkFyjWM
WqA2KkzEDshsCjpD1oAh3E5G541d9x4lhjbcKxJdq8BYOk253uxIz6tMahCaQADiCzqJqaSQhpEm
RiNFYM09RfASudXKFEFio6CrKFjbrNg3OLQkuR30VsjbOU3czu6gIhqUaJyy6SlWlXh11kMOO+9F
nSufC4dKIhmOisz0wGP95uziR92Bj0pPUjQDFJqd1A+gk9DsubrDkCVjCWjzqd7mJ/5kVIkY/Jh0
DRyMkTPpVQl/ALslh+zr067d5u+zsYDf53MM7mJllcWNIiWtF7DtXLDpqcsIbA+lIb2csxshv6Fp
pii9IBhvMsVCUSwcRrqH9NLZPBFd0N9fopE0Sib9XYHt4dfPXGfqidz4rpwVP/t8nOSE8iZYjYfU
JVl0vgLa18WfYMkH69HBD9CcVDBZNbKz1klgkq+1IsLZmhO/yTrcVYCBfrjvP2WeKqBv6556I+4q
mV2xHrana4B0jc9mpGoqInWzlUijU7p+eVRyzgP5UtO/SIGROWfeAv75l1qUnm/1QtvbpFze9dQX
Katt7fcl9mT1kVl6ns2m2vRVY9cmWXX3iYaZX0JFPN6DxFHV4ou1u+0cRfQpIUp97zzZlDNJeWi0
8BONq2z1IVYyudW15r+9K54hRW8BfE/vXepwDtykFz0A6C4ctjS2zDElib2hie1Za/OuReOJpo2S
tcZ6k6oIWMgqpyQ3ffRtXxb/ryyB0C8WyFRrBth9xHjnZkBtQ2STzi6+FwsMNzg6jLI8dmoh5+aP
39VgP5fGOOQgf5H2O7+BZm7QCKl6kLmPO8WO3tn2HlNne8s+N7aFCp8eZC4so7Ap1gzwqeMunptr
6A9sYz6uzNvm0s3zgFSaPTZVnJ/WpzgMyKv7JivXQjC3PT2TxY9tt+JJ7B8EbmQ/C6vf6FeMfUEa
mJ9ntCou3j4YKv6bDnjuJoYM6Gg2rm7eXKmJQtP0cX4VZ2KSv4xavG9kaGiemEzkY0lPyFwbZJpv
xnrosWKzpqF6yJrznlbr4tbw2SkTtpW3sCrWh3LM0ZhnxEp3zMOH3ZIVZu3N085vChWhyUR+Zco2
BDloz8tc134WA/9k7qveXxPUojA4NCYDw8RPh2j5L30MJz4+4Agbs0MhvfmbKr6tBnTglpoaSEf+
qQgSwbl1UmaA7sfsUxnHj0XCXM4LNOHjh+KOf9NJYA/rM1GOr2pb4WwEc1yIbcYSK679IkY0r4gs
VF6ZuGE7aCm5wky6n82GfoBsyViWlDJ8onG/PVj6+qcLsu69goEIDOJ85Ri0tJtJmj0zV87awQvr
Eut4/7mSiB5kflEW4F/lfigcMjniaWoTe5S2sip/X/Va7IYdo4Ux0tgDkGwsHCFF7Ppyhossxb+3
XmTdeovQDanvr7rxLR8Q414wydDq0+L+oVLDfYD95p2AISZrhl9McJcg+QLY++en+qPTXYshbo5K
cTeAxN773QBjjv4ZZIUOihwYW0omVCnVjTc6d6Px2z8YkOhhWRJC0tpCEmghqsn1sSeya2A2GoI1
WgqIo9niuGAZBNjVEmACRPR4qUTkSJ38vMElKzKsIuwJyjb8ZTz/VHw7o+ATuTMZI1yaCV7cjDhS
Pb4XgpwuJwbRCWQQox3lGe1AAoMz7/5oCDAXNoICpOE+MPc0HJ1UmFyTdkKx7p8yFyqJ+MdWuvMg
oWzr/oA1yDs8MZ1vtGOrTuNg5+vF6MSjQnTDlg5jiVnJAqUC5A+i71a9ceoeF3byUdR+yWctKJh6
SoMSxP2tiUn7wYVc5jFRr9bVTkKHTJOazYykivFQWShrgO5iZgnf4PCurImF9JuM2vM/CTO4viHU
9qejMmmG+3OX6QIidTcGgdQBTTU91TpgBaxF423kjjYi3YN2ZbNs1rr5mHkpG8/EZ6IzWTlPsFhS
i7WrqRdg1qcNQg25a2K+QSlXf1FAOoIdX/wLHovtKqtFE0XwlEHjrV4NgXuqCmDhKMXuO2i7yy4T
WML7rbY4ifD4M+EqrYygxEldaUF2NFoXD3f1NK+n/E5p5xsdLI4mg0xLAn8tRvLjl3KPzDfOj3c1
cxnDRK+yI6Ek3EhhQj4ggprRHuEdipLcdFhC7tbgiwzG4X/wJZRUSB0Z2ubikDDUZdWEdXXLiart
f6qDvEuDDj5eq64QyK28YbrfbwTfjSTcJjTK4KhCYRyhEqkyw7GHMK4L3veAAdrCCDNk3huFZjoS
ZohpqXzRW7UKuPPdz22OhE6OhqC9+hpMQUYKV0IK9aZz0ypqsP0iDkzrvyc8wCfR59bqOAOO0Nm5
7I4xwH8xH5STxVKiynDH/hJuTaZyZPv2ZyeuJoFV3BZCvcZVmXtRpgdN7hIfOGH37m22G/mSvYKg
mnzxBmest7Y+HRzHhJLo37d/Eswiyp08E8dfEfjPJzG+mmNG25s9O+e7A5dduwzFnupMIt+GftBW
nlV0nvyS8Dw8SwKzAelIZlNxyoP9434QWk4KEjxdF2ZE1MUJ/49MQb2NY8htifcvZIKkW+heJZp0
EklIquYBSPbB39pZQjUZHw4vW3dsLoq2MY+/x1qXwVuVi8Su6F1ObmD8dJxytrgHXMCwygpqnirx
hktbGSAc/aOM8JN1yw8X0Dp++hvy1698Jc+SBvfF1P4xDYplMOzWUzCLM4YchI16t1ab0myz4xXD
Uq0OZrVuXMktG2l8fv8dfeJwe75tL03Uzea9zGNpd6IRNrAvOkPm64pV6GYcuU5JvC5vUAGLO0j8
EtkpM163RhvGkhFm2lnzaGO7vgILj+NDzs4Smyyz9HZwj88fp/jNLGbuJyrlrWWXh8uFuDyQpPL6
kbnzWjELR3qmj8mS2ZndgbKOjt5JxUUwKnmvpsFqRKq/7Lo1LSfoXfiD1SsdRk2uJoN2UJrMSM1Q
loK2DEV02c1PSIbsAqTG4UlKw+gVSpm/qSPG1wzCA24AuVrt8uuriobByJWItoIC6ub5GuPN6xZR
fe8KtuKHb5FFE5aEPsANqg5zyB23VukAfjxBqiJ3h9AaBeHUXutLp6h64VDavucCuZ1Vj7CmtW2p
HS1N96JCYIsys7IzDBFFG2ph2SCvuhiv8/6NS0qDsBKXBW+zzzWiLfFYdknzGeFrnbWcVMlNZ+qO
a/ojAJ+sIxet0SF10CkKTD+hPBxX0qql8EadTkQ2mwZutk7JKOY5e1f2QiBoKEHxBiaq7Gdj0SpQ
bg1iFcCRcmt4t7nU+PTA5m9L2+hhcah+W/Yn4vkMlbhB7QTLC+RiWTg8+xxNO3pw/YMqNvVBfROZ
hAMHKlm8qPxvoE5FMTpnxbdTuGeZmxC++HJT8C5gARlqLADBZC/i04VIrBC1YCzisZm9cxJtZggZ
kqA4QIJpzrrdv8YrwsxzEBnue+Y76uCfwSpwCWkL7o8yfBIUbutVBgldkRZgfSXdcNjcA1/etXjL
9J0fv5oVE7abLgDIxxhFNMldepaBxWSGSAOBXtD6j4LDdZxUBCPldAlknaWioN7kJjNcPU3Ej+iP
kQU58UU23yyB3+tmgpCYOvGcx3977wrylbY/IDCllLwUl3b4gfF3hQ6fgdvA3G4uujuW083FY5ad
wl4pbj89KR39wK4/SyFrD+yn3yEqWKRfhqaMkU1TvA5JmTATpC3cilrqhCo8KuLeMAkQL5P59mTK
NyjoK2f8USZethfWQ4gOpAcpG4I4ZbTd7n+OouFN4v4UwitNMxLtZ6lwZtDWt168DhwDpkBUTvHf
VcVdqKu4OcTVg1ENykdH/QZbZ12lNuL7Wu30c+WzXwka1Pz1r2VF+OuIwGmBx5KldXG6xdCDhQCJ
5fNSjhYSssguBsG6TPcOiEttCGmKsAP8Vbtct+a1rq2GnLGrLWay5UJP6c1jeXds6TWxOU5S8lBI
fCuYuBV5TwSQfXflLnTO0876sVpgRo1x4zeLwMzQ1iNgiKXFxpHJ1ICOHJwIft95f9b8YEGaKMsZ
aYzsJkJgLArjEJaJImZk8GNb7KsLxoEfPz3Wt80T16n4A+n/5nlyjMmRbXDRd+S8dZl3dyRl+qH3
9BooDLBYX36UjlfIjLfrUoCTVV2WN5vDpPAVcsSMUdUk+oMwiY4Fki8f050IxLINO+mLUx5kW4uH
1rn/4e5dHrAn9mNLsedM/atRaODzPuRL0hAILam2/lpYRNXXyMnsrMnzCT3K+CAvHDR9q0RYaNhd
73Bat1N6gzbh8D+IqFZ4p0QoASMFy5qodKjytjppdQ6dFwmo4gqbesUERwbH44t8NsPR2wtXasz4
XcOE3gQCVmBGOUCZdv6hdBULXCVjvrqvLnwF15pM91CmNrde1lZFsPfaeErJgqLeCYvBF7mQCtvB
Z3XfzmzRNfiwORtADfCJmJLn3Fwe+2mTjvyleNGCnvS3YQZxm6cE4xgnkKFQnpW/V3jK+l//ZG3v
fHQfDTtTlUx9u0fRMnCGaemwlvbGBGFJNA6axADTTcDsL+tS1PxFkC7Pyi6niCIccYlEZLyBy+lk
TZ3cAVHD9FeSVOSsyTZxZ0ZVB+D2Gr/mzt2rjkkwME1mUaM78uKpVGpeacoWb8q/+x2wbpQawVr4
3JugoesSgmHNmDulvwBoKlXt1DZ3ClFgLpv1phDhQG6rtFd+E71/e+wlVkgFI5YF1h5B2BiMPw61
tYCfo6zP1DQaet6I++bnMt+fLYcMYSCwmsaDb+o2rma/ukNV8CGS1NrEGIMLpPr/XcbKhUT5BD7X
9+APl5R8/+ZDAxkBMP1fMtOO4GxlJZ7pWiihUAPX5/G7hZxTLdLL100DnfpW/0IfS5u3sfdMJSuc
k4u7vRsTCUjPZMa8zhQG+n+gfddE4b9m+cFggNJRY0rwROEV+NHao6IP9wFGlUXPbdExyZqOjU/j
FnYQuoeeRHkXe9cuLeB7+mgh8biZA9Y1a9FHLyEZpcIOu8zitCdKe4jiVfYENktu13lzyuFfhuj6
2e14stTikwE+ZISWZMJsxSgZ17YVJu2UB+NJbuns/GklOWGDzBd2BbgTVy7S4fOrOZRdStIsidKP
CMDPG6mIMiLdoSSKDzh3CwjAEJ3om2UJLWhufAbKfImkVSwxCbk7gm5I589lB8ov2wvqMkMXsaO9
689LZDg9Z2OAuMiqGonBAzU5FpNhKrLkYp0Mgn37imebN6mI96fgDuzpg4BDo4sybwLLR4iT7Ku2
Or6F6PVnVUwuAXp0UL62CS8RXgwUcu4vibj6jwOSPsKHIeLN+EYd22ZKclo+zPgSaL1MkMK5s5j6
X4p0INJb9WndzWndfcNcbx+MWrTrn5g16LO+LPXuh8IMBHPBDd8K+wA7SCckRNx8UYOM7R2JEf4H
uCPwQXJyvCW5WbCTVveB0sM9ZV/gjP4XM9ew2XOmq1KNz2J5kO1ci91SV+S50YwHAuiXxvry91bH
CGTPYpZWNiQZjE2ZVOIwJgQ1LDOmnmGiTX7TevmjMXfNat3KakdlzIMFVMldyZMUGnXQO28nx9b7
q/pn7s0N2CDfKJySoTZ1SLxxQzncDdNpk/AGqWxZAQOLqMX8VtSSYDRuRv4nA7XIVeTbUTdAV/wV
PBHeKdI7mGSLieCXSZbzZm+58L4WVkT1iJl3Uu7qB/XvMnEd6PPM2fK9tRlkkEi5We9y4ZJtxV2+
uquhZsjfpj8b8031nfFXDlYOpVQ5I9FFKvHJXEiIA12k1UXPZLjEemM/nsK7NaQVxsPfc+gWnMpO
UfD5TxdLQHgQLkBvEGz3N4dtYBcVzvQ03W79pE8nmHdT35wPr3OEwNsLLQtp7LCbWD53/PShZNw8
xlcYKq6boavHtagTKM8bpIaeRfXsOION+4/aHNpLrMW3qJks0DTL4FDwsOvK9M0Z2Oiw0sSSJrxl
qZT7MQQkYFT787CAvJBI08znQpOkTmlkXYOBg5spTwzxaaq+juKBHau+8zbYM4VCAlZZi+mmR+FE
d/ta2+tza0ZNpnJQoR4LEgsjl0HCa2Ph83YahgAvND02VMRXPUDu3yBPv6Zln5B9eFo+0YSmqNwP
DKX1uzi0VNxkIA1APsGRRbdzFYt5vD0MAM7LC4APpqKDApsh5Jk0F54qc+WjoT9HrYPrXxN+W4dy
/bQyds835XxoyS89Q/roNj0DonzJyhXgti4TtSirmasvzbI8NA/6BgTzdtuxFqV3n6NyZpM6w6Ko
HSmj9lUimGpstQwiHKGmpGxBdNiJ3hJ7bbcyuD1ILnJSKYbvF3eYL1SyUuUUy/lrpUam0n8OxvMs
L0kWUWzDjJtjGu1CVGkdiiC7+f8sMxnP0TUg/mA86gf+lMzAFbTi0HkgJZrupG7bWznelXR+Q0M1
Pbuqd3co2y6p5G2UxykyUKMhOlHg0tArOLOeEvAZOwFQ5lODNL9JNskFlleyluUpsQZlZGJLOadX
R2Vz12K9JAw24UivXQxhyYFr/unZ5uT07QVaD5ZZB+WcTn1wev0O6afkVGMzSaSXPseBW+nj6TG3
ZSKXEQwa8gklrs7XpAGOWuKZZF2BW9wZzV06QlcsllCpk5FNZGFV0GDTId6Kr5mfcaRTHJ7pHpNf
W2d6xqnCxtOj8iVQCECm/jO1wTJ8jVHk+V55m9ktt1d74llvhVlooCf57ht4VDnHp2S6lDsndlwp
HmZrT8S1M3BItSlGN67h4+SYTZ729U6Er1+wUmbnimjxJ0eglJ3FE/JV9/2kD7mmS+DPur9J7eVP
p9af9JeSTt8oT+egIoV13YzX3Hp76FSGfN8M4EFWXjjD6cPdOsAm0WcNCTDWvDZ3Du3ZWsxjIkEg
/A43HvDn/ol+8xxUPkLo15V/T0x+9Bkf7+bFx6vLDcevO5Ouh0KkaJSZoULV7r9noRKHT08ha2dj
VJYL5Yn0yzW4bbHtYZ0Mwiys+yrgP33Gwmus6sO8F9NLfo0oYHqNh1pVUq0vFiV5xcbAc07qv5Nm
YXArkuigz8APF+gL79RGAOPWU0oUqynsKCugNcaBxHD644NmGvGRqQLLLEXHdiZgz7kWpuWQYnI2
ndwWMk7Zhasw2nodImrsq+AbtT3XjNz7QOVZEgDhFxjaJr9W2RSEg2W5Y3MFgVu6mz5hVtszEGq6
hkYgRH0bFav8MQWyNThCM8ugrCOc9plKtlT/sun3ieurOf7ZLh8vyV13i6lnUrnJpddXZSzQAsMJ
Nr2ep7zM9AE/Qt00gUjGwACUM8RgD33CFSJgImoraDT8//Qe7y151QEx48+DtxhsX3KbZldxQwsM
mF1UvhJWehtZEWLiV87MxApXYb3JD7ayWVkOSpdetEVjaccOFLDFv1+9EyD1+ZxxNbJSKQ+MUB3R
Va0Kluq8A1xHQBdCf3//EhzyzMBz1I5uL9C6e6Oc4au7NuoXZ7gEnsWdGYXiz5X7VPVzqpkF7VVK
y/WIp4w0Pz2rCXWJylJX5htiTB8CGMPmxBG3d0Bm0qzfQe71scja8X570PLN4ZN8Q9R0lX5UNvGM
tTYyeOTJaxzIGI4bRJ8lgwxIiE3wI7h1st7PEzS1JXAoTFuP0e/10CJ/EYNhDF2p6O6rdq5ZFpez
iU63NIFvb/tWQuvVlbAoTuZH29JHIHzIa+zOwxAc9j5qVlE3glJbJGYUxhKKOBEDVtYzqu3Y5D8J
EbsNetc9EAs7L5xU/SgPmApUwiQ9Qb+ntxBfwYs72tXL0DLZm5fovaR7zw+HNZbUEhmmcvXM8oyy
SpEJ5NeSVr4hF74+8yHM4JGNb7rVgRA3hF6sjv0xQPT6dHuqwr8aPFQDRg9nyDcNHO3249yu52qJ
pL40sJKQW3nNq5l1Y6h9ausdC5t/VntoPCkvdcgbr8tMFINNLR9jHzfio5uG3JsO0GzSbVoOq9cU
nIP5EwpKquUEzV7PQ7ysnT4ABW5Xh7JCkOYFw5jkVygyQYyISqmhQp526Dpvl2LXf+Nu5Vf7Uo3y
caepCF9zztczgS2/5ayWbT/6y2hg3K8Brd6Q/129/OKF/Yic7LF+Azkw4HG0aI00rZC67AsICpPA
K2s4XkO9BVSKn3txEF5fG8MN1woc8ueEgida2i7bNGAV56cakgDmNXeMyf0SMwsSO+2+rEjcQ0tc
cZbONJU4s9WdZi8WgQ9wMdonCYNyp2m3bx5FOV2Oj7/DL2x87gIyKB7ZFeWRomcNXqb1poKjyQzF
/KxM7xQ+2RE89PNIOYtXsw5E8yqMYDlT/EulorqIybO05Lqr+lNFCVRSD2d6OkCzqwEn47DAVyy/
qfccvIMwfbvaRz8IpPxI4W2ntoJKXeEWcT11eGnqfpmd3g3dkRkLD9fdXFlCF40U0WCoemL6U6Ww
eC6h7KqKfzQ0k1h/RqsoVU7sUs9RHjyM2v/ZoCa0tdy403IJRWrtATgY5UXsgPYKuyVe2TsFN5M7
T5hcC7oI+wRjKWS95zb0GEDIlZ7mGv5iwz3x9jDTTnxZDR18pe8ntXCmltk44WCQUZboFmmOvGSa
/LsboAnUgQm/pi8y7qiRIjkVTE7LI3IFVZ6lq6tDWwr9jeH2pNeW9ZFVHlCvZHrwLKtE9RVujUqz
LyKrz7nKXQAnXWjGE7Dy3Kw4/nM+OhvnvyxA1WoY8vPjp23Yk8Y4qL8TsCejqUPUPWyQcHurJeU0
02R3Lz0Y3AQmRLOlrGpbl63pL6RIjfbWbRCqo2wla8sIm1KvHo8DTO+IrbMZrt3mvJ9xTYnjfUkG
QfpaPr4acvu9/+t67s63ydleeX1MYxjsbQ1TDAg5u9h6vNmK9GfoFeSKfsWEZhbae43i6ooyX+Ef
8Vvct0eBbVeEjbd0Il8KVXBpDwFPw3bqrxV1wYFaZG8IsXX9td4HiRGt4DTBtOGakIf3jTih2G30
xu4RyHH0zwVemoXj11BwjqTxRGwPrxsbSReJjH8ih4NEFQPmnaUhvT6smC3hR5/s2bWLZMckkn14
4ecAbkCOsq6ieZ+KJl5GPZxnMO16LPdNy5F2Hqb0CcDnje51ok5wQD+2MdyTPfMmkmOIFlDIIEUh
/lyaxWJyQYOYSDpY0/Grvc20ACG09RFt45BBljNAf/6C++Q7Qcpqk6DEyd3mh9muXHUCovtMb5Gz
nP+a4z4AObvDzOEd82VFgQuar5mQYKOx3w1CL8BzggUSNSzZzwVqYod0kLaEM/Eo12JKAR6lQOz7
KrZzaJCDQsxXdKRiFrCIWSMIMUYBxgxKUGGqb7dqTaUADb0EyNBHRD5MAJe+OYDiwSTRrDSSw+eM
Lh2IWv/vTAgHyp0mNs7Sm/k2oNFbPbM2ldvYlXJzAkrORU5XHs3Dk+f+OeFEnVPgP9x5qBsdVvxA
KW5MSygHtG93nrqqYX9p24nA7TST89thQpHtcgKMY6Hxim8iY35gkJHG/94Cj6UW1X17ewRq9hJ/
SYfgbVqgaK6RoFdbakyA755z8gtFOV+bepSjgRBeLEPNobKKcs3A/LwGhKvcGrWup1Wq2rH/ek3/
FMqcq4dfxajZOWTJWiWhUFQPcD2wmag06Dq462E+wkaKYNGVzE1Wgrn+B5Qk8UIneQn3iI6D6vTD
w+ZBomfKRs8BF0oXBjrEQtkiWxlTX5A2GkRYLV0NxzCrktcOYExvWrd8wlnW368B13QKjMqsFITA
TqgUiIAZTwlxGLEAccf4SteysLrcFmdbuIlcZKBHniktLwyBAWLMMGcKFq4yvpe8Y/d7clzVa3dZ
+NhG5qgTQYsU309Frxo/LSk7xGa8l5xU95mWp92E6RZt/pOlWtOy0wsIQIbO5pAvuEkp4jWIDSjI
utBy19Ssql2conuXpbLXagBo+74Yh0u3yMnPc3wuJnTtKy7EsPK3lXd22KeG7LG14av2xT0+G9h4
QZjZZ2lCZslZAMBqj+dEn5HBxvZ/z087CVdbR8VPQ+wIg2SozTYeqIsDw0qlxZ54Eni4dKooTKmh
6U1Z/h5vtGSGuxS8qb8BlzKPRxg+RqGJw0JU+dJTiY6jyOf5RcXz6Te2JXoyMKUZCOjUeTq4VcUl
R9WBJxl3sGbqNMGv/pORClgS1TVPHTZ1i+PyJYj/CVYI+A+xRHW2H1/wJHgBYDDHdKnAHcqPEAnk
85exwufwA1MoTZiuwwYuQrLflP1sU2Mj2MWVUFmivzYIBm5R43Be7WflrcWKONNiqLt7G7S5j6ww
jiEzLxt+7K3H+oPjBd1HxmqAMbbMyHwszg/gFjBDsdSwfg1oiYXox3TEwO4+Bg15P+Z9MrJk8HDO
ZK9rng3GPZReFDKWZm7bLzOvwV062SB/gVzF2tq5FCu+mtCA/rSRbyH4kTQm+KOzupqmoI148/AK
UuLmHV6EwQYlOvUXV8EXMxF4oeMsPyrHdJZ9epNaqA4VrI8RQ78rkmeHrjBkRtvQBkRzugT8b2oa
SczORFD5raw6iWrNyfwItcB8bCQBYh4qq3t5MRQKuGuen/yogJKVnAD3OiaJbknoWJAh+ypyh57d
XOfO2ol3rrzQxz9jBNh2Xo6TDEuZBWuAuVp9CkY1QOZ3klk5c+33MQsgu4/PRGHWebk5NkQIxAwy
bapIHCFrvkhYAnpA/ZQEy48IRnGs7x/NI0KfvE0535YTVHAce3ogdFzponF4POcATj++8tEQUR9I
2O/5tfd4Be5qEfgo2L/g1dlCz84VsJtKIvTwpJomwKCaAPzFCXz+MGBtohwO6y/abmnZzjiB7V8S
NEMdVWmGAr6/MtkCfQL8UKxM0zloTX9gJ9TpVl7u+a1WFas/BXn8GNh4sCuOmQclfBVH8dow6t2R
nV0KuyOS0QGWVGKzpBJvGBTHA3RzkzjpQjhpu540INI4mfHPDWmmO8l5M50ZldrwL/A1LeEs695Q
DaogyY8hXx1ImuHh4jD5/1u0m67Q8DXYrDDhQVOWILdKS3y3+5jaoeIBvwnk5vf+FKNi2cXHaMLQ
JFcMQcFx1/xXchvq5F1Tjs3gCJ7wRRYNgkuiUHpbUXyDdeVVY3H8Vj5+k2HN7CwaLGeC4XGipSVC
Ad6fi4rPMZ3ppQj7xaV7uRT4kiwH+4/4OFY40p1MKHiQh/4/dxQfjRvRu8OxtBo6Yj0741+T5uTB
dh7yu62BGnXMgEC9dxViPBiyQW5cU0OEOjBbyEI268b8QS3v6p2fGBloEkAOmY9T6wVrg9dB4dYe
OYNH7izJRG2WjNK6jdrS3jEndz++gSrw9Tx0YNrfcxMmUf2p458uEVBZ2bkFBFcy71OB3PriRpXN
iekvalq9Q2qbxQvAriYwrsN8nWl03/aBDVhSbrzMNUqHvWvUsyCCooXupxry0FyXfSvij04s3Vjd
9jUVxqhSAuX5CyXYQgPqofOHbBodnGMj/dgZznrf2WnNRtSlSmZ6wnO7uFJ0ZNlQ1Y6Y/s77pV1K
5LSzP3Qn87ZejGBvhFG4gQC4MAgccI63w5H6GDaYCQL80dEaYnkbfqt3Q56tjHFd/ZQm5w2DO6rA
8u6AE8tJnw6VV8sX/TqaLATIyPAJvtUjGmprj/QymYNbgWQpIne7CSydu0IAnY5i7B+vMKvztt/m
6YkpeCcJXYjUGi03yvjIN0Pqgl16XCAxs9AReHGXC+6qSHcpv3h1oznJma/5ex5LL45xpicSZ4f+
ZyF8cqp/tSgFo98GwqAEWle+NwO2hBocTzJWr1ucSnr6L1zL0EaaXt6lfxh47BgPJXvMVVicI9zU
6+8sjYs7mSkaZqHmf+RZ8PQOLu/PMf96j2ZChkmvRWR6OuUtTE/x81WznZP+y++c15hRjNgd/XV4
tSqgp5xBWYQ8uTJSMuNGLbSP81i13RAzkkdpKUmN9lw3are9moQOsaDYSEw2Y9iJE2dEGcC8UY/h
t7uM2Wn5+OZRRYc1f27hA6eJrEHLBmGip3i5ZeGqfW5xY2f/4RhW617mvSASdhN/Rp819hzte83l
tVHo/YAQla/CCTZJs80gHJ5SIQIY58jyPm6OZ3Rs1AqdEhQNDOKyZa9vg3P2oBIM3tHqS8WcpMRV
uDyYFTwxV/QfyHR90sdZ8zTR+qaFvYAwifJOvvEQYTdv8LNjwU3rWhCpC0YuLiq6lL8gPfz5t7+/
D7F4UDKFZHu5jQEz3rt7d5iQTXRPWpZYZpJQW9khezXR4n9jxVkG3ax2as9g2qU8RcbRlyL+2df9
b47jXo6lZ5qdjrjcXolJiZHgCmP95c7rH8ICdAfH0xmbXlkMYMpZ7EgYd5z2VTef1scbMZN1lAuk
V3vlfmUrCOpv7XlyddWcsnQW8Ql1DxG4PUQUyUESTS321BkYn5NzaofwTaSY2BkKmaGqS2HOBCOF
eOZH6tT/rUPNvMM+3WCx7BfDkjYhk1QlRE9K+/Af6apkWZcflRl/hekW26JyOJv7QGdf2sYEZBvi
TtzM7FKGQxVf47mspyK8yu2wJNlL5A6wBnxtHDuwgSZeVsmnpmo/bZT2NpUAVhgUAxaE5gheqGDu
HoULL3Cn+MPWs3G7vFg8THCkMr6rEuNoQsZ7bRJ0GjWKczWHILx/Fbj0m+FFf2nZDVqSthQ7EjSf
qM2bBZdZ/ls7DgZgOSAqUDyYwJ9W5v8ZSzxQ33PALwdzHSnt/3dXmryoAWJhdrlipjYTe5ElykO+
Rczw9jlY043fFiiFbrfG/2cABxAQsR2Nmgbk4ZaCokFw++LNVLs9dFvB3ls+j+JkjZRLZbY30uKz
nbYuf8coyW66EHiqT+NT1NK2kj+5q5R0YgJSoc7Ns6SnXE+BlLiS/AmOqT0CmKvsKPiOdS6qQHQ3
UizOIGN9Q9dHJjWaerSoaRsny5Q2SfkhCksom2j8tuwDae55EXcCIwlablgmWZrVyGajstzcEbyk
L12TMW3FiCqD+DIxC82OcB8kFAoS+P2B2xK0onr77UUftWPuTgfWemRM88evH1irL0c2mp5nUsVJ
f9+hwkKCfd8CBwPD1fMfvCw3KWGYTmVVSgXAXADqQ55yRWbTBg5T7gM+hRAW5t+xMHJZOc/yPY/Q
sXAQP6tqwIriVTsUemoXVlkc22QNrf5NP+KoHDWDdhUjpN/2hJdVQQk8+F6UReKbYAcA/uqlhQVL
mSZDW/dpmywgv7FbBfpoqmv7PXmgTwQroNAT1a12iKk2KzEcWFsqXunTpTcft0DjuPPGMWjkFWUj
CEZHkTzjC7s1YsCgkEtlLEbxPub8x52YLh+5+68XC6ToDWSzy7qfNw6F138ZW2xiK70LhkncNkzO
Zb22STi/9Tv9EK4OtHHpQrb/8UXIN3pB+Rj7Ux9pYDFqGhgevC9d4AGqqt5v9LAKQH4K2PKJLq6m
bvDq80OcSnTEQBFf27JTpLpIP/zbHN6ig1SR5j0LCjAY0HxGxR/WGTPOGkyUjDk52Fw/DszPwDUf
Im6G5PTvtHahJ40IEpEl6w+GXyE+vbRzNi2r/wZuweA7Hk4PQfoHh4O05hQVIpHMOB8DWOByNaoL
VBiEHxXKxZ8YvNzY6895anwss38vZArSN/ZNu9CuI/9AbSfPyJT4wawP9Qf8oqSIMuXpAOOd2dzK
qmrjltyZ3OSDUHAcV47vAbLxNmbZT0Wp2z7Q28G+PVgfsqXYUk5/0hBn9Y16NWjF8zgX9yuTw1NL
U0rYn4qE8+0Uj52+D7fImkL4H6NZ6DkMVoPGsHozOprPGeWagOp/+udWMgeIGBtEAt0Y99pR0uvK
PAKgCqtuDqWQhbRcaEGp3GdDEDB2pyltgOJLGhWSieBJsxmWzNOtRocXJ9+4kzy84OZe76CD/8KX
EWJXULcvTA1+Ih9V+S3tY73LMVpDEBhXmaYgLs/Q3QzR6pgm6k07lZzOPtymRxpUMBujk/wUWBfK
5fAdZ+IvWfzWICrcE7pNbOrif8m/nUnnyR+46JXKYUpO+FtZb7JJBEc/gxjCkDJardKt2xCGI127
pSf8qGUxreFIgSBui+S3+RdX3QZWpz4w+YyjR9eS5jnx0v5GQg5/gogHmEkwMhqpW+z23QArVYYS
DqZEdvyjS3riGiSOvSZSwJw/58nEC2jiuYMRhPoQ4CuUzqVN4F87MR42Ym705UtVvsLyylHXGu1z
LmGxThwuMxfoFJ1ZSPCShvhBMGtDK5gxjieuRmWJSOo/bj0VDgz5OR0WxE61lonhpYKR6huGdKdO
pvetqlA0iQzccefTDNeWWRo2eoSF+dT3KTlJ0+u3dVP2BS4/ASTpLT3p8E/kebnfgmjvJlZWwWxi
R8Exw/5AqwptWKvMkScL07Ml8Y4XA4/u12XL/nBpLHDXtpy4uKEoVFTlq2zDomGNEkCg6ETZPkHe
vAaY7BGYkF6QyuXm1hTHyFS9r8qPZYpkurrWYh5puDUdISp1IbASbYmMCo+/rwnpfEbGp8714Tac
4tLHCsKF6V9x+9LNNUXZ8T9cqE48aKXMdaQNAgK4pXCLF+zBHMpPISx/hGZESvnqW4JGT5BZuhHR
V9xLxLgXSS/xlcHhmWEhPnSx5pjj2JOCUHCZa0e9dl7FhJFM0bqfbNcCUxNs+WI2csGIn0gX0saL
wsI52c3+1UWlx0/9UJy78lDSw5emkBwtlXfKBKv8OLMi2dt3ghuEbW5aRpQHquxLjJFqFWletGeS
Kpr7KIOkMyZFBza4Z1JWJwebPZhcK5HM1ZZvHI6KcaI1IkPjItYS1mPe3eMre6bZ/SkDzl+7MhAr
1AJRkRaRrD6BU60Abfby7bDm2EPAHEkeDNfROtmXFJRg3bQ4mWeQpa9G/sj+lBGkILy8+Cah2bTL
UamEDkIeMH1roGlOjpkHkThZjZOp1PoOsTjEGmiJACKOeMHkO481eUMRBXUgTsbpGoO24XJuxrLw
KJwDZHQeJG623gQN+6zqkDcYfGgMHIYT1cczqNXlZ3ZxxzFoYEwuAaY/tXIsSvd79c/wHNf9n+Rh
xhKiF7fFlF4BiSGMBEeOHZ1sel+5XW1UGtF6zFr2BEici8iajnZt4NALw91HJHeTkPC36GVOWEh3
Fj8962fpO0YV71LB1djZY8HG7SHWz8kmIRVoFa+Ughp3kiAsvQkhzNLScFSOf7K+FuA0qL9LhR4l
5Ekj9asInvH0DP4bgv1CBOugg5zNjda6znESoAsR+G5+KRc5iTG7W7EYNSfMJUD5ahunvubWq05R
m5cFT6ekMg9fVUHkdI0JB6cDJIVfoTW/vWTKGSxLib0SVdYg0ZxT+9CIQhtBwtNNZXjw+ZHAILpm
gfozISDs7wBt3mtd+e+lQMXJlfHMg1mhpQASJ7girUHCHpvKScmePGEi9+a/Exkrmd+MVhJh2vBu
J6XdbMHn7wAlng3SFbhpDYmqz4opanjnZEo6bfUax4k9qYLZF2ZkiHo4I4zMU9bJKf/DlMapvsPR
oSPrFA3VZY/hqnFd2bNfeCY3S9HfVYSNjjGRCqHCLEWfex8oZewxaphJg/dLfjTqtvot/HQgvaOC
X97QmkKI8fIdDsRGdGcxdBekACGg7m6OWOIVzr1NuGTcw1Z9osYLRo+lCxTVjGW+KfChF9AOmiw5
Y1MnlhP0+lJF1efCU6yIgwqEIYk8l8Bwv9SlEZM0Pf3ZvmyIBV+ur9hWapzfMo50nD0edl1hCsSB
bGlOXpq6ceRIBn0Ap3f9vXSP5lC++6JEeHKY51DXFJj+OfS0S+MQmKTQJZeXWihq4VsmIRcLOebp
uJ74cQO+wThlmOMmwfDuC4DYxvYnSkhtePF0t4BcBzhqkPIs1pLQRbLdMWv11GqVZjmkOIKF0xDT
/1J0lkprzU4yPnb/GybYHwY8c2sV2mPyrC+JIBWRm0pyZ+vx1aD3GY3RNFYnkEDlmEscFbyIyFVX
oQEqdEICkgy/OGugESdu3dbbzKrodXYjdWAcxzPy6t8Lcyj1kzJJCDZ4DJsh8RRVIQ7k/fMutugr
WRw6SqzcvWeBO/BaS7LgG3tP/aqfBCSo285o5aFvFc/UMhVFvep2sXvzmY9u4moWLB2hSQv7aGJk
koIdA/dUosJAvscNKjxFGQXTr5hKXgrJaJ2XPvQbsfcDTCzlFovnpQgnbloTOpv2WjdJfT9hpbKn
kbLACKJxgsdeEtC5yVFl3ggReyxe+ccy4H0a5jRKg0HxTy4UNaE2+ImnVgrLJlRv62DQ8AIc4iKF
qjupQokLfHpLoOzkCzaY1tIiXXTXGc5wBTJdWD34jOuXfDO+8Jtari4T1i1wgFX6/a/8hOqU3scU
3QlC0UOmX7rCyhupsoA0sZBjONRjC4YrfEfIKmRRew+JY7YcpM14uGYoyrUDO+uKfWDIff8iuxVE
sUiqncJlh3pTF328RJtHc6YmqUhRGU37UcdDsY4OlKMUmRjrlfgsO5ZMegD43zf5RH3fQzyYf8cO
ClZkcysTQNicFov5nQPG/YaGolnOqUUozzRrqf/lwatSSui+RVlYVHyTsc4QeHz5Mw3aet6A2n1O
NLpBzz1AFz/SLQq5KorzxsbeWSVvpKDPndYUyb4npBhOHBcwsuE/jmDYeOGWiiQotYj6aLMxxfvt
B8gRwawLe7jBEtgseaxghEOaAz1EOTn0KjAghzFnZobUM4vShVFWoDnmGE2Vod64Z1nGGI0obJgT
2vVkp2R6TPWZWHQ2VEayYRil4o5fUzflezsQmlWfwcFmkPmKwBV1xy9Fev16TGxYOyDmUBdvOFjc
wNCDporJbdhfvas2pV+82v/z1/6ltOCdRGzGhcVHga1h8ZLPFMkTp0Bac49CjyyFzpQ7Zmhevu+V
dOhWU3D9Sj1//hSvmUu4jqD037242lH0M98asuy/vsy/kb4WVxv3tRaJzg8pmxVr80gx8Xtt5S72
pA8kdI0L17blTurxBvNex7UtGKSDDSEiFV+UskBalkZhg/ylZUCeYJpdWFJzmpsUl+EWkTbRFFDS
QtdtznFPnHIYDbKaV/2zmB6kkcfHbv5UPkp1Z8fM/lY9mmcXqBxDMCDLmp9tUGCxvOW8+W70N2i/
wxlWK//OzLSm7AOQWdRHFun3sptm2UxIHJYbWMGXXBryeDieaT0vRHMsQywUsl02L1oslB8ecgyu
o8zmHdSUH5g/PaIR3KQxAHUdwHB4ZAtvspzemoi9QAetiu3ExsYnZAZdtw1yq71CqBA/eXg/yC1W
yk6bl4TQEZRfm/em7Wj71fQRCCBNFihsEyVQESK4kssbQMfYzh27lF5lO6XCllqnytjk2+OGa8n9
4WNnp0hgHB0dYaxOcjBQausJ74qA0BErWeL3KML6sSFYTo9uMB6KQOYdNmcegDlRMyafPOlr/sDN
nwhTRi1yZX9yC4fztt709gzRFKOHXQvYIY00YfvFJ5cQhxpvawrJI254G+IQLk9ga+lXF87oem+7
Q6JjaTtV5j6grBrlwvEcH17RqC8G8X/D5XZ1qOm0TxUCpjiYU0ebiPYIigO1PTs6K2Kqj2MxeWje
pHuag6C/9RZtgLawdPLN93M/Q/zSUokYmAfdxGZ35G9G17tuVNWbEn9tCRV9JetOaK9TWh1/zFbl
8dQgLS74+9QLzixRzIy4nXo65ImpYMsGiTklcfaPaSQUH0gWJgIl/EOff/jZzsrxSnrcflp4+fKo
dvZ9F+T95sBrVhrp1qUay03CYBSWbQkvL0FfLo+Tf11fCf7BPLk2aPt/Uu9nAVpPz18vWdYs92ct
RSVTyVIHtpolqR7x+3VG8TzMQeqolXddy3TCSwayNXST9CUsH3esLvi64KildI3oMJZQYLxUlJD6
r+ItZCu3BIwOrlq3WPVlOjVcRosQieP8OSdfVWfxrlaSsXm5ulmx31yBmuTp2KirKv8SkbyD6U61
NNwy7ePtA7r8ywHOKIm/YSn39O8w4rMwOR37CAIYAv16ESJ8LykQjlwVHXw/luMjF9q640vPSR8x
c6XFdDvOA2JgbtuJqviaiYgeUSWSQwvrok9zyYaPOIN9u6zj2JG/Dyi0kRZ9YTBqBYURZRWMCIsm
DRZILLGuSJyNLXAQR+IRMiQVrC+zqKdO48Bme8p2I7HhtwJoFPDmL4qlxDERvOmkLZxBPmL7lMBj
TPpBm3TbKW4htjx5EmFJB3WzvMWSP4jHAOoV+IBUXKtM8RUBlhK8mszVM/6aKAA00zi6uQ8l0ffo
gXOHLOEQ4aowkkbjtkXldjQpfoUQo3VWS4fD7gvTcJG+Veta1Np1h7Z7hRVEplwOH2TYFmQsG5bM
dGatPltmwd6bdpStqFiM45C8M8h0EYUFHepm1Ths3C2LdkiHMSNRREk1Z+nKUXmfxaQLAynG4bI8
Ubp1eob4eIeUvtXvu8wUD3voFFhHPHe1Hcnb1otaFGfALgXC6OfOIqR/v9TRQCqY/Ym6f6spoako
zyhqLnKs/DZZq//FhFOvWGoDp4VjzxyKw27RfpdI/1XGT6pZO3DrUYxAjDtT3q5GbXQ+b5XNfo5W
8DxVzzuyTsXb6/fIV9LAnZgdixmHap6PQ4PSoZBFl/WGk0Oyz7wLMyiLl7xbb4mywYKV4yI6iXiz
0Rrl39vEFBdW3+30QWzj9dU7GcN284KZErJxCsIVL4C//AjBdTGLCA6tzV8qrYSiPxkWxYwANlCs
f0PWXPuyO77EAb/PIuKYOETtyjJEQ2mni7ihNvpcuT0SCevtcUr8Rcvzv0qJ+LUfek0IFMPVS9Vu
XTP4x37QVVNcR1CuSnOni2z2gntx4/ennHZeF7fPlDRTIZiC1cDaaOtkMio/ZMiLg/1p8DqDJ6g1
VbOGd51wuNEjBIxjtM9SF3h9BnhByjEwxFlJDXln9HtWo38Wo7T029W6vrrb+9oYsqZgj6+uYHBu
s5YJfxQLqBInfzIITOFz1ftAlxbdxXtlzxWmbgyk5cTP7PEJQid4hZEFOSGx5V1FPS07vm17ClhZ
pPCGR+RHBAUDMvq4A2O5wFapWhtKxW8BuRCdeWdmUYTeAG6/4N5pHcDxVHcieT4/+gCMJ/xstX0X
I5Ly1X43vIf2wtr2IFZcT7/kiw5+uJjAI740PnUIAsE3VY3MoJhNb2TLQpP0bT1J/+KBwQI0Y5Fs
a73Z9FpCldyS0ZnC7wZRdVEoNC7OppBr2S5V3yxLHBJlcPVnE7+l06hmC3qMSgwiAf+g987dzRee
BO0hCRVQaJ5wDLBqCpugddBvtVNdGn2uyir0PrpAl+4jhNEbPTawhBxWiTkAEMRqGD8uhYKjioJn
EJaVLjbdsI5rw6h00kdxmUmLktEvjkPYh8Xr9z+3pLsAhkBdWFvmPU/9cN8YQI7KFhZMTafqsxGD
wyRBePsNa1+cobHnOAZPgOpbk/WBQymPB1Edh1WzaGX3aNG1sUK3X8S+sDTF0UzlmDY120Gk3QB8
RlWgCnvUpJnee8KeRmZErX9BLRix07oVRq1/iMzIrHz+Pgvjx3q7bpPLfuREqJsoLnu+EN+DzFHa
0aE0oE9YS1v2n2mIRdhF8ReMpEC2WgxxU3cGxdMDjamQ+Yxzu3Cd3wB0IOataXbtXf5RZCgyPzSw
iGzYlo9e6OXug1EFGWQ6E/LVjgOGbZyO6jALq8SXgw6RO4Y6bU8zgaPd4MTeEmhAI+jf1VoJXWyT
Te5f2Ob/UHEDT+CVsvdm9oR8RnT/GcuwH1kvqGLWbQbZVxCviBJ+jpCm3fFuRFntB2J+viZPCvHV
4RHlYJOVv8gUbmc6wysTVnYduA5fLb8+BBXaf8DP7oP9dyvJQIoVf5Y7u2RBkLd/vtfdYKz6tfZl
Nd5IdBRJAXGL92QI6vs7w45fU2QOLbdD3KKzIQZY8d4VIDr7g7zU0LLxA1fNvz9QyPtLzApRpMaD
2QBU4YUUBUesHv3GEdZQpYUHuHVCj4pckrxbxnuFK++wjggLMAGLi5CYczbBYs32Csw+RPYZqZHU
szsc9ziLSUnFwj8+RNREMPbR/sWWvntoMFglJVzL9N22M2LIRXPL/dEbz+JTmsXCSFQcokUvKv3b
rnhnorlG0HsyJvyaP3Y4a8cO6oV98KnjL3zwE/FI5qdVUtWtqglpzWz0xvV+PaGWdSEkYYXbSa6v
9VNoRQT19xnC+medwOX4W4933ujVCNgDVHndbriQvrj+oO2pfnVp5kq0YhT1gENr3Gpk38NQcWbC
hNHOD7JJyQtLkwaMOCAVmg25XmCvDsfQj0GHdSjccQ6nqo+wGHJFupTj4Px1T3HHyrwHH/au7LTr
gkmz6lwuzPnAd5dNUczU4WC1B0yx2nD9IWbxi+Ja+sq2ggwF2oqu/Hq2JnLhaPUoVUrMVuC+zPWq
8Pf1/v5/VhTGpzFqwfCauCgS25G7O+s+KOxQO0mdMUsNc8YoU1k9QxO6kLU5PCTj2giCiFzpYocu
gn9CDFW2+Vwg9cwCUd2mh6ZUa+TYXvRPcqSscBpieDYx4axwT1bxdq/tR07y36Hr+Uh4xBo+WvrD
j9VHG4AvmDBdCbRncbeP1lFwE0BYvk2MWKUx60LISegfM2m1lUv3VtqHgYok7mWUD9NnSqwNVSfG
Voc6aHKVseU0OYjhowz7TTMSDwdi9QGuXk+8+1z9fGd8KmNX0cp2C5bIKc89Lp70Xl+etgKALJoi
dXbmGq6m7lweeVGCStsvd+463E9JX6AZkHXCvTqu/P7h1VSFGYimb5Og9iU4PX9xmZgPVis0kZZu
vOYnsjoY/CZ1hesSvVSiVGiy+kzPym/j7ILvQb7SmxfYob8VjxIye1BA5WX+XBgid7irRHrs9Vde
hgSn+fAtkvVIEOlJjCLswV/3mOa/DBmlB3YVDN3I8FOMUarv51m1xG4eu3BbS5tm+1h9smQmcFqK
Ov5AAw4xC+AcNsB6nJ46jR7tW2X//7rUBd3ojL2GXHxFZR3QOqqwKj+kZkqQ1PlQ59UKFP3jD2F5
SI7p3AUbY4+xRCbmTKeiWsowit7PDIzMzfYQc/wjCjesm/MwSzTcf8qN3HW4O2w6ZvKCMNXJbjEu
vdbGRAYmnmymDYarSTCaGXCKjG5bMPaRpG8wbMVtA7SnBdSVJIlK3guFnjzyq5vvUuIjImrR6zZC
8OsN6qamfEcfDybGeM5hHd4qTJP0JHdBtdvTTMUXczogJX30+h8zObNhbAYwspNkgsV5e2ZFdh5W
fsJg+o99dm0ddi02ETvYacoXMiqsnvpRqusg5RS0PlmNqNOgWJDUQHGFEu89rvugyn3SD1GBw+C9
Z0acoe+Z+jC8B1Q3rt8fUlNvGwtbkEvnCyCsDh6UUBQaLtCDTHrChq0Hnq4+hseXZIsI5P38WVZH
bFfuO8MTgvDhJt2B9d9NnUag0e6yEFv+wOOUJGIjh7MtwhwhvEmmSIhIPgWbKXPYy0Jxa9VXgOk5
tbqk7NRybdotYE5UMHi/N7gDP1PEPGMYDEW1dLlP9DfzNTAbqwEiwcmEx9HMFCMlRncEUgrnVV5q
eLpWIlQRhXfgcvCed7ZPS40BmXsKmCFdInjQwMWjr83Ium/sVfNVuzQTyKYc0bj6Ki4JuWDbjwzq
u2thhDZ3Frs0/ft8xwvDFLgl0iyTYLcxukg3V/N6+FAfeoxqzmSkaUoN62MXIV72E10bEfMzIA95
R4TgzEo4iuAs5SJxzWWWLhVlJOtcIa5T2MG5jf8go3zlrpNxSjK6gxNBb4YaaI5URlGUdaeSiA6V
CAAbiIbxfzLaun0E89EjvdqUCZsZiW4qy7Rz+C1Om8VKEdCY/tjf9UbyldCEy8JqYQFz5zj4pH4P
xEbaluujQ9UEgW0t2+qFc96IXiCXInVuUP8R00cezLsRRpQXUZG4WHjADPzMu44C09yYJ8gqZbhS
52ig//A6fRumtKq4P+1r+ABArjTJAIYM4gOxihM0NFrCtZz3u4lEvgVNzG/gb3pxMolI2ODZ67+O
hspwNcEevfY25oYJGkJ/Gr5QB/D05xR7sS8iCENppfp013tQci0k5UkziPt3Of/e4oXENOr0TNVR
aI1dD46FtAy+Uz4na+8TOQSJXZ1Oo8pH7k6DoS6YlfZ1ntTO0N3EXs5cCbRj8bF/yG9IVfcJ2Gui
PViD/gnuwhpMu7EOgzQDnf73mIvgilgHu0VcQr9gdXFbxGbEgfMUXxuAe/XPAE6i5eHgeXLbTIOQ
JAAP12Y6ZZwbyE2rYpumDVqcK6nNci5B/7XOSyHEeV0kdPd+geSHTNHwhuD2WVfTuCycmWUkj4Gs
04CIinttg74fZanpGx5ZRXFbyyk8rzCmYA79l7SgHU3tDVYTw5xEfMxEUXLD58I8KHhZROWouFnv
355mHpuT5+Pwqeu0qX4KJ+tTXX9ZGIjppIpGRlgUsY3Trxc9Hvoqsgi6Q0AF+ij26Mt9az/+DCjY
yiZRozZQ1Y9c/TLniOr65QCwuui9YtnurcXzKAFAmYPB+Zu33dBKfdK7kO4iAB6ksbToY8yfOAkw
NkHgLmt77KsWecccpDVRGuGmFRPKY+bM0zaO4aZDlnPwzTHaktQwYqeRaYG+6dqf9Qs5/3SpLPrn
OJwvBUctfOYeSD5lq3CQZl5xjJtFKitSw4UYxEGD+g6p17tgI4im383NqEod7flPyCh7gx+Xjbx6
mLJH3IPi7PqHijx2G8oFthRXTcpL87bddqOfUkEzno8lik+UrtkMxzn4h2dypJz6I0ir0/cWLx+j
sFPeAwPrn7iOnkrjBJSLHZrBwf3hflGDp8q2GHxUEf9Os1ZYHZDmhccdeSbBDGmZR30RLhqylgd9
MTQ0zZ7nNl6XLXp75wFerznKlXLmVt7dFQSdjauacqwIq4e+he3+DRTewEardAh5DB8QB7CV8oEY
POpBAOmpLZAW+X0+5qFLQJEITxd5AOmyoRj0+KoX0GNnjn8eQHLY2zfcQXitaFluNlHQeU4seyIs
dsC5ZAgvub8Hc/d13T/Ol5mwOhDO34cfmda3pnwaohlRFNQ+Af/0oyaiKaNH022gXI20Taf/OuD+
/4tNsEeP4QqQsGtp9RucsnZcmL9OpfA1YgRWfs38vKkgv/gWyxFg4HRlpwuLwZIX09g6K+DFbV/V
NqeV01qkztUKqsiCmZwlBJQQRNrzDvmAEVVi8KsKFOU00NpvYyzL95Pt+bwWJ3zriaOu6X2Dir6t
zCOGkhcZEEknhjnXulxqNJQCgBVhQbg50z/lHireq42BuoJIaBsnX6gvTajjbLx9qVc/XNLUQVNu
sbZchJL/tGOXmLcujlO4bO23rsHkztl4QMW+ZIzILTjlfL0BOiFcoEng+5vBLJ2RbodzpT7GBahN
fUtkHBkNmsUy4ZhZM1nwLHmIyuicc8KKLMI2IWHbwZToxoaMfgqgErKp1Ux7WEaU1xX8KsoOY0NC
3K3CWW5RZcbDxlyYq2qQBhP5r0OkwF5kSQfk9/qqQfariU3d1hEfA1Xzb+k9xYeuWPcLNjsImf0T
N9f6ZHhCP9W0q1Tx7CBIIHe4NJfhXhAlXT36Uz6gSkUVpvswnqg4sbIHLAlfV7AXjufccUyqfJJS
JqGs8eoPLlD4vn19Ia0R/Af5cDJXwiNnSgWIYpVis+ChAk1okxJIKWzK3emKci63LCtgbWez8VO4
hN6OhGmgI7V5oQEvmKqja0TOkqJOsyggTVYtatLJRVTpJOrcFIn9Etcfp6rOeHLB0qZ8BJip8bf+
EHQN4h1GW1MNhQ1+En4aGaCZfsEyMRYXSSS6cQwkJSwTlgwHKHX8S0icUE6GHDtApt43idDD6gnR
b7pQcjTvTDLsGxoP83ORhuICHeVPH3r0nxZj20S/cWcfw+gOYj5EftmMaXnxtlmLpjESYM3fpKTb
UUeWJtxpytQjI6svsJAbdPv1PpSbVWk6ZfW9DP65GicI2WyOG3/rSYljwGlCs2q/fON6kMJhjP3N
oK2WHPvJdgrHHgyBD2A2rO6U+y2Dcp5E9054FUtOq7wLJuKaraQdr2crXRTfmYeiLh86KPFy0A4q
PFSU5ADdK96l8rIGWl0cLNmHfP50/f3bHLWdGouBsgHDUHgH5INCd0Q1SuZxhsMJ5qvoJcGKqhTc
rdUIdx7OGC0x1fOOA74mvQXi62F1wR48qyFjvOCzQuClrIGILhA+tsNyHxjgXa6c8BrcRwAR8NFc
6xoGP++dJZYP6llAnOmiStDQd4XHPDZPk6SzmEN/T9Tbehqpv6XTTbzA061Icu4oAo+kDnAOvPwj
Dunw9aRtwIQqRuwAwHNnCQG3B2Yyyp1J6xxHPykUd5RWDGnKYMStWLCeiE5mITM4oU6Mv5Qcl2w/
fOyuEACndB5U7tK8CYuKt3gZkmwjdQv3dHi6SkmvJWmKhT1KMVJOFiDSkN2v/uIhPwjouMolzUR4
x7HqNjHiKg3+qJGvtety432FRZHjesld7t2vmZZnAzKhly36WCqSLYtWXFIU2EsWcu0XI55YgNCo
AiJgbfW6+fsyAhd7MzmGjag0c+dLbAsLofkb0bZ9AH4B6AUrpPHQXdTD+hqrB9BgL7EfkBoYRUDB
PhyT8/Vdv75y3uP2bRElJ1REVjVXEHYX1tNgC5k2A113FPp3lhq47qqaJr1yRA/zFGxZLt6icy1u
/h/USS4CdCd8oue9NKvaFQ3dHaSILiBG/3bnnRuNok0KE/AxbfFcbmogvzbjlJgCokpc1p4ikx1/
ex7tz/nRpwDQHHOmKb9buoXWGa2RoXUlEGKSLq5Xex9H/tLCxoDYQqySEd8Rx7XBOc5W4Q0uYc5U
PXckFsscNbmtKstd/uP+Ovax3EGHogXWA6OBfysaQoI4a/YvIX1HQVaRiEiBFwsvvhxk50Ym+Hn1
hbaWMXcnTa7NGdUfBGAJhkAVfrdKSauclclBQ1NVlpkz+Y/IBnZXNOaoXLCDaHUG0PuK3/LF77RA
eUFBCYRATpaBQLIOFvdQINjgHRHHO2KE7RIoLc0NI/9YMhfDXe2iAtwAr8WW7oo7NXVMJKkXFKYc
n3w4STLn0B7T5U5kEpQE0NQwZlHxCl3Fm+Pd+76lxKIFUfJl9BU65hSv7RlNYUQBZZpVtb+uJ0yP
kcpqAsFtK0YIPV6d7w9nPXFoEqTlQccf/7mouNQGzRGTkIHDrdnL5jNWBTtZL2fxbQmpI/zxp0D2
wQwphewW+h+mtEiHIIOhyxehTsdIAf0yvRsB30LwxjnYK5BnnxmvpYaCj/rpg+ZgeUunq1rIaMe6
PkJx1/51F2Ntk1wSz7ixhwrwBs0ky/g8fFk6tk7B0XHT8NbJtTpd4Zed7H6eZqPXubYMYyEhEA4L
jUUq8p/gq2wBzGwmC6rlvPWUBvOOsZMumRPMqr251PYdnmQU8ieMgyOs/WS0lIc88vTwgpLexz8g
R649ab6gYy9Jz7a8ZeeUw2+DdfhyJRBtMmCppjJn7pRrOCt7eWtIPAArPYne7R8otdE1Lg1YUZuE
RAX1UQTA4KPiIHOCOCZ0usinQETTuqfRvFRCaewU3YjqfqLB+v2xvxrZNkp+Wd09P4sz21HhtKUm
7evc9p3cTMhp9jatjyE5Mx4h2WyZQ5jRiYzqtaIykr7UbQA8jMWwl4zgZCi86gckeZhlqIpjWuet
yFQI6NtacPsTck2a5AI3VjfvlmWgV5z6Pa8XWo7wcJD3eKVV8YT2kqQzHBw/mWqHMrR4eUUl1OF2
WcN/fa8iQNS/AhnjAaDQAvWkEwncm9FscGkGEC+kP3YXsJ2AAVd8C/7DZOoyzuK06W/IUWh1+8xW
TGWjOZZmM1Ncq8lpHBfxYD4D+Y/rxI0OelHJamjmqcVL8e299kZ1sba137LOqNj+PNH/SbHJlH7C
vYtBK00pBmchtu8INKTacilFVcRbLsUJcQM1h2R0simCVDGHZ363ATxl7dfQff9NEubVjsA4aDaU
b1T8WyWnkDQg6RsbO1+YOuljseOqMP3tozvSTjZhIziy108MKYctOLeybC44hJB86RpmNqvqwYzs
WCTVOEEhpS0rI+fyTvq41eZno/dI+QyZBLLEDXoXSBMmYpFzKs2S7/pTjVDY2LE+7RoUJmwTHQ8S
0i0k7ml6tuIWx66F1wee7Y/vxunCkHj5LsrNIoPHR1+FVDvt+/hAmC51TbMfCVSItMc4yYKlpDWs
NtV+cjVutIQfhczPYQYjOiqt1YFOKgwhuaTwFqCfsLXpkUEKQCEqGCJs9k//GAo5u7Yry6fuR8Kj
MA/BcGDzlAILLfwtfgz2oDcR3DZFTT2TKnRzUU2vZ4EdpkjjWyy7Pc2LN+FqmohCyz2lYpkV+9ez
YopVKMBrwuBVeVfPIqU4dZqCLOc+Ikz0yVcoK9KsYXrCpQ5W7d5LgUgdQgzAsN9r4/nqMQqdZCMK
Oz/Cwi/CsDPlBdK8R16DOLI/Zl/oR3H/ZTucrE+5eforEUZUEjfbhOZ37T+lkw3HI7ZHh8hwnamg
td4EoYcqRifnBOnfKRD4kFQxM9RLtNow6hCPtrrH6LQv0+IlNIrqxXOEDTfY6H5gv6/Wk5cEsKCq
gGb7DQaGPTVpyLcI4bNX2BLNbGtYWDT0RjKkPekXK5WFCZbppzYfR7wBmKlbh5GYlTPoLy5x9KU+
YjHReKuRfvlnVUfO9zPbImKKGjqLnAvOMd/ulojPlwC1/FKb7ZXIgNrJx7FNVdtwYxV/2WAUMC9r
CXK4u77PPlbeuYvfJOURFqMP/yJhQu0GV95F2PAId4JLUT4jzLoIMsHC0/1zSK2uWkTrh3Tmaubs
SMPdf2RsfpCSwkFUx38bJ06Im5VRUF5yXKMZc7qUjXwqa/RYq0hZbxJkn6D2ul1Siaqi1YshRwNR
E4I5tSHN5h/wr99xFseTKdZjwMwzg8Pfz+PWhf/EdL1K+ghV2im647Rq/VGGXvCv3T+esLr3L6Cp
2+6ygTeW4muGnvRLlGp5ohjloq4Qs08QhBfCzfNZiUIef+EI/j2U6mxzXDpLdwSUOXta7JhaGGwG
xIl0n9rkaxzPrq1yCLzeFFUqmyNy3AVgL7bPKnwR44PqzvZNZAzJpsdd09sB1TCvdAjJrrjdUAW8
Jhx1T3bKKk/B0hyiaCqg4KBU0DEwEuWNlBoRMkcOVlNGtmzIwwDk7/kDhAt12+Yobv+QauVREuUW
jVIwpaMjKLh3nmLGBmKDWK7IV41OTWRUuvn9BJczkexd1wpvASwyx7qcs5zEc+UjDRYEtzE9XiNY
KC4gCq+TrJChay9HsiAKjayyuEEWb4QPBry+182drgWRRxlzDEsA9FC1Iiv25RsI9WesZbH8jE1j
deVvWwUSzUl77nKHH0ZD/Hqo+1xJVIVdA1MSgbDlwpMOdpnRpiP9y9q0ok/5K2mdCnOpULFYgFJP
tIBomEJ62MS2903L3EZLw1hJpMdk46OMcIamXOyGEIatXkN3lAzcASD4Qsl6uSBJkegVYvExRd2d
4RRJ8WgLQi34cQJO+yV78zIscl7Fpne0flulQls6SN/3KdA5IM9gTmLqBNKXYNulAWndFZORxasR
icR+gf5xzWxxrLR+BzQh26Mo2arcjKhdnyxcF4ozb/7pP0ZZGkeyAnz6X0RdQK2YriOdZxG0TNRF
oma/2f9JwykaFSRGqig44oluM6W/k8iQbMftjDKK5XHT+tJzVSHZg8e2Z7a8P9fcfPGtrdL8Xtls
Wd+DoIqXVwfvjm2BEFsHr5DSuDrJlaLD3rY6Vulz1/Ok2rL0s/WtIASVRCAxZPPTsGuph6t9h7cn
gMmdNF5e6iZ/4bHliHwmoi94qZdBMHgKNU9UNoX0eFpxuDvcSXLPwgo2y4kSOBTT5PI6H1TCORhy
vKSWnTn4BzwlhWQpsqWgaxZsom7H84gNx7Ri6XcqoeNwkcz2c4CHZhrniVYrUh7SlVRQ8BA5XpRU
/+YTZj1hkveLBHR97Pl2iTn85I1JQmPnnboXLSRvbnvX3BHYTMVhOd7tmFOKkiSV84N3IMpYjJCr
pUqj0ShiqIxN3WaTrMlryP7XBbI/vX5Ws6/gdVo7NGj2kiQgTKPK1fyRBrM/BhSX/eyF54MHnvI/
/fmXbA87Ko6WkgOcTXSPcaImiZXYRi3xOBYTAp5pD+1RGXLrGCTzp2WwoA+u+TF+H5h7+UVmNcaS
mCvIoUbimW/3eva44E4kmMMYu4/9ziwKnG0E2P8WyPjU/Ejfl/LdYPW6xGiPVWBJLZoUwcVE2oTD
USnEuEHT75WTrXaxzhNFv/rNTZ0NKgJ5U+yd+wDGp9MVnxaKneXF3xbQLrGMhTWnqf1jCYcQsi1r
2LCzWY+zK24SKXnz1lxvN7T51SrD4p8oEee/OoHvrYvT1vQxvA8So+ocE1wxGGaZGhud0EmNO8dD
z93nJF9C5lQurTNCdCHHLTJMowQztdRSGkfg/zXktXy0BqAuvwDLQ4hRCKwLk7tog4oBLx6BHA09
m/9aX7F/9YS4YV8VWhI7jzrihReO4QUemfh6oWxF7EWNMjIy1qIIyQfuayqzfjTq5DkHBf4C6J1E
8ETeYrNyY3NTcDbJwrgx7wQM49QybNcFX5w9dcqT6VwV280PbgUE3bUpD4c4TsZk682LbVrZWcuy
VOJKq18AeOWFBeKFapqxl4vQ5D+MNgYN5RY3id+rZm9ybKoV9/SNI4eGq+7alvimwijgbr2zhdov
MXmhmK4W97aYOh4h7GRksdSP1bXl1nTvgPiv0oXJXdDgp8Y9DsTYBa5Xd2fa2jKTa/ldy+VPstFY
1F7/oRMPR9SIT1Lil55N3WPn6CDyIXWys9js8aZomvdITprIFHhSpTuv4VuEVy+GdFxg3OWBwW7W
ken4wxSlr+v2b63Gg8zcEMWu2JCmJ9Pf0jHGcKiyXcw7c2toJVmQlI0m3s3xiNtaFmyn+dL6olfv
55ADowFRvl05cyL7lVPqRZz3Yx6cwDnXHmwW5/putPnqR3pE5S9CTL/29Z7QB/39iC5qK11ymqdb
9XgR7xvgoQ9CssNMJKSemlslyGRjAsNQMnqKzP2rG2VtQHV55+6y1sUW1bqTNOOnxt76Nx7bVGGv
WY9lY40DuQ/znGD4mAOjVB0UpE7dj5B1Bd/iKKG783K4hGSVsWXt9cwZSKf5GOFHe45S0td8wGOa
Lxr9wtNsxou688bnfscjVgwPF/Y4pG/+SmD3J9szSipw2djDZ/pMMbR0FsM7kjwANJab1ZUXxsr+
mn8D3fXZ+Nux5uf+j5zS8ZsZ1NA8SDGxaCdPxIZRoaOTfVwmHidRcCPFjINuUsOyu38XqHUjtayo
vhDUTVVJoUwKPxL8A2/lr8vBV/YKCEPH1GmkIR0w/JXBSLGww8cjDCS9wxouwDDyl/EFgcXqx+45
9gfouqsmietr8Wpu6/RBGlkTF9V1My+5h/7WDej3lUg3oeQU9EojfoTgGYZ4RuvuElhkQ3BpW3+v
rwfLEuDMGXwH4k1lewF9gk0tYxxZuVQW3Qwbp0RV960pAy59fIXXZO2kknUu0OPpQGUJpCLNTpPk
zaAhVM+vUQNyV7ku+JYou/rYnujEVG1X1A7fkGhPWijehM9GPn2VbTwY91Vl74qUDbEiF4iy6Tvd
j4C6mLrht91l6c8TH7K+9xMm1Aidh9kc8/WAi5NGyuKNiRGpQm1H/+kliyGOWSmorIn62t/ev2jG
oUmsdLzI/OHdStrAECAigwNmW4EnjsDAO8UtGZiMB9IcAXFLZbZUtsEI650VsOWrhNG7SVy0JeqF
47XyJ9Y3LitjyHO964yAMhd7BqYqMyOuONLPsAAVkLEDJ/0VqY002uiTl6dcCssenwCeTCiG3MSF
FXQV2P9ro6Biw8qx+4NDcFx0wMkbnqmzGJCwWFXz2kRFFs7co1mJV6e2azBpa7LKY0NCGaYoLiOa
0AcXLL0odw3bENfk58HjY7uXSk1YEcSUTT49jnpNlrANqTPX2h3pLNAvXcdrCige9s9BPI5pGl17
Em4s8p6OLJgX8H0yaaq1L5+GsNXF8q8HZTEonynPxOnC5D+NA6SsXhx3InjoJsfAcYwCIKKL8kbT
DxSr25ahRtteJ29GfNRgT/CiFZRRH5q854G1jP1gWD3J490NYV4hopMDoYcNCAuSPP6YZRzn3YpH
U6pYj2CSS7ngKLLey0qJg84y0gf0LmGVO9Xqe5LbnapTt7K8zgTaYjVLwaX00j9doEwf4odK5UgY
3b9rwK0XqyX2SaCz1unPQjmrRO+jsrZWxAs7eYgnl/94+wwWMgXJT78X5KITyY4hKUIEMCfvJ/i9
SODWfW2VSnKXY61Lw1BDXpi/Z8KMuhUt+AKCn49NPMVyVVGiRn3uWXyoOTLwfGYz55hWazQwkayn
YjGLYCr3CVRRkuInzRgWWFeldE+8r8Rh8AcIvx/g5rYKU9TA3LNqVVcQikqmiYO/1fUkaTdYpk7v
hY+jZNrtA00YsG5KLu5BZRrXn+n0RNaq//LUtsHFVc/KKzmbq/pS5adoEL41wJ2dL7ZCQDWylTkd
sLxSZBupLbfwMHQol4StGoSzeTQZ3CYW9UIaYwftYSRBXCJ0YVWzj0aIQDEqOQRtPRN2iafiA/n9
s4LoxXRdAyT5gFaP+2m+BEQ5IKaL02hibvecFCxNTYDrKpemY2HXqBSrOTgIFmkpYtMR/wtcaTtu
qCoFZtj4XRwgAtzMF8LySfd+zcLAghVd7HVnPLk2rh0HfMQNOnpGf3ppPCQuCKeXSlwGqSxiCrGP
B2WMsy4x48QFphGfhje5695pqhyHhInzTYzd/EhkVAEp48EYf3cb8XXNrWJGvg9HZ9K5EkDnIlh5
7vhB7vJzsT56FhHRLdqM3i94tjey81vkOvtTnSgjJpVahlcAutwSOiKKIdFcCLiHIKyxVK/E1b/e
xeXudUmDiCNTTvtwZoNZOBd9kKMHKeUtDKCBp692TdblWb4YtRE7cJWnf9ieSwaiD5c/2dlnbn04
dTwSyLHkdx4g/k8vX7+amn7xVYLDBo3GfaTr8DPMrvxIu0UfIMctib1y9eno+Sv13z7aa+oxdUR5
MRzYGVTv37tC2HxHQc7xbB/BpjQ+5Adb1TMmm5lNkkFN4gUJ9PPPrQkVSXWRvL0jR/4/SBq1GUP8
J2ZG+5cuCKOlIIjqLzhHpOc2dyoJRTANsdsoAn2tFt6fe3KutqLOkt8b6r6tx7Fa7Zb86w58eOpd
fg+RKLkAUQbMyK5R3WqIpHUlia7WRLkmMXioTGSQh3YRoRDTxNMTDMATp0JxXKMSZECxR1SGvF8a
J4s2u2awce0yYKueZkB6IQLxyCmskSt9KjqgKMpeq09Dwa02STmClRcsyzR1+7WRy0A3qKi3HIzp
e7TWMfHF1ptmBFe8XoEWq4jrFllR80aOKzDicPJ9DZt4Q+SX/oe3IWHUJgbMCNDKyXb0rP/3iB19
j3TT1U2/U6azOm5zCU/bWCceIC0XjnH6M2UsN9J/3v5ij3WQUwZQZ60Obr9/wXdir+YOVCuDS9B3
Lj5Z0hKSQ9NBHjjMGP/9HlMzdvnxrX+xEPe5rZaLpr36aSD7Kkfez391Ac8e0qKxxlRI3FbpK2T/
uID85wgRjh2Zj/uLxomxpHTjxSPDKSjzruWBr5Ch3rrjh2udy+PhkyuXQQmTc9zEdnL5zUXsoBIY
EdRerG9/viaOLx1xhmfzLS0DkatvjNNoJTKTtJfEW9DzCJGHI4yP3SiD7oI/OyIJt1Y9fD3/7Xd7
1yEdJPAseV50y2GpP5hqQIerhunui9OkQ8NtMWXjwZt+rOIgNw8wz91hBRmRcQnpzTAhfWjf2Ses
UUcDFhirDZRmt7tzu3yDKuF7dzb9PlcsbJn5aB53ncYuddt1QriCZnmNyDCjYpf2EVmy9fpVoFKp
x53JMKxeHkbkvljBndON2vVhn97yFSUawbyrrMEh8ODDF7deiY/3sePVnvF1vB1P7Ya21K447+jW
kFOzTBazkwUpMYjj9AZENWhIW7olkzNss7iax5pCvCXdaA8iXUO/V1lxsuE9eKv5jaZAmS/gIE8h
WpeMRFyYq9tSqihoEZqdRXKSBb5XnCsozJV9Ghg4NZrxFu8djjSvz2hXOVgISmL4HG51bGFFswqz
ALk0o+LMvpY74csjxmUq6rFbWfiTbIMS3SA2Q/jK92/YB7Z8O7ZQ++rxPO4sC9VQ3xRa7212jD4H
2hAvPmKdjfmskP+2+r4XSzz7CbPsVvjo3WdZw+WvJ3njSsMk8RJAdmwZca83HNiPVWtJcib5KO+5
038IF27mLGcsfmi84sBNj9zfX8g0w44HliBN/RnDnJzA9Gv86bln3JnPlsvRJvjmss40InB8yjs8
tHHPVS/jFZrgub/+5tFl9UHTR0PNI4175ECgA5A8RYZ15fFhoLngSRiohCBlYncXKX+NQroikiD6
zMCKIwDV6PhXnO21EB/A9E9R2qTwmmQXz2ApHwSp+xOTwLgrgToelzu4cZ38TZ7hkpPSgtE7Re7p
K1w9nAQ5IhwSnHH/+5Bn6DHqXyfnEzCOuJSwNfyPN+ZhxOYfVxLUTQ0dGXXEYxI4r68FwzcN2eLD
MqNjGLJU5dRgRbqubQEHwq4Sbpck7kraupgCWWkvN6dY2Bd0Qc0p/lDGPQyfgp4w+JWWLAXRO5oG
PD4edISzyL+2VwUmzy6zJ3OpAocHKU47fluOKncTrrGoY/BDTnFt2AcTenNdEp5iNxf/N2/TlFyu
DYOJlNSGWFO2ynyJrwKJOfgh/CJZKyKhe+fDwxy7Kjr7KYjJck13BcQjaxDIBc4u03sadWq/etww
2S1TBoc15VZFU+osccR2xdTy8I5ZhG4eny0pMtNL7muSZDbEJP5DPXr4avWameT9KgjHgMKZAiIj
LDa49rRtd+1FymqGzJhPuxDRWPySs9SXthMeCQT7z2mcRwY+YICcNqX8FYqixo73v1bKWWVM+n13
F3PCC4p7wr3BGbl/6daqtNhhg9KfYiTBuszGWeqCMLx2Bo1ZvjAAgZOUA6xfOySfHB7HWZTn/VH7
rHPUWY6fxgH96/rkLSYxXEQ0rcUnSMCThQ8V+rd0pqCiXpXWMWDRVXYaL/IyAegqC5L3oXcu21I7
HlZlxCEyWExir5WFMlxQ64L9lUs0dJ53ffIaQ28nJkCPFmLFqkiq4MdPbrZvw3gacPQQooffqK/s
K2eLeoHqE6kfsmYD9fEbrsxryAoTdZgFWkHGSDfO6Q9Ufb+JKR7ZB/Rbi/pFW1LoDCw0xsAer9G3
GgeGfF6ntZLUDwoT4jObjyMu7jK7sIh6B/7LB0DhEC1JWiH8zvMKOBuiAwHaAC6kmfW6bA5OZuLc
mfFa6e53cDakkgriD8IQ1gagG1Zlj4YrampTvDfxJUDUh7xZNINxvvSFlsDslJEOKCvIF0fqHCbS
Vx7OThfXNdGf2TjG1/0dJuKCb/E/4pXiM00PgELtsTdaX54ZObYu2FkUgbluGA07d+z90VJNW55g
Xn8l8Yw7Bc566V8SJVeWbFNyQEYb8G8gwdM7qP5e8iG5qEsSI9vrUR3ze3bP/QHoABZtF5HZSsL3
Fk0BjW3LzMC3gTCykc+i8vSQghAg221Pc4Pk7iachb3VNqVKPcSL9kGrVpVcuqHrwoSzvxPYR6GX
LCXdst0WMio/jVkLmbz1fU9Crd0KOUo8mSOAB5LNQz8+akaXBC2DuV8yZ06bk8yd2EOemN5gF9jl
WCZSCrVNu+KsXzf9t1K10K6B6ixk/QuHpAahXl7ar3sL0LsKms3F9qTgpO1Fv28/vj0lp8xETgNS
a4p4B5HWngWtnbdH/9w5SqB6dsiNoAR0ED9q9rsy5JlpK9HUwr11kWpnxyc/YLZThaqJMYb1P4ac
Ry/KwfF5RqeWNc5QE6zqOUrExlVyxYErXfGPuTxLm0eRk4owQAKxnx84ZL+dBVLB/EM1Dp2PNZYz
r5FZWQcPevc2ZefCKV6g6Gt4Fujxa7IaKScfdtQcFewi79T2+jmuhA7Kvoq7O8IkuIPzEHSpw8+W
bsTjM794u9GzDUEupWguLxTixel/6xcIDyZ8XkwuW9fhE4VUbrp+Vu/VaE6VK+WkGXNAnqwNFOWn
18VHkXBsL729vazaZugztdriAiN8szAR5tB+sHBzSO+iCtsP8nUINE5+KwnqyHMQpVOQUNyTpQd8
nnuDShb0pXG/aEonkHwCXJ9qiqEk6MJWA1EvOUyEEo39cZ7JOhYfCdeC8WAklaZHsxgBinqu+MF/
DFpXGoX5LlDxPyPNMSA1sI05VOHv3JGBOwneQI0A66gJSiK7sNe6H8uEuTqOTafCWfQyWwkpsBly
qOCLyHknn3g19O4WA0Cw65wXrUlnDgXAyYMWyLNtnLI8kJFnKdRFVdc4DsOfzbI6XiUD4q2fwd2i
wNIZKSaGCMeH5qURdx2fEevpflIHDK3rN5A5YbapZtjC6j2mtHSOpnhbPC8CwlIRoaaTNxIREvZh
RZwth5v6lSCHrAN33bYg2nAVt9q489TQi+TWEw5biOcdvMhv+LAlDE7ULharTA+Xk+j1uailVy+t
D5RDx+tBUXQsy+hN+G/PODo/1QZ/Y4gqxvdOvS1sOEiH/wKoEUeeSOAQipDkudoB6IvTiJr1bB12
mrLfYc061YNnsNiokfJu9kU8xhSk3H+hbGblf7tt5SbFOxCujzxdwZCbuCXa1u5gCQIPCnPVFqou
eGXUxQiufWvHjuVYQRcKtD6u2UWuQ2u1lDyN04oeMm1gcDRz5e9j3PBwtJQ2w76oZa7nQrD17l+m
5rnDwhcDJwA3gqVLxdJfAg455S+Sj2GAn1gE8LtTb97c6OTu97oBjFmoRI+wFwO0Dxbe3XtLjbmO
uRyuitF4Wtr8dKhWz//eQ/GkZy4gkgcUY26ilNzQqpmFuyeHmdhBTEiSdwCkSRFlAC6NMVijcUKK
/C5StR/u/uUYHhfUYGrOmnwP7wAcPKRrH+fzhFUFbE/fKhyjtekJ2ZL5cAGPQwmRtdEhxEUy63Dh
X1aB/e2EU36pwPAJXA976DCy/5C06q4naCrcxZ+q4gY52/V9BxH2QSdo9/On7zTGtK+kOJ+joqDU
p0q8fR778EpT4WdqCUEFLiuoxI9rqtrhKbY52D5hjv6g0FXuv/Vgr/3oZMjkQ5MvF1eAnV9O6LdT
mAfKzwQIY7pdDHv+mdMTzAhv6YBDGD/2sLtBJa1RXT8hWK23y/sJdYjM46atA004PhHF2bOMW4Te
7fISPR9g/IGU7m+LjJ2/AE5IWJDSLmJtHS2I3xJuE/L6pXrE39mPfvYVZmGYnRv3HghadoRAy3M+
SwWV23f1h9o5y0CFEaiylBvU60vBJ60j5vnqGR2zitZ3+ccpKtVWAPXFERXatE2ZwMvj2+ix76cG
Izl3oQ5UNB2H2gsrRrqxpqwo/zN7fRx3HVVGhSG98WR9yKBdu8PnCR/AiW/LTBRlREtzFsn6bHYJ
ElRV4uHHMMZHEAGx7o6S2poFtIee2UgBMangBdkvozwWGiGJ0GCNG1TG8n4h/ffuqfdotwelPXpL
g0BtVdiuXpgNZdTWPw+Vk1Ggjq6XUVI9ObFSNY0seovrH6DkdRpwBx2FEwP1gDpN5O+NqeO5sv6X
qvmLSTHyflImA/W4n8GuERkUauESfbxs+OdAiqxXE/mtcZ72+FAFTFtsXzqYOXQfk7TNwSWrk7mO
d6gq8z4Ii4JqBpqksQdodcUp4maay8lIgFMMVzwynjYG/75IotvBKBSW5XOeQpbKSdBNjdudNCIo
B6yeEqSLi/WZbphCyYRa7rgdcilr8fd+Z5mnIDH6c+iE/hQoMIIdRHc6LvfvG7f09leYg4/98T6Q
AT7o3hBtxwO72/5rFHBs1YpEE2EkrysjeMaW1aZDO6ayxjtWGhjfSIzErWS+t6SXsOWQ6mJ+2Eyt
98Cdh2nNw98/CZ9iFIB5WIEqBTj8caqhdJmt7PeOSyd7auc1HDg7dQPWZDfGolraIBsJfC3JW9mN
xboetPkdasWjJg3Kr8IITiy33T8xBm42E0FswGFI2i8LEyqZDt/RcK1d7prxuhlkXzZXn4znaaHA
itlHv9MmDqSlXR2njrgXJXONm8tfhD/FGVUvILVmb7RK/xZyzpK7xUj5YN9ugrgYDacJ+uCEHZ21
7SgoryIS1uHx3NylRFSzK1GIG/mAPYZ1PsC2iFVZVr3BA0SOZR53ie7/TFc2DqrVlyQYAy+ytl2U
0jLN9BXTVanmDzh36v3dZ9bv6jNYyCJE4McMM7zch810TA3T0TcvZZVEmapLgH5xWZw12oiD3Awx
ytTxFDPGg1viqzMxCYZTMw3Q3d7vlysac7xxHKcmY2az/CODdi8YWxQOsI6gr9JLlqBParAmO9Fm
nf4S6DzsFGebmOFM1PgyK794wlYuRB4s6+tGw83pEyTRydPs0E1cMz8dKzGb7nI2rgttllDWqO+c
yTheyno011QCEhB1YLU6rDdnsR7n5spCRX9g2O8FKox+LGbemzqWX/2gbPLh5Vi/v6JF4ggGGBr3
enpjbMXoN8fQ150iFFbbw/McSd+agyOTRUxdW2uzKCzg3aBMTfR+u8Mdk1BjrXxHAIE4H10AKTSb
NZzn73f/9rbcnK2kQ+QxlCb/RQNatb6tMPLH1f+an4SDEXzLO0q8AiNPA9ITJ4uzZOx5HZtSjuFI
P5kJKIZVqO4Q/C7vJVS8nlULppa+Jt6aBpqSxgJOYh9PHL3XWvTcYmFdSs0HjOO1pKrdiZ7z5QQ6
7PIJxsQgn6cFMi+SvRjJFR8TmZ1nrIZ3KAfI4ppzoKW/WFZ+VTraQilQseTyMgnfJbFfhxdzhhw4
V5ta0r4YiII+LtZ4Z9x2pbcTjHXo8WQJwdLgLinSL6ES3LHqzHjF9L6lMcw4YwsorKcyJTx8Gjqx
Ru1Ua4oDiGMAff4+AKrqB+Yh/QVXkrTwzpTHlevuMOikWpyUE3y9DWvYvRwCnj/mUSk981Gr8FV0
HkcUjdLYhvXpxX829+R5f12I174WWJWSGHIUwbEGMNfdGfENjyIbwJlppdfMItj+Zic1PD6y9GDy
vm1tZFFmIuwY6AzKorCQmdSe02XYZlK0q+aP2WO2u4bC3BBgIbsbD8v4fu2YirVEi7eCURc5XgPz
SxZmbJbvEsl6FZ4b7/54AW372l+6DHAYL7uYtVoX3fX3nEPNeEtfoTHX6JZaMeq8sBvt7zjg/Hzz
jdbuHJZP3rii+sAANKq2Q+XPNhsjPQDOHPNBDPkTOaeTc/23laMEUKwDr+QbnMQZdz408kDyGLOd
vAwOEJw/VfihAAWK30iDm8/826CPGzeGttf2Ek8FjXi2rVG8pDpTcNSAmcyw1QHhsd2GhvnC+4Vn
MiexgrQODwYBTlH4sDX1fI135WRArStnxb9LUYM/VqJ6tjljFUM3EofYPjm/N4Zw8UBMiZJVQbx+
YLZUhMhx7g/HzSUiIHwlgTwZPczkru1hDY8w+fQMy2v+OX0K3sTqIgLDWksqkHGvM1OdciQ7fEiO
GRlAIEq7JMMChAPwPHcTwALQNNukF9QU2RG4vViMRd57GDv2xiZ9tlbBsVpotPiO9rU0z9+uJIlo
uQGBpdrjAtXbfbqFm2epwl1oz4qHrrnsuDshMi4MxlVeZZtKLz43EcXV8JPzLUfex3KUqdltasnp
SRJ3Ixb2WMXZPQkLq3HOxnbFIsKflAGikTYI6pBf5xqcisBFAGSEEklt4YK6byF1L7GsuNFt4cgD
PVKS1/h6f9TrG9/BnSwMKBfAy096CE/nNcIVziieskJcoZw7npraDWlfOYN+h281UJNOQHiuMnPt
XPjLXmtmtZVCJYYmFaSS+PfeIH+sCzO9oUOG8cuJ+HBUfMcKbk9+qdovqukGNXQhHbzkSm+KI0ft
I4JXsynKk1xGI5OVZ74X8yozamwJNoP7aYOAH/pPaxt4FMl4c7vW9dEyMXYgUVeuLT76dbf+tsxn
VcLOFHs+b6FuoDQDFjv2uCcScQ2fCaaGbhFnQXndqMAgZYWcn7YUg92Y1VluzETDD1U2xKtYzV/1
wiJ3m7ESe/3zPHyah/ZhpoVUbklczsNm0MHtB4zsAlZBBkTpeV+RtEi/eBDm8248e5KgDSziBHjM
6d4ZP/mfEa2yxueBhi/zi0ynjP6EOCvhUZ/fj1WFvf4fSCi84Hk7bqmj+YV923+dVkxOQfEgzZKu
UT4k5oQpPXSeDNY8MZWDQF/qbo1EVjM7OOGse73L6IXISDw+lS6yNBeAwJR/sGMilnVutU8jVIg5
59GikDQi0Qg+PswUJIH11HMDIAe0JsGS8LPQuPuIjymTRk3NYvEHMLyyki2HTn2KKKLm6naA8iNb
ROdWW2xD9S56Wo195ItkIoR3LvrIzhvEb3RYkmLGdRbpw5sVorPgmgantjExNbwcLc1pFyHMx/5U
3POUPzBo2+kEAGoa/eYJXB2jxcTj3dSSCWvztrqsGbnvcMZRnbV8fWFybapcsvFQvdSRRvBzyXjP
hGAK5KoI8oPj44XuCsNP6vVz7UCJN5A+WkI51h4wWmPTMQoT9P1n0s4Xsmv4zrJNeeqrTiMII+uW
hk7ZJBh+U/adwT9p63FUFIARDKh9XqBJoXjCllX4s+jdes2gXfIzoJjT+uHXIbm/JuyknHLHU81i
HJG18SScIt6RgjUnYxB0j4XAmTMfN92Pc8S75AE67p7Zr1Y5omsmxELOvK2ZxB9t09O4K0s7Rghp
v1R9s+Qc/WfzR1FVmHRWm2NsAUg70YfkOxoRwNxgapFEv+w9umac/sdeqGUcs1e7VkiDQLR++O9a
8lLghjYfzNe7tCDaAZ0mZuUwZoIckH9m+L0XQpaR3HPXr04pGcROswRKa3+5R8HV7I27q1cYi+H5
ymB1CB+CvF83tAJ3PvrRcvU6teupeVpaU9FYnW28I7FTcvyKWyUqLNPuE9V0gzkUwBVwbCA+POR5
yfVw/4r6QVQILri5mRpHZvsQvDLgkyo+n/yMPpPe5221XcyZwZOkgfBcX1zxjyu1ejH0vJcJzelM
v2Xp/h7L8p+jbEkeGOc7B44AY1uB3jE3sV1r2mdulUF4d0IE2esJWom2I6Pi1dWyjF2cUECh520g
LcksM4+bWj9hopxXNYz8YkKICr5/V/Fb4S+CkD/VdH8EdjEgo/chlMj996+vpj0sx6/TR5kAkVgd
O7FYXSXE0llT2aUGdWqMxW/D07N0Ek0ADn2Xfw/YTKj3ggl7+aleiFmexE0Z1nQ4909zKTJ8rNsv
SOFGWamYO5W9i5go9w6ojVG0QeRJFpuJKeYyQfPMr1b4HH1z97TlL26CRJmwCoxivTErZx8f2kkI
5P6ZyXQOP25wBJKsjmJd/NJGyVv5RwnZoaGHjqpwl92WMlKG5hPLlkDJytaa5ZDIU3Xi5UWnY7iI
T7GhM9Y2DJMGI3btAoLt4FR5oz0pcBADoyvC7CUlmZNI58gV7CHGtniRHeBRY+pyek4wqQ169xIj
2l1p4aQscOX5FIMqlYTn5+opBeC8ri7Gvy2CpmhRj1a22ZwBoTVUMePr5tFfuun/2/JwUc3+WSoX
/gnlWdr1+XUgT5stLI/SVZiA+pf2kmDyGB4/sslVjvN/zJHqwBznmyBiPluzd5LhE7adrkguXAFG
HZmwHOsEsIYfbwq73yZa3sLMKCNzJTEN+1ty6FnkIW25CMFdVMF8MdtQMXIhbCTwD4yQ3i3LJkd1
fZD1hXK16j3Bq1rXRc1jTRyI0xVmR4KEfpPvOIe09wGPELvW+BbCJxX40MnVuOq/qExwBYXXwTyl
mdOPe5PqgNgUM98T8W3Qzer2luIk/f1PHCIcEJOfC76tQ1wmPKyqXpUh5pyIWKV2VPjxWmggz9/U
M42WGBCIkOO/bCTBBjaC3PVq7eNbtr2Uv0yFEIssKjhnH8LyVrD7m7vdBFa2pEQG65ccV+igO46D
R7QGxddCUOLXHsdFVugi/ZyJT0f4Bbj5J0vJ+iSz3/0FPsEcwB9/rusT5k0Jhrc2kluIsVb7hrRx
ywvVqK0ccUS9A9yg9kh458rmsv31xjxj1NTy8lmiHq6TLvpG0ls706nwCXRc4i0rlVW5xX5/4Riv
zlgdyJc8Mwv7AxAgboOp6soKxRvj/z95CUujX7OmJ3Wmp/+fWHbsSJr0ZLLGNAUQaqAekbFQK55l
LMMlkJSGT+RmUKKxF8vvFtt5SCgoqDCZWKQ4RumEf2B7ZehtEvLqBcvjU4KF7GctcW6LXq3Ger6j
+WveY+WAQBaeiWO50Ij3wGmTrADz5gNGZFKxkWKeKIfYVX9tpMxZqIb47GitVCj66Pqs16wzeniA
GSuQT4YtRHQ+y7jChf322MyaaQnsxp9GbdCkGzRuKZ0sFMlibrvxeOOIXJPvPW8ON918oUGxzJbD
QOVvT5AkaLlliJPkyMPQgRqFd3TNcOKDFRPeZ3wBDkM5Fj/DwyKxNjDarJM44llMtBI89JtGQVRo
K7+q1H0J56Gy1Is4XsN1271czl09t/4L2xzDn0k26H0LcpjtNn2XpGjVUVNpXQBFEz+brgW02Nui
CEaacHXMx3sAzVmSzYMUlKTGqY2a00niweYB8YPjdLhu8JwG1AxbDbEUrHJT8kWwXS5GjbRkP/Up
WjS+hI4I9/gLiMkxDkXv3kIvL0U6A2a/LsTaQqHhWT1xXetZNKCCCS6+mcgBsbywuQ0uo5oDCSW6
pd6sxDet5Od5lMdolO521OCXaJI8/qBWXZfy71MYOYVp+zKQD6UOva6W7l1/Amq6NfaqKVq6AdeT
R51223U+7faQCQPrbgZcSXUsQhMatBPx96/wj0OwWYhGmY2r5iLx0LtVa3YhjcRn+YNo2syJQBWU
w4NXgiQogLCkJzeBG1XM4AHItGGUgy5UH24mJs86YrrJn9nCSXmYEBdIlDKiBJEffyxzbvQ9Ox2f
UvIH+2DP/J025ynIpC678GyFB6nuw+FgyuTvXK6bxLjdFJFXR5NCd78tb0qgWgfegnNbPDeugQfS
FPngWPwqdHNHH6XqLKB4r83hpwjN1Sp3ZzRGwTrUs9dRRnCJSfbcUhdNTpGYu9/wbrXK+ZiRxpCb
ErSB2X7ZtRDQsv6rgZuygKpW5UD3DPA3NtsoWax85Pd0lqPIUyBOZQJXGVQwkCDY+gZRkWqkuYBz
T892e7Yjr7TrDkx48sLtheM7dgBsVatvgUb4DE7YT59xhq9/E2+IgJ0Z5SXF6yrfyMWUByErvip6
KD2KyCo1RNhG7JvwmezAnRhGacn1S7GblXaJ03oUzJ5YeIaYSlipBPZgq7Ew6SFuTF3cv11aiijG
5s0bVHJz6w5/lYI3ZJ0arcW067MHlkCJ0VrK5DJlvoTa4woSKuK8d4hOybkkraxi7NZ+aRU85DfM
OnXpLgVPHnsVdushF0ctnD/zs2IvZ4NBYz8PMW/jiPxTfXRAhR2XIUtF8NXBEfkedt4OQTzdVs/9
qzutvSvA2RhOfeokdSbq+VTS8+igmLE+m+IqUJP95HT/yBiZfC0O85sB0Nr6GgfmT6gOZsevF5we
H9EoeT5rrbaYS6i2Iq+eqDARDJQxBtlUyqadCt/bSwoYzlFz4ba5yyrnVv7hxzQfMrl/WTQlMoCa
heTEOavTmBlrgHhy7mrVG8bm8RwMSI4hoE4vKvb2rf/FOKoN1uzuqgrqEX5CcicVPWHSVlQ4j9Zc
OYlqmpQqy/wAor0cId0Q9wnN6RHLj4L04c9CGrmJrnGi9DwhlkT9zrzuwX0wQyM9GVBwqATQIjUw
Cvlglvbf/LHt2jBAWw/txgiZpVANjydmudJiroJ7wxFnlBpuvaGAV6BIyFzwTgJBVXWz0d9a24Ve
mwG2SgpeQfojkv670q1+H9XnFnHSQtXM38Dt+WDnUS02wf8gH0/rSf1F9qlisDri+MTNPGR2RLcJ
wq69Fys5QCsULRoq8QGPw35+b9gAWEqKnqtU+iA0uvKCcYkNcG/3LCeZgL5RueQ9Uhm6QhnkBIV5
kgqk3XWCBJT5oTbQrmI8ePwAzbzGvBowzCwAp/bUXTkL4GuLki8wUGttHL50R5vioJ8SwtfPJQrL
TptEydySemmpM3i9R1Bj/ArNQ6+O0HAkL6Q8r8iYK4rGqu7QKygkv/zVYCszG/81+nuvWZwxnmM5
tWVbYmr+4q5Xeja9/n2zb+LBQyNp1FyKTYO7CKzRtChhAZpKp7AhtVgHKKWc0LK9Zy20qD7Ohqhz
YxOMxGLJPUzASbjJfFK/zQzqprtKZEJsIBQdZSGXHrUNJHqeR1DqFO1iWQ6XSBoi74Mrnc2VnY+7
/JpqGlP6LMswwDuLbi5dRP39PEZWHa2F85xH33BtHFlotpWNQU12eH2adqO7GkzzLixjwlV5ptkv
hbPrbz8r0I+lQlJDEW59SC7HEVkDQqaCixBj0DsSf5d13/g9Rfg1nkDklkHmE8LE1UBPDHd/AdPI
gw83FtfWaihGEopdiGWbQKqEkQEZ8yPPMPmICwCUPgyJeqRKUCZ1ZMQvN42LCmmmcp2zupfLCg/w
S98kCpN7vEmQXam1cFjAfjwImIuKvVKFTgpskWFTag8hx1pJ/AKB2b6pprSlDM6A32CI3eZBzFOM
SNct2ATAIY+xITjyf1hVf50EPCDHDv6/SOSU3htojhubcZvXxhsbYlQ/M5AE3Z/PuiWHFt1mhh1m
wYu+Nm2AvlACpRqiLV9g6TUCienet9Fp6cGsorp8iZNIvU+X4JhjSRKmwApQ/IENtPBUedHN8ijK
S+kQdodqDDC9VA0zbcYgMUdY9cw5+p51uKH/Ol7X/eMcqANiLjmBZAmBh8p7TrsGbSHjUqabuzND
Q4faYwhSvKxTwOvXTbAX42ltNWTU/pGy0OzzOs1nSmYfvBWxkwHagofmnTSIL9VednEdyQG1p0IG
TPNUL7Vlg/+BH6yWztuVOy250FtA6bSoTnFntPHn6XLjn3vIxxNeHHsxU/L4ZfofEFBnnHjI9+K7
6yYdlyERCxLk+E6wHzT+ev+IfWnFnZzu+wZGwuUrKyN8c94wJ28muh9AhOHc35h/Pn7ym/TgWi0A
hxnNLcMxlsaFqvtNFZpiSzD7RPutFgpvI7YZzd9zvfGc56mLWwzhgGGEDuqDMVlD7zunRnehLIW9
9QTEWQKa2POOAj7TK3Xvh8tsRTsx6L307SSTu7Y1zYoS3wgf65GM49l2ffzX+n1vvgQmnhRaSSTO
44i/azAHTJfzfoSIe4ojtnjjmkzHmJzYBaJQBSS/ZqxON8gIOV20HHUatN2C+sYS7lWGR6JgWU05
rYMwuBi8bvFyg2f2EHyXMGQtWHMhYxMdVVH/+t6qOIhsci1LwV0njAlxFhluEOQrSztyIIzfiIo2
SyuRrKpRp5qPD3XrRI+5pFvjhN7XuWUltIlp83XSWkjylY2k1LhkL6uEnoN8P40P8YDpST/mTN3/
XNoWEovu4jDwuWOmLv0CwAW039CibPo2y+zAu4yjAIsL2MonoafTTqvumj6bof2wK2Zbd2WeETgU
uqrvR94S86ieopqWn9aQ96akgHxCOi9sv1FC89L6JDZa2IumgLoIgoBriNCWfftTMzchOXvR8BBn
FBFgI4FSGfCWnlhIfZtiirgNEJz4np26GvWSYo+BZBKLSGtnaJNLNEUhN4REsLSU+mw4Hnx83swi
enrD7KAuyHbQE+e45VUWcQZ3/KGbuMiV+Po61pKcw/uwNVMkjn1SYEj8IrMrnyE4lDQ1TGbvp+If
HDZbhFJ7ElgpokfzVHxfY4IPNi8VNnpRqMu6z+qB6QKFWmauhUKY0HjiATwSti01lg13gWzQwAwb
Dp7uTJMo4GUw8fSspLdTZNlLgff8GZTFcZZu/QBoMNEewN71Ka365zG7ASEkd5wCUJIY57qqImu4
FQz3YyrVskPFUwiR5lQqpkHxDE/ATTspvq/z3oMuX0jROU13MBGF0U2L3tiQLmrNR4fjY+7tZpGN
JlqQv2Z3MuY3TwD/tht2rm/zaQrLwlNVB9ccLsGxeUlZ+ytEaO3sNtcNvsf6HlvBGty6b2d2+4Hy
uhPoiD4X8W08Prac/1pQoa/nnYElN86ERahjTdPK64LrzAah1suXN10QQ10R+KGfkRONNnELqaaA
lwy1MmeTED+W0+7yYhWtU1MfFSJvwqKUpbVQgQC7juocd8DRM1FQRXtXETgRBOOF5st86arqBxt7
UlaLQrxg++Cbr7MkSWtfuZ37DjgEh4fadzt95QHsumxGmxI0AH2RikPBjDoYXuyjOUhEandGKdnu
kssiPGPpks/LrNv9y0ng2q8Dokp8QhKlogFy3L9ud5nw3/Io65SUKbrTH9hEYed09pdpmDcU2Wvk
8ivapUsysrqfppW8mfdOyKWCwLQvxf5ukdSLJgvbSwB45d8rG5rZg8ylfwIdbq7N9ubXqibjYWwb
5g+tiOeV3mk1jRhYW/8swTb2op+oLJqOne5E1pQQWl8hJjdzToS9idH4BVOipuVnuHes8646iple
M72xnVGA+BiYg869nAAP5AGjIUfIausl4QZ44NxIH3OTBbdMfUvSQuWVV4Ny9WtKuKTS3CKjuGMU
CoaRywTKubDU4nMg9Jn4l4B1WWV0jDvfrJ2he8q00PuDLvXP9fxtHyEAOU9eU7YACljpdaVugpXZ
adjurdmDDZ5RmCyWVkbyvmz4ARKk6moS0qPTXZZEkC2evhVBFAgNYGNRTHnrtcw1aiPbv+fE4dOb
LDicqQJCoTvF6aqNpp0njiuFj2OHdnVi3cjYp67O6UrWxStZCpwtQYpqB4Q+KkIbeE0MAP11r+cm
WNOWLdf0QHRWz+/mTzURWjbAK61uoiMhIfbFV8QAur6nUDPfV7MCH1ppyA9VcZO3cRsOSrJqjQrt
xEgFtAJHnHe+HOozLJelNOEhHVZSs8R0Q/LtJWIeBszt6MNQP7vyQYyZ7t/GWQGEA79O6eH+YrsZ
EzPcHvKP6mmwAdhcS4phHWCZa+uPxhQ02TTaQ4qurmKrdQ8x3p8UoTwiVco93EMcxu8PrqrDB1Wz
8RStWL9NplVMlhWYD9RjZiavVbR/Mej0lBmG1pBWvkpp+ldFM2KAlLvHsWfzK/hhkFMtblHTVtO8
pRinXWHCeBQcu2TCIkRU9nSzQ0m4kmTsdgUOfhRcrhtZJ1N0Po+KpGcuSeE7G/7yk9lBbDXUxm+b
5IMTsHw5MCB1RQd5rMT7DaSf6Lx9R6uffzjyKZw8KE1zjFAc5+SurZyn5LO7rfN0tPALgRYheRLa
fg5lxRxenov4ZBu/1FtlSq+lRRWd1q9hOTy2unREvqBBiVFvioZ1NXj8//r1DkcP4hCxF8h73Dq3
vecaryh3jXPiLXNVp8X3hdyyXY8NV13ydtFnGawGn4QtaXgEkj/0LNFaTttxLrhagvs7nXRxC8jE
1PIqhv6c/px2k4rxry/mqIA5fUkjEL38+N9m0WdDMyxEKWznT1AaL7uoP9zx4CYiy4EHa9CffcdU
jRWeDyiueQp7c25ufDFQjVG2fh9tc8/Moomx9Tapt3a92beIEknU+a1ut5Sb0JOifw6VU5O83xVY
6KEGhyasP7JBtDvyAl/rRzPybuvbD12LU6KPzTY8Xp+I1DoPImhHgZVcfBcpWTCVfvWpi5q5kN2k
6kPd1a9+WKfQjhOPzJtpdmDDIvPkVqQtCOG/TnSaqQv0p7Jj4Y/clbVzPJ4dFm/zv+o0ENWTWLJa
KArs340AWPuUBZ/zSkg66GCYrKXnlv4fsbUImWwlvMGuMyXh8X2iwenD0BkhBbtrYoeaEXZ2BsG8
9GN+BzmYS76KrVcZE+uVdgjka2TV5tv2n0N496Vy6F4wPyGX5JwaXfjcERXUuwBlzevjtwRjQ6t4
H3An1pTLbBVQejCMQdYmaPN1OwlcLMXcPB9jfHlFMdbt7ly5KOD0zzWYvZqhgU+RkHkEzYkb9Dyc
NJfohd+wuLGeOgfL33tNhG+ImGwYMMJDEYvepCV/uX6Y/SkPnQ/FVwY1/zhPLGim3wipNUbEarln
qS8B2/8XQSKpkGU869SUZIOlflYEdjuV9pcU3RTmj8OEUzhhQpK6hmWaAn3rE3IBsujB4JdV/QCW
FUFtKxXXkLuI9QuyLaDFe82HkKhd81FYGrDEfofrRY3HuXAl7s8myDlgvJ2mfImXz7vNfxeI6QR+
qwUdDel0gpyF8NUzXPvpakX4FR3jPMKvfnq/y50lOBhmmCrjcc9DwCnEojVqvMaQMQCRLVKOdZLc
hB9IYMuXyMCC4wAP+O1NlJm40IF2Q/eFAH4ISSFeYKiymJ9bXTqyYYuxYHotcg1V904MRBSqfonc
wUoBhr3SD3a+sA7NqHjnO22ERLvuPEbXv76uwZwfFWKw3+UeYE3Bj1JdfYb4TJ/Ci08zcab7qN3f
S1kRMMu1vPi8FJ/2rdTAUcm3iayqeVWxqP707T0siq7a8L48Efph+eWAwC9jalslO7Xc9y0yUdlS
DJB7m1As2QlwDgBIj3t8+TOSVRwtFsn/iTvIWqw6UlOcjWW5IKaqqMCiw8k/v4+INeoOMXS381S5
sbzeZNaimt/zQhaGi56v4pHff/CV4DE19gh07wJco4EI+gUWjZQpxKdVKzbhsO6h131JE/3uqeZn
Qza7Y1y9//6w0LAcn7SQmGCq7IHq5xAAqJfTeBvVea62ZLuDTIKApZmlAy5hMNf3J4H/mVUiDzx7
PrZL6DzxRsVxdSgRk6mxrSX1FcGTf/dV4h6kb1i2lDZjlF2POE95KwAGzhtzJbHEMukgh1xX1vmS
5iQqc9mSgi/eJN4w8ag+SOO8v6oRLoJ7+r5cOSfdDOS/QLRAcS4uLf4HeHtU3aMKmaQnq0Hf5auh
FJVSFGAOwbR6o7TVMiEysd6CCcRMllj/PMk9NvWagmi9BcfdcHMg7P+RpK1J9BIsCBPTCnhb13iB
IzaISlhK1sLO0UtUCVzGAd9hqQiSiNWRdUfaIKFuSid37BpqtlQYlhqCI+bvvfi/Yas5x8H+U9wq
x5e4Nk1qy6IvICfasV4Uh2rr8fmR6aDxSBQ5R9Y3A8d3exWFzk1tKQRA4LWLQmxA6h5by/tMfe2F
1MtrSvvljcomHvPKzXJp99S1woduX2+0N/wOQwlx8K33KQeRyiX3ybBaWZk1M+HckN8RuxQ2oxH0
nAWe+mPgH71p/lKxzNTUplC/6q6V6pi5SqkyTsV9NY11WX/odnghUUJAm8iRcJAVUphhf81zRTF2
lek7QGRgFF4PpER5NF8kPM8K09zvyWdmP4s/sDN6ocYhWHfwuytAvOau9BY4r/4NhV435j6yd388
824cAn2ui4xVZk3MKNVQpYKLGLOn6uMxKE9L1tmsKvXKdpDnOUoG+yvMfQdmN7TY3n6wGxPH788K
qPv8P15cu2IKcDfndZ6DLXZrrpzmCgIK2Ezj2+rW1QbzTX/VynO64CRUipVcd4v6fwsMbW+yaaXS
jIFKk2OlGOoXDKV/dZwOZczEmHJLmyu34g5by0jF7Q378s6/6eRG2qIsB8HOfXRjGO/ThP70QiQI
BHgol+ajsndLBTov7tnbjDabRmpuMi0u48Tv5bUrkeapM33zj19eFhZZvNAIVhN6Aijl0QVPyGrE
ghDy6WCvSvgUy/myLVZD/TbfNdMQoMcN2tdUGEsCwSi0uZgqTXQ0iSBccMJupIBx9NgFojVj3gt2
NC1r/EILi96KCNFORWEOISQPioUkQ+7l6BVM5oyzzWSrDV47CU1aAEpGsRTohZiHTzDuvNXRkwNH
qthVH/XJ8yZCF59/IrCWD1gIxjfVp3knQQCBPEz3wWel0rxeK+FFwgodnr2YIR4NvL7R2hoF5XJh
A2yWGXILsYe1nB3LDfuk8W9/j2S8OMqqBeIfMq4ZbPmtmNhW5eZqnQUzLKTgnGGJmusoAKruoB8R
utb/s7ek5kW9L0zhyOTp0iMXzDC9ySPBtdIZSRCIOHoYsZTF79wLwrUTIyksA0QxCM1ZqSFGIKci
nE4JOX+NGyk9znmgo32uOZ1Cl80ZHFul8oY7TIF46g7312i8sMsH9Z0w2ZNlu4FI/WqG6vZ7YTvk
ssXlIB+Ley8JUocCIUv8tYSucV4k465tfyIgHNVIF1hCuz1JsG57ZoANxuGGaMoWsMYO3eBh0Cmq
qGqBfW7DZ4LNzEGSXoNYoZ6lNPvdEd0xsG2hEyYnuII6rMQXUd1GmvYNwJYGcx0/IR+E4Ur+jxYt
3z+w+eEBe1lMvJ18GK60Xx2vNVdjxwup7usERE4qx2pnrMNs+fDFJxcCWYzwxkFfbeBtqWTkGdta
okf0egi51xCZIZPBw/UQIG0hv0ZV3Y84QfhbxtBeoAcMwiqR19FPU+yEOs78j/muBrAfDyfxG9Xz
a43csnzFAAILWw+kb1aTx8y84GXaC4+GH33vc4J93AysutZNrfei6M0RtMQYekcp/OPWubXKGvQQ
T8EPfURLpkjjuK3SJ2Gs926dioLZP6Xh0TfttoPRiVkRBJQkDcdMQZB6APGZaFmls39wwa+G47EA
FbSiIvA1U7TwcwoUnviqkFqXc8XyejDJBamGHZtFOoVz/k/Ql+wBz4CptVN/ZZLNL08D0RmTDTO4
9vttWPbDKSO8MG0HWrOpeFRykQ9w6V1Kadec2OUArLiVP8QsA3bNgYKq+sYmO+Hu+awbkU9ga6HP
qXp7COtzsc9ijqPfSp6YM7/INmXkOQUFT5cx7NX+gnAr58CKTWPfFCRBmLxwh8lA9ZEL0cVocfGr
FdN4g4ei401WsSR5/15xLdZh79LI0UcQwdrwVSqlCNSHI1V5YeQYrSypRImsa5s2KCD6P2YK7/sI
ZhF1kLrtDQxO0p//wKJlmiOaduJZXAjYDNPPHfZq1L8qadrGEiFT+LkgI44KDFaSsv3rCXB4kbcN
SE3RfXFi18hDPuOm8Sr/R6rGnVr7LYMADwTL7F5KZIEi7ZcQ9v1dbHj3fQhhmAd3ipnQrZFpVqbv
FgqUXx4ueoQYqEg67Tp4Clydk8PbxEBoYOtM3pRcjPxtSQCInLDk1XcR/v4cw2y53dGOkxadSLnF
tLoK0MRfDZgIpr+eZFMY/yKygr7fSOAjHFkaiuAgmwA/8Q1LnBFhkJIjK1e4Sx7w8fSQg3dMCxir
t/d5ZC0QH3+1MrrSwsCBSKuNIftwbUx6bRPCzBKHncSbBr8/jAUTvK9KC1CNzp0jMt/yfBOHXcGa
FBPpP7ykJtvYrGtSSOObaOLw+pCkVLfK+31fBt/uJvfbtp+DHc9yfhfFkcNNazx7t+5Dbm4+MQ1z
G3xoFJcdH+kINzvXtKwv3KqYL+StKSdyLahvhf9KHlKFHmlyNCRkE8RCcVwE9DJCezSCVQBVF2/k
NVIb8WkINPpVIfYD8vLup0UuEYHGKDOVzZdS1hJGHJfL6TaT9KR+BXD5vg35WwucAlw0Ubws2ZxS
Mqb8cLefvyGwKq3IjiaLKnTyugaXJrDMejmiRgLwirwzrL9iGIrPZK4WAjVtNKh0DsVY5dzVvFkb
tRzyJUSgZaG/UHbX68wG1g9RhFUWgCJbLxiphAkIwAqzkBv3ayv8LaYcl/KACw6hu3xx1hRGImQT
fQEgRG1oEreqAl/3tQF6njGxmt4xylR6Tm8hpqQ5f3Rv2VodTDfVmIk5SGt/yIwZoR2PLl7zTpwX
oBHnSYFfwKliBdx23GAdN7g86SIBfN6qLBpSBRyzDNh4+fgBm6NWYM46KWH6xqcm1mP5WM9/5ziU
TYTn7DdzJ1fbBldQsCqVg0d7a09mp+tHYVqUSrDajnxEWCY1OdVCcesbZVCr0i79UC8go/n/C8uv
kB9yllqyt6ko5BNQ0X7VAUjeZNtI39lnRZUm3B9h7NUDnwaFK4PIexZNCe09ASVbFXXQgrHIeed8
1juAqE1L3jgQp5Xv6+3UO7j99ZNdrfcefTsygkD3hIccfhscay4JK1L7+kYDHuUa3L5FPOHdskNo
xL1x8rXA+/Fd4pS4AWQKIJrUnrpsNCnI8aVCsAssh3lMbeWEpSgxBd+KXRKmFKvTvfSCc64hKz0p
D1RnhULhGfhPBqAJQEpcAAKzCoEvyB8fry9opONqW1h/QFJnMksBFxpZ2j7nN79I7d9msdrX4blO
KJ2ZOU881DHY7Gy5YBy+KW6UZ/SlLPjboPZD0LiOC4FEMrQmBcbben1If0680xbYadjEWSiUXTNL
quslak7oXtADMViipijMH2Zg9QoDf7tQ3D4iAqO8PHptF9ZyFuKeUlgI1QelE3wcBY3puvdVrvx9
YxwT3dLDMuOVaoG14gtZrd7MOcO8kYWwCBqYokYB2Q3uY3i02SJij/dRBaa+KOiLEQBFhLARo2Rw
0D3hMN6H4et00nZsHaSb2rij9S88jwqVjcnLzvmADau61+xQTKY4B86LZ+EPeJKaP0zLL6PiepSp
cd5esjmoqxaywSHFedkOKlOSmIm7EsqPCuJAfN61Ss477JWp+vM9ceBpUdwC8Ay7U4VJEoe106sW
gCfGEdk2x9AjN6PVoGBN2cLNmOb6q5cAtaCps0++LnLs1zDVq2SR8D0VuAvWbVznrbZHu+eX3OAq
kEs3hgZFTmv30GG9sSvSmngV5NzYlon40ob/K+EOtv4CLhKv8gzlNt85m1jSLKuVLDd81EuHnJFb
77XIlc1r7ig2gafqavuM8AJNFiAgS3ePVT8awrJsvY4vdQq0cN43Xu49IRpwEknEkG5t648Iv2Pz
mwlqkcgos8bZZBg3xjkA/XBgpan3vzFwrw/VCVms/yC8SbY31xXMo2849KPdgCvU+/4QMGmwgn88
yYQAzGDYOaB8I8x1vNh8RkmCC7SCJjAHJJJZPepONK5XQ6YgJXC5X37IHiUQY36FMUUEoPGQc3Zh
jtJaUq6mHGLlk7HILPZ2uemMkNsfZoMBdBVxDLYoBukhQGPgy1wTuaxOm+qd1zGgzG0eoIHhUOw6
GVauD7kjiE7bI9nqPfSKvxaUgGaB/B2UCclnFhb19sg+F+sJVGqKQh2hzSUFYWwd6TQSKJ8g1mxe
StTSD4cGNTkLs1qO525udCpNqZEZ5SogBUaxv8v9A3Rd+a8h850FA6feMr5RCOxXx/MFE9Q1azvr
Pv9l0i5dcAq8WoTu9gLmLgi+V3gZDptRjGH1BXEpaVu4ak4GRhCCye7tMdpYJewLZftBNbKgMuNI
Hm7iKu2vgwPUz4xHQDGRlYhc/tzXdHgLeJkEJ2SOUERSUbPppfXCyzI09VvBXr+4M5pbM9ursYoV
l/vmnoHHd5qV3fdJpW2lalIqb31tOd7SFDRC5lD5GOxTH7qhQ2zLY7KL+162hsarf5qakZ3rS+Op
f4blcfyNMiYbpBGvz0ZA5XC/GoIoUVTgp+IjwfE8E+zIQFnbE6ZrcunoV46vx/OMKuxv9sH7dUaX
JXlSNbum03QOex3Bom9G3Ns6hc3JubEfNtoFhwDfqIm/G5OH6qN+y4RxqyXrrOxKmTBabvvoxOF/
TrPPj03nu3paHX2rOkq1/V7sphcPlD8IZPuEJd0jW6jyOPO0+VkhTNCeG1f42yRgoytASuycZo4g
Ivx+R10UXj1xGXWTBE2+sRFjvIQb7LLHGzbFFP4S1fgejyVltstajisHjPvpo6uTxBEdXtLBdt6Q
ECgGbWxgWDc4laPSjosSw/xAqeSUY31VZ/MdypD8Z/uNoWf8oIo8f8PRRRDE1B/UcHJ3gy4WN5f3
0pCYdKEABq2+Zg0HUp8gLw+i6Qa1UZy9onwsmljyVrmJ6ZDw5Tyg9JaGf89hg89+Nd/FJSq5oixR
e+uN7l0VF9ie6mhqKT6gBnY5f7BOlCwuHJ6f5M1ke4DM2RSx1nwz2WjwRXrgTSfySAn9kNZvQXQK
pUfmR8U4qxrATjH3+rnjj1XmOxZyWhEg6w5mR0tiYDwLeY3UCLI9lTDK3YOUAfuAdu9OTUyn/eq3
Q042hl6d5LrBV6clbUs6jssO2pfeMfKZ1KaqsZixBsyZuWTPXVHq3osw7PPvR1+uPaFz/IIlb0iM
KcbrFq/b+oVAXv2OdLyzaHtEf1yvEsi/MBQs8OHbOMf9HNvQnECdK2B2UbsTzKwAQNGT8Oq2LGPf
5CyZbWPBY/ZwTJF8Mpvq5NJYAh0URmfyN2n4LERQKu+12E6+WqqZzk+x0sYUy+J7GRnF+LdiExp0
NEW3/yDjGfjoHRXoelRD90BgmLOnKu43PSzyPSIB8OZRw/LacMqtosqJjt/OIWNhyBooiAPymSQk
uLvyX4MGTOV0j5s6X+HCW63cOPfvQs9fikZeHMexADdSRPCTfTXdDwdoT06F2Cv4TCB3gyYspBUY
PnXfv77uHDmG5s3WFqkGPH2JZ9HJxqJwRTKoH3wz2oKYv84OqbpWkhJ/1qNHb2HOJ0nQMI5jin+u
4/jijMZgsFizLvHRT9C9P+p1/MOaXt88RZWjkPZlJBSAL3u/jR9hHHhjyRzZSk4YH6FoGZx7Rlqq
IpNsrD5sGHoDgoAub/bAvJC6yolBzp+15HGalp8AQQrNWCfyye5czaJJxPkyyi7v2m1bveLzOH5+
ortyxjvxl0yxd44ClKMJFpF4y0lC3gT4fJkTyshZb96CGGP2Lb2hCK8OEmwIyKMjUAPkK1jzD+G1
7wT12KMe6UNeFqV0KMu1qZ7QDGieV9CupLgUhB1F4XSgGWPADqnbZTviTXBWkCJECIo9WvhoB2Kl
Ihnp0beHh1+Or3hVEjPIgR2tT7LXi6SmYwco1eOVb6QyWbol/CxARmNhFlVLZ+h/sgQfCegpHUoa
qGUHMU+8yNEUcoAqUS1/5M0YS/s9fZMCf8tujvwLV+q1vy8BVlOgRm+FAQIzx0rW9XHLtplhjKMB
xQ0Ia63xO5PjEjM3H+yNc3BkMl8vKvyfMf4Fg9N/jbmC+gI/LQ5HgZt0WeNwfHxu/tHuLEBaa9cE
RPA0jCqwDqL1sOWNGUGXq7xfKokSOZutPRHvlUjfrlcs85ErSVdXcmF6aTX+kqIA2CmMIkBLlpP/
n7piMik0J0XSXRKgbLDK1eq1nG0F/MDf61jSw1JexW6SnxdAPuWPtJXACErQtuQmTh1G8hM5ZwnB
YKomyhxiuM6rm7HbTjQKhCUcx6HrJvkqd5ROsS6zzUqXDUw9MAsOF3b7uegplBYnNoc4Gnc/6eHv
9B+5vJjYDv5UHCCEc7ks3n45x0aVly7SC7nS8se3ASTVk+wdzp9sBRSSd2lxBQxrfC3mZggQrYK3
CmdzcwcYWKTPCf/h5UrQ2kTcJTkcZu/kjP7Jn0FuL0TZOlvLgD2SbjLJkteKxJ7Ln2ioG0q77OAQ
QpRb8MOxV6ua8sZ+fEUnaiGKvdaEEEFuOrtNaaDbvt6KLaIBut+fcYAAzB4JWFa/I05r90YVzFxT
M93DUzxo4X0v7LAdT6/51SVPtDfXza41RTENpnRxZHBGW5FtMOIFLRD87PYZfmRDZePcy1sAF5+w
G0/93uCC+xF4feLS4TF+ncHFpmXMNcXo/cVVNvbt6YmjAaLahVxxONEJUGeuNUx1m8rtai9rUNup
VXWa2E40x3AE91WH4wheiCbBE3IfYDOeklB8ve+aJ8xSkpiktSDCPIYVQ/X1j1QPO97brcT5fXa2
HjAERHU6KTCdaKpnhys6IVr0wN273V8QotOoP/lylpr75zE/ITheAfduxUYeal5tiYeR4tmaMt9q
YvhfQshWIP65mhMruVXln4s9afAgEAeA8MqhSxdQYyJYTfbApQa2WohsvTMzEUvfbZE4grFaxgK9
lEizSjsIu7qj9PfMPybiE53I/tZD/eEc+7ZTwXB0Ai4FKZiVq2AJTkN5uAm2dy4VneBbJUmmLGQg
C4rf+l2Hv/6DWUKRwcXvlnMPawaA+WcsMwyPKx3lI0L7U8MD531ufhSQQVJaR88Av1QQZ6oP6SCS
X8Gm9qcBNCVsJrKbZzfHSz/2LDlyd1MJs2I3VLu22ZLuVfqCKMPXWOb/SMSeoUsD9Or8Uo6okLUc
qmPuyNwIydDTCLphtS95K0FzYVe9vmg4paXJHUipd8caR7kOtfs7vgoPlp0YOznOMDoBkUQ6/iji
GAobB9HlDSQGqOYSKRQzw5ygcp2Jh/oLtnuLuPsyQgs2XwBiq28POsTQCYbpiEZkHMs75QQ69Sbm
OHuAq+n3UonezXycS3VRnNDK/dv9EV//VnLQzXyTyNB9B/h84dTY1nJwrz4QJtQU0o2IHRs6xi52
njhEGrFufsnqPHWDRPNdxlgRnhNpuutJDkIf2iYJQbcHq0XC/mbXXxNcfybh3SPO4dgWtibER/G2
AgT7aP8v6MyH46QQY+4FbcZndadkxHolGr4aHrsxP7vwhgg9IiXPPEctxHooRG/YkhH77Bcqrx7H
9lPGlti6Pn/pULaBcmsT3ZKSBm6A9pxbtOCIn8x9RAoi8AuZ7WyIBMV/SCj04zd9x42JYt5xlYhG
BvwgPYLXDxxpmVL6tY0UqZOPWHPUO/NfdQnddqZX1CMG+TAAfp5EIBKIIrXBEku5r/8mN2GAQMH4
DgR+vMx6U5HpGg1I+w23HCLSenUP42OD3QSWLMq2ms0aimL8T98eKCQVUQPySafFfCk6xnh00Y+E
K4zrBk+kkQ8ZscdAPTNRq0rAIbw3HhtAu6XQF3wEvlAovi7Xe3Z0y3VfZPiq4rHiyfaFsnuu+w9E
33cDxNj1wM8OKjunv+Ot3scTATWpUlvuHRlDVyVtNZE6cR96mDk3VvzkZ0UYIS/9nwX6Gaci50+4
jMnlxXs/u8MuExAlllDQaKtXqMcbu7jFoAXEbOYR/gSH7TH9avtEX4iRyZXjtQii0U0A9nSuLQUP
XqC2JGJgjWFTqUZOHLLixIgBXf2fq4t7+sMGcJsNd3hJG+Hy6RA9GYYAkVXxl+ROgw6H2eRB/tfD
fc7vrfrIMRfeAIoZbLuDUQcGqlIYokfTggYNTq3pVOtFnbgF48QTSzq+NruQeqO36y6WYfE3CBIK
TwP/uYT6cHWXsTYCcwDATfWVhaWqvAR3vy4r36+2gzE4VnjJwY5+05/o3xPNHiNNuU7LAC2CZN7W
OBPjy5kTqR7l05Oy8gFS6jfipZdfaVVFvAw/a+88mxNLJJVmhzoAdzMzDyIkUbC4HBpx1qm0xnfV
xvjehMXDQ1EO0aDaa6i7qRHA4LAy5A+/J1649JovZDur6AKnLeQ/74cMrJwW5PNVjQyZ8dBCwa/z
bFhL7Mdq0S3mM193FRNorMkJlxvi6+QxAwtsECrHanRSmvX48S6223WleuMgNqTtmnLY+pgOlv1Y
AEHiUUtdFNtVEIJclhwH+iFNcF3nKWT5FrzqVuczacmOIWMCkT5WYbQ3oFtvRJwEIczIcdefY4JP
LMMHZTV9Tz5ZNu0JniyTqtHgo081Cubu3inC2PGJ9Pcstj4MT/g5gkcO/GJSoaH907NJi40yufpp
WESOSBukS2GbRb998eo+gMTmgvCAXbF6CY6BIiI2p92Q+yC7fUGJ8a2wdcvqyKxMI/P3VXKVHmPH
W4GIizNMr4T/lmF2KhEWysPQJJ/pfRZMR5MEGn3oOe/jzmNjtOq2aSDh0k0U7Njvl9P108rLOqcz
jByAUb86DkZhjF3nDLgyly8zo76dAxxVGPAMDycNtaM1A84gYI1+1raeLgCxStcVql2zXLBV4Fbn
NWaPcx/Nf9zif0WeFXoKzcmF/d3Ngiz3iiEYOtp+SVXfQ/opMSQcNV4kN5XxF2UJI7HSnhb3HWW+
bkQK1Bgjoq/Mf9vlbsalKnMoLOhVtSWCZnrcHrGvVMbgoG5I/djiygSX6WUJT5+7IiCmbsaEI+us
qYDJlg1C6SEHWFIS1sop6MOyxHfx2cQT1cZCaBwRzE7RZNSEee/BeRupBcs/xefhw0OQM1S5RYGE
ZPh0wGJW7o0b6t1bhldm7RTQioWHjEOgiR22v2rlj33r33cZ8IyYx1uLcbZHpShpREi5/O1ZPS0H
eoUvvr82rXyaHGlWutkmcf1g/JI4oYsCbTJdU6QfeEY/QYGQMAvyiia0NmxGKvHwuBiepcDAuqdB
tUBGJH4oWJKS/3gmegdhcwHGIQgvmbF7l2wmEyTtJNfBc+gM3SvCnNiMnwfdv/g0EnLOdBIBdw9p
9MQArq5AiIKnxCI1HRL4ZEz6KGGJC56amDiWBz0rgNYPJedmP+n3p1WISjwVBPXfYY4gc96AHg7F
FEwq/xRsrTPfUnwMQbXfE5uyOFh0bJqL/itjfahdX4894wkv6PBXWHtvB2DuY1Sjd0gZqwtR0kJP
2DaPFk7rJ0rEUE9TTET/64Su5y1VVJAju3ntwwQCeP0CK2Fc6bb5LynNwSA4A+wcKuaZEsXf90BJ
cwahXOtQ7mK88cyM4/gHzEO6OjRs0svNNipvSpKNJ1Q4zsy5Lf9ypGBZfV1i+Bfqr50aYrjeyfUs
1gNxdTzmkMOCE9/eTTrup6eArCvdLWVl3KGrhDnwBdJuGYC2jsy2pPESFqJdjYu0jEvegcvBAsWL
IZM3CgyF7pANR1hdQjBCVl/ICjNS+cbKW9OLvxeLdHLx686u85hCvzy/AB/Jabl9lAbVMJH5JdIT
wazf6UVpkcr7Qtr2zHL3tLU+tqvyGKIduQ0OEMRwyRWHI4hYImnzBdkKTuqJz2ClqLz904zql+TJ
Gfhq19zaa2XtvRQgD8wUtvtVcv55wsVtZ0TEJ3DCak7GVKR0409HS/0hRlNwPiUaCGd1WlSyr8Jd
9C40UfPf597kUhoBm7b+nOKD9bj76PiQjGTMkIF7qwVuQx7rbV6z4lbMD5IEhEXPD1dnKdpN4ula
8KowdQlri3ZiLFdWO3HGoNuTy/A0QQGtfAGbk7smxlokEoe76CggEY1SwXrjSMHMg3ou3m4ERNF0
wxOCB9G5YNSc9Uz8JsH3TdlU5g5Ed2pEFExiz0XifPoPQjjEwL4V9Em9GPq2lJV5n2dyTYM7nAcN
dkJLSxeau6+/ZKYpjS25Fya2Vye6pkLpFzryZZy080Xzg0yK1QfH2ViLfkWTOr5su6BABS040GBN
qDXo+KlbPqqjaHGxqRjOQWpwbrPvifDQYr0+E/tATB3akXt/G3D+3KdcIrRJVpBH+Uf4oSLiMufo
psrCbnAcrS0l11VuBXB9wtgx75VkbhThoj/KQUFQdkC1smTPdiq22jwFBAEGqEmj/geUW0D7IVTS
+LulQvH6nQsP1PWU/JoW33GI+Fmr6kAg4obbGyLipWVDeYDdUsCkg8kQBHNdC3iN5iAmKwLfBdLu
eo8TmrR6aPjybcAEIHaP3OcenF2BY0364GcnLDxkUBtN4fmcr/oN4YLT/vKroiYO2GTIaWUVnCgc
158AHk1m6EuRUFLcSN2rMudVFNF8F2ASkBVLdV6bgzARPD+VBAR6myZSXL3Zrio7VGDUpMnU57Z1
Muz25GMt7ymU2pF63rlRHccDerwliVWOt6csvjpGYpwz8it0EpVlyDdxUzpRcBl2wgQ/3NNWVKQw
1KNhwo4cYfw1KOOkzR1WeaI1oxbK2ktfihhbX01enekkgHgPz00zgeb2viND/6euzS8QDQiZJBTG
W/5FjNt75YyXbGkBLupAheHGz41Arob5VDefOjQl8syCf3BG+ZyeH02dSL7WAuH59l2sfkMmZcsZ
/80WR3Ken58mr6Q1Fz3g7sOmdqLBdbpmlP5/O8zKnWA+qtsELVCS1kL/elkbMQwAeQ41CEdfwD4w
wZsW5Afpf/OjcRSw/ohA1urLzYyDLa9Sp3ERhp3Ff7zN44/yLIchM2hQaIbsO3EbJUn1Rb4nmcKM
phCyAwE28pMx2GoK3rvgY33kPH4Po67IPAIpiFkh3lScpkl/rLKqP8aM3QfVi1UeOKici10mlA4o
z4rggeirklozI2L7klriREnoGsH/2BacJNK3Qo5DAUaeW882e81920Z82y8dQRPwt7gowCGPNbPW
zVujDj6iYAmLTUWUA0mMzcSlDussWToGMe8t5uLvwsYVufR7+vbN/2gszD5dJwmGS69t0xk5GL6J
C2+LBY05mX6FHBUoRTKCY+DW7aZOixs5pE8I6r9CISCKln+zYkIo3XgmjqK4MF6Rr4I8erAnYKAR
Uac1puj9OjepXDC0z9odmvmUmTi9Ki9iARps4oK6f8BeYqH3YWYr+ipB4/zGOkors5WRXm1oFieg
2Mwy0VluW2caUzvvK+UvLTAuPWi9VR6RDl6f9m8LfuXnaT2wfT11dVkHhQ3WceIDUnBt8i39hEeE
QlF06Q07n5bhuNH4LMqG0wuD9ouKJCT6jmNBN4Ih+Mjs1YWH5FkjoZUWLrNPMgCna2VP+x4CP+L2
KYsVB3XWcBzlc/N4yf3wUMkqpnx7/bJ1Hi9oR4sy5Vl6I3dnkpgmStmBvFv/bPNvmiQhBhngQA83
DEflwTzwiquzLSFA/1aREu7c/3Y5hKXdlM5Na0nghr5rLuQyhyerJvFi8ZMW9TIEM0S7UbuRyOLR
Hf8AjRYCeo9GVc/kpYmQ+imvokTlThx/HeiQMX3xtvQB1W1fy75W6UYpZtwSG1J+TVpskRot5660
9B6BzsYS77rajnSEMp1h5maet0KQSbY2A0sN3n76ZdkkWw+ySrl+/g+B0dkVdFOt9uYrtKp/ATw8
OyZC4XwIbXVvJ9sLasf4OtPlbapOjpCXhdRFUiVqRARynAIShToo3guQZYWWolmzv5G52imAghJQ
4/mP9lAWCFCfu/S5htJSZYxYv0xWG22yj4IwltWkpnWICBIRYa5FDalQPK6I5f4VmO2gTrVPS11e
/INWCLqD6IiNBd3u0iFi2p2wY6e4Jsp3BVLxrwrvEYrYHpeveL6MAZZjJXqqsbVjK/HCyCO3zxe9
IDDnYDp/lrGEn7VwZ2L8iKLRCWlnYMfz8tgcQ1N3c8R2hk+MXD5rf+OBtkf7gacgS6Qh3gFv9qdM
IwSvNjqGTvWp3cI3JLKEDcUqugOrTbd/3BDKD+mk/uWg/YCZ1uX62MuguYmbRi+V32XzKDqjjfAL
CwwuBkireeKesfrHxAZE39emf/zlbjgLLYi36M/ju7lUu6TBNClm3HAyMTKGNARdUtf32cOzQcU/
2LVrwrf45p4T623svJWOnhHzoWzJSB7FQ/T/5jLJKbqlDC24GPoDfvmKS8/+NdyCXXseNr+XL19p
wieRVFeH9TPjbBFxne7jPlHJ9lVycAZNaQ1m9UD2xtQ3NcWYjShqFCpXbN95pX2dVkZwaxaEsXEC
h/S6PmRiyLNemu+/z6SJJU3iTjRHZ9YDqTkDbJpnDpv3zyR9+gJh7Hg4aTkkX2fCspxsFGoTcR7Q
EGyVo40Gn+S9+8Hni3cIXlWQq4t3AdobNOIWcusF2njZ4gfF8bVajCvA4MQEvrllWNSgbs9rF93+
/bS2jkBj9XOzTAkqiB7YqX2VKT6ecGsY13hJQt10nnrA48jIPBtphnvVFdSgBMJlRehKZ8/v07R7
sMMJ3p99qVrqXfgxoJ13YEl6d9AjVNQBR+VHyUjXDKvM7IiWUdYPDsIIPH7J0VD861SsTZTaH4Ip
K1F+hnOwMy7x4DBN5iEmEf4n0EqIWpjUEOr/HEEYLz9yDq4xLsiDErFAV75omtc/VyEVcwaVBFnB
ei93on3c4sVLnRCjL99sRxMo0YyG3kOu3zRHWsHuiDYBOWDpUtXfn9puY8SUwdXOTJkll9Vxfskg
ve7rVHIvp9GaXtRqpTSxABeTLWCM7tTxVbFnKIsD4Ou503CKWQ+eKnYooPoeKZmd6x11derbL7rj
ygtrkPT0jpNyGxKoMu1EPCdBLSlxurlbqDRpymHUu30qbvzJ3evb/bsmsZSeZo8ATGribLzpRFl3
z02Yma0rrTJJoMacj+E9nTIZkuoqz/93pMzBq8QVySn9ImduIf4rZ+0d4Gl/mqWQdCiLqbOvxduh
eTqUxt4u9BCmQuFep3ji4q1pvZk7LnALhiOEjfcoXuHMnYUi088bp9KVH8AUyjYrLWa0jHaHOYGS
Ps5hG62AMmF5VcXptjC506+lamopOjLaURjqs3X6j+V//cBdM5zeKiM1v18cjYBiQqakxCw+c756
vQUc53XGkR0pkEI9afR+ZmbbD6DQ2iLoWPrsTO1cG2jU1i+fdV35OZtXVRHpLgiaBj+RgQOB+kJd
GeWic8wzKUjMFOHsGaYYcuJ5TWjZZaRbjsBygbVFc7LTaNL7F47Dw5EiwMH6NjxSaOFROdi6FAsG
Hoe7u/rAYNVop9zJbjYIyBwO5yvPIMUqbzPqZCJK9cBpVrQ9Bw6NfkSE0f8odMCEq9yHIRZkN2UX
IPPk1Lhg1B89mLX/GMLtogXA+ihpkqtSQM4Jw60j7RSOW1+g4Bs+81TTXShw0gvEeJDQ27CLyyIt
dkqKgQgKhF1g0LABo7Y0lspCTeKIoGhZ72L1QfPUWfA9J61jVKr/Qhy8d7ItKCaOXee1+IfVAdtO
xQEWuW+511WlVVqoxoc82wWuej3uCynqUWsRiy7Hs59g7aniffi3RUdynRr0AxR9Gedyp6qVAo8u
68Dyv/cWbFCBRqBPBHhBYh7AMceS2n6eLa6jTi/dOLGtCQTvA44fuH6Rqzjh3uDUo5rQ/ikOSNHj
J5bA+yjhrXybhg0V/7obLqL40E/Faj9hiYUHkQmbc5URxS2Ojc8qhRNcbG0v4P1EE2K6HXfoQurw
4LoaoLiuK1S/mZ8O5YLrFVtEjKAJ5yvuJREJCmIb9/mdpPEWgJe51ks4/clE9STcoyJMQgoWAzi7
qvV8kfjjYZq1bOG1cmYpRZjGmNl4mHo1qY8U5e1voacGTbz/D8aZW+z/Z9opZtCihWTe8wlef+jx
gydGlCnfG49XdFNC8mIzn3bKqMXxRGsOkIMkqXyijudAcM0Zv6FFiYfNJ6/C8+x+a6E8b/R4/jL4
XWf9EXU6MUn2n8JnYUmEp6BVPm7RUMIPh2kH6fdsWfyqhumBR1QHqbxquJK0vLmgELALZW5MDWyZ
hQ5arcSOG6p4NinKK2zNxplIfni+OqnVK4rwGncGtY5etCz1utrH14LcLT7Kz02pqTTLWMBxidZ4
9visQMGl+/qbnGiUliOPXeZbYzkb9hgwW2USFiSwCI6rZD5EVuH5wQs7mTKo+/y7wNWPFgXw/HKL
HBxwQ4Ss40caYENRhP5UpgeSttw5/VdwrkhLK/gcFQuo/VfywzpeWPkfba8/Xtu2rc8MgV+CInBL
sHPczFgQoy6ubyQY0j7O6uwgxMJQQ+HHuh+3hYsvbVpuiQxJomH0gf+7XvfA0BXSAjldk++Rmcjx
eraX0F3z47vhcz4rMCpDvOfMnvAvk0w85ivANEvjeG1PuZ5EmYWg+YSDpqhK8g1Xt2LVnz44DOcA
xo6qSborbvXrrRFc8CchBYoq7BWGmZu7EN6TFTX7tSmz1MHJ0JRZmK8Ithsp400K7+yb7cIfvkYz
ZoVHxaojbrViyEzw1vqrtqhLsS8AOrwJMVyvrGp1qDXjND9QMFgzRWvHogGXXCUVZzvwTPImUeMq
uOF/xw5fdYSwYyzFhW06TcEjME1bqrLJZpu4unPxl1DK/3O0J8HUqqvLnU0v+dVgEf072q7D6D4H
U0ybUw2lDOyp88mEfdpnJByWNtibLdo0bfhKveVhPPG/ZsD5XTb0ZqFuk+TxvV6xsRMvA3Uqe1xu
9mLcH6oB+OoWCvKgBIRg7SfYetUeH2mg2JE7zvBfsJnQJkxKSqzfK82iT5x+Vv7LSGPONBHLzY1E
XTNzqYiGERJgEOOE2OEFZhpRm3zojfbW+9uKK0SWfRnusVEthaF+XNw2adO0fva6ep0kZrPm30tr
guZL086uF9IILHtrF0kK3ah3Q+qwnTcx7AGg1hUFX++m97NRFQnYUdztwi7FzVJVI8GFiTnY3ghV
UMazoZbVAEdLTnU++zrH7Y0E3p+l9HAt7/z0OsILoAt+WyiZIuyS/RudV8BkPFi5uOrLUVhVCdR9
IlG0Wal9r8RfbxltPyUQj5KteqM+2oehvi+hraeOsuoTxg4GHTxiLzkMXRWeSPu2q013L95R760Q
Efie7EOlc48G4H8vmjPKuNIIGzwWcM/2aHZIMxhh2FcUM+Gy3eQ7GhohuYDg8yzyx59dbTN3Ybb2
4j2jrM6q4UPwaGJgZ2JTpJA9US4WfK7XdhjY1ZbbO+25cJDQXzfSxxiifC0gkpwaMKyjr5BrHsC5
obpR6AmjCLUkayI4NuwOGn0FhIvBQr2aeMFpeAPogWwsBEDoq1qknCIasdO30i150EZ1/vSMkCrS
qXoZHBYyIkEFDtgkzTZFbK6+ge7XnFu5d981A1KQIZnMQLpr3mK1elZnEfLmLLe3InQe76SURabQ
KLvqg4GiMWaWs497k2bDMK+Ee1gpEWZU+NpB8Z9+fzh4uaFu20bj58ZunBysHKOVXxq5eEvgQHcL
71gjENGnWgS7HW7XMMwpsPUeqLTaeEol/i53nrIPnxHdqYILLFedAaQOULpkf/yPZbRhwQ/YTInZ
bI7ukzju2/jaE9c+TMkkojLYxi7Ki9vO56dBJjThMst4QKBWed0mILK50FfDlxuB2Hb2kxRmeN++
88jTcPYS5Q7JQ+QDc+UljPiWsGtiv8btNW9F8JmYXUkoWdqhiWC2dc/vZmFW+QSAWZobqEtnPvut
3CzUGYAahPdKWAPaC5cw2i6p0LSw/eXDFqXD9fIFqP0KlDusDLKepK7Vut9V2M67ufk4G+R2E0EM
3XBVMvVIyRiDAC504kYsINaBP5d0VmmsAJV5DVGjmL9bMHenGENWuXp9yDgYF0bYXOHcLkf+Ryvh
CcNQvEKl+cnTlKIahL7X4h1xOvrW5hca4g/RhuD87SoDViHsPFLaYPZJSbJQgU3cH6cTv9UnfYK7
+04IyFk441wJWrqyZ7tdPu4lrbkZlxO+yldzWVo/TFKcr7p2X5zegB66hz8lIjrrMo/dk/DU0lw0
93Pdc7xADF4BItYYupMAHnXeWFGwPkSOZxosG9MP2JMvvz2o96EdzXbLtwR6vrUBWWC8gJU4Hhqa
AyYXTOj+jRo/iD+JUJlpgMhxlAyd8IXunGG3aershSj0hYk8yCHINorjGYwR56+HI2HXSPncGJdw
O6RmkKX4UJMx8Q/GTNNSTeqXAjYj0pGil/QSR9vi6R6oBv4hB9eWd4z97TzK5wgpu1iNE7Kwo7GJ
CXzjWNTBmFaovcZhBfwmOOrBy9W9DRXY/MKk04iEzT+3/UJ3SYwhTqgLRQ+EuCklrVg72kuevDFh
dd7NZIjGS/RGW+VHpUO5gUyiVkq32FAXVIIfQCnZOB2l5DoqvCu+yDwwuttHGudzGiHKVKDEd00s
eI+4qC7b/NW/zp1gs5P0v46/7ySym//RjKGByp6f1l3Vas1DCWt9KM1g9XPWA6boWrg4f1ViPv3h
vvednTbGi7tqWM9PoFYFVcz6ZtRGCQU0mssmCGjDZ+kNrNJmOWPIbyYJ/dEUYa6K7fuHG0nB1VEy
wPz+GKS3dQEYRYrAuhX9NLA2rsEYvqD7WjPPiV7E35yi4vR45BcdJHNsG+KhIGQPTXzCGDVDQWV4
3SflCHj/mYwJLGoNyKH3IUNSW8N0Ml9GsSX6tqRqZBAdKOzP2LtZaBItI+ngOWhgnOyM2ivhRYKo
iBciNhaKpAL14GhJDy4KnM8+/C3yna5N4B2wGr3vfIiDAuTAq3yDp71LA/1Bfnyfc/MeyIz9t6HQ
tI0x1M+dzK+HXJnbtwARs2A5E6NCa2+Gi23wCQk7RYH8wz4h+Vs4Nm4GT6+A+5NhL2UJJhZ13P66
bK5FAheq9DBkPS+zhkIxDCk4IoUji7JXUdaWFpg5D5KvU3I5D3PKkQXAYPFmIB5e7T8RfnqbT2sg
kf6P86ZMKXGy3/Tpr45EWY/9CSL7e5fgouUSW7jU5aXXLeGZw7jC+SysSQmYbxmw5wRw+XPxnCFQ
T5rB2XsY5YGHYs31ntA8xdUAtKLsF92tsfaTspFIAphQ4Uf09t7LQzXAqwcDeN69dLV1zZ46kOkI
KQ+l7xLqezIrhoG9mKAqyvpS/P5BZUBhJYifTXB5O0Kjcjy86PN+QpXMa9d/FRkELMM/6c+y/LJo
KH14MIE1vBpWuycwrFn0guPSQ2bCz6sg3uRYFwmvM4h0LBo60CLrdGYvz/uptd0uOYNkqos5aIyo
Bb5uLaKYFogu+qLg56AunZcv6lubg/2Imv40BlwbVEUhVbWM5OEwlDW1zv1jmMFmExkHLTlvy+Fo
GoIUMHSIBWom6MAcmGtGNk3AfPWMAF3YCCYbCrS9RlFCNPWE82STWOISi7C6gkLjO9MB3BwKI6q2
Uz4B+RKnfSCgL7Q+3Ptk2UbEdz5qpWWqosMnthB4vjxp/IQlUFE1VQ3d91G3oQAthOTFwW8uVqni
2LQJc+g9urCVvtcGue+ix6fKigLAk+ocFY0B1XQNrppv1nWCWeNI9VOdM8SCbMgpQkI0GhjXAYgG
PuUH0NexQDJNTUlB74sCFVVZGIx2PQecsYF3JPn0TcEo1h6qPNF+4uLlk9naaMT9l54asv3efhM/
b7PH+IiPVVZQh/G5wq46dsiPXsxQLGGQBpeNwC9J4WFyXkZb/Ayb8TmGemSgvlFx7U9BV7JRuCuE
A4+CRF1L69E1/kh38vQCTkeRs7yP+/43xEoQVrOa0UGACvE/VCrycc70xmUbgQ6BYWoWHnPfjmwj
5axNd4+QhRwwhh69EtaKY1nLMb0dWTHspiyUqEUfW7visyUXRM7I49Swbg/AKIrHgu0F++daxpHP
oKTuyXO8sdhl1zlZeK23kYPLrp8Lee3Fcdk7YzCoEJJuj+f8IylAE17KzqZHpO5bhLBDQW8ubggf
IQbwnT83uSWrD3/KuFEpmX5O3xH5JFhln3hn5vvkAiKis4CVHV5wPd7yl8HrN5cTvinliXydnXC2
WwE1YIlsNXG1ENAi2Cn6SYzG2TcB/uOki//aIyWSRGUv9R7peLbQNFua2xSPMSzicajoROQn0M5K
q15FVITsiwy7V+5K3262GDSzpJ+lQlDeetvj/HwmwSB+FgKQuVuFWZ/TWDeKYDGrCciq8O/uQMRb
siqx4TPQaDKaMLxjBN9uqh21SvC08kU7f+CIaP3iNVgGPa5xDjFl+xkyOtgIifOh7Gfw+ks4JwNK
XQ3mbqXwVgA/pFTtGEfI4meXNwrGZZm0bya2fLfWzd/akdHnxFlKEdZq0RjKG8NdrMPZk+HbaYbz
JQaCKxCFxineMCcZI/bCsdX8pGRNaFyQj1t6VdKTdsE9Tii9fgPjfWXhkYGTsWF/AqQhXiWEs1GJ
VLvzWSBiteTThUPdV7/42jaDLusyunczUbD4+UPnMHDvdc0cWpLExqmR3JeHPhOa+UXYHqB0O4dA
s2fNa1PQNeR8CN8/cnIk7Js64kDv80MJ/s7bCQ132jm/mUzNKEuYdufNItfxHP4sRviW4hAZJ+zs
eZXqQE2x1TwJoCDjh561wnGquMPtk4G9d3AiOkTFDy/yuY+Og8ll6lDJaVH13vN5JK1BI5JXN1aK
qmXApG+XV+OpXEBufbLPlJZS74rVv7+qLVFKqfCJ5IrR8vBgqbfzMQz+I2eiJjS6TiUP7F0bK8zt
WEJWCmY32/rzAUv1JfiUuUctwrRblKVMRMEjMW2rSey8SvP5FguRqx7W+9XdDtGXpW2sDeLbUkxF
LfwTFpETR0YgmxzGg5xLC8qKhALYcZ8z9+xUDZO2J3HSukT4oQeQ1rBNXSc5qrhc1hUQOCRHCjJc
y0s88hvz9JUURhyiJWR6EwXTfCN7kuYvD3EBFJxiFSYXCJJnbgX65BVzrnzCXAO2jPP7tO59dpKF
GzRSPfrHAuEajZu9hoTQD+0EYSJJA4R0TAXOPWFlxHgzbK35q0TPGQ3iMmJFjwdfRAuKglBX+oM0
rhAs94ENhi20NgWPNCBUeTew2Fyo6p0/75JSzvAUHdLM3lQ/qDJ/vw+YDL9TasMxkojRDHxKn7tr
1N2eRxkibNSx/nlHmH136Zy+DC53y99R5wuG1UYVnOBYz3Y+Biw+9GrX94WopgjHpJRTmGcC4TmS
do7l/zymD2MypHzydYRTvxtaKw0xwnZMZUpXL42ETGxPHe3emH2kv0LA3uRGCnjiPKk7HWQt21GX
I1areSxgp6I3L+TArmSlOXsL0ug97M3K6x3MMopwhzYJvISB1JJUXRXgKeCt8wJ0x63cDXccqYqn
SLjV8vvk777URKmLQVJWJXsgNmTMavp8sOuKsthOGR5laODfOeIjdrvKlTAgoI7ckpW/3tA50nyv
lgSKOV6tvrqym/9kctjxzXB6CtJdyux0dxSfIY++BQq+pzMejiych51vbekAHvl2ZBjKdbYf3BJA
rWvvTia6IuHIcsaJ6JcFeuQxqoq0AMCJeaE4umJNOBuPGPNoM45Z9jvt2MTK8lfbafJGAYhA6/eu
RA29PAzO/xZW3U/s4vZgkXJeaaZwRRom9R3EBzaevGIjUf9rJqrclvS3pREnOnVld1SS7NQYHWGa
zlOiEkL9iN4Yowrq8rk+d+6HDiSTpeQvKco/Kof4jz8d6tyA8sysJyEZ+0ZKyn8CtjbFg1RQRnt5
v9eHALp2eU9hUYwGd5xfzXuRivXfdfxzOCUTznobqmFg/+0BjMnb9Ct3Q0tRuPkpqRFwHxQFMl+y
Ivo8xhAscP2mFgrsvzIfSGI8SU8erMQ61LCoKzbVuYETjnSHjuFCQEmqO2sWcY69LJWA/Ne5poDk
jtatTWfqkrbHmiMS6zznfmpUntQS6uNpYlpMVijWUee1rQZ102isyjzq98XmbvaoOfjjI5VT6X2J
aeonp0I00k4UZGMojbwiV/BYGyvs8JZC7FFSJthu2tHh0jKlNADJAN7ZUsmZnsQbks2L69Z+BR0d
PQrdaobiyE8JMOt/oKGGSIP7Pjz3asnKR4HT3aFpamlh7fQO6Op4k6A8GrAxcvRcMR3EJIKVGBCX
/2/mZIVkF5/1Sizr+43fpMLIkEvK2YI+qBuZTkAKz+0HKJDJLVrBY8fdOirQH1nscbpZ6xdBg575
r0X+oY2OTgtZdLD6HX+v0bBRasnJeFWVD1aKENMMh3KikSk3lUIKqMVtdOSjPJ9OKrv9rAIS8vPJ
lrmcg1tEeuHf7q7KPECShz85vlvY+nyrH2LLaN5mXwSkM4JpOy4u1V8swvtpHibnIjF/J//lD9U/
lWxsOYarIR09RcEVtnUMbvPUc2WyHjYkrWVUMs2B7fsJ7aj4CjHs5jk1ARI9Id4J/5DjoUR7FiYh
ugsNV9byGcG87ieI6I0RBXuDVsHY89Wp5KzwTYqSPCcdQow0gklnowG6HEDHDjPlLrL8cMKewnJY
sj9ZAnrA/j/ktCS0PWwZ1SXc14fx4RiM6p+236Ojz1aA3dAgjh8ezVeK0V0u+7D5PeOKHd9yTLig
W7mP8eyyE229xNFVPEWkmRBEAVHZYU+ojdDEdMPrLznXmEJWPbfXETgWTjYw+00rvPE/T+q6c0Xf
ZxAZchLHFPB9Nzr5Br9OLLD+ld2h+/N0lCf99JHM5KOmKBCg0Kz4Ylmbw/jL5TWgNEi3fviZkAUG
NwOHNje8QX81P7Piyy/AGy/R5kRckCzdGgz1dDQkGfgDKxaKnDubSFsO8HCcPXVlCtMy3BQfxoiv
VA98NqRzzbnNpH/LUvWem9l+VAShKHSd0Mf6NYvjx3K6AGJtvIZJOOGxTMjDqGs5TaUA39jFKD8L
ttdAqdZmMQtaloQwIOP371yX0TsnYl46qV9fzJGgbxBOmbvIJJmaqFXs4FZzBOV4wF2/AqoiaDyd
eO2bh0hnSEpeKRUrZNQvN8BJnwjeosjfwoBVZ38w/iYaEjgDl7DIF/rXfO8tGdTYzFUHXrz1IBX4
PwzGEaM1sGPYn0pKPgyCNMqeadzj6zS3mNxVnYGa2s8HvnGtE7CzmBjKOkgUNBQfov9ycjUzZ+Rn
VzSQlm033FHGmcBdASNne3ZJk6ET+P46WBJFAHJFcsBy8kWpVQ7WkqoF/GAGvflxQ/bXITWmowDn
kNuNaUEe3JiiNXLU9T8ATJx8TGTc5oJbnYTacAtnVo9Ga+7qNesMtGkyElGO7Guo3STOiY+r+rtE
QL0ldYToUalQoKj7xtuNjeuuJQiV6eRGsninuQzlvsdl0g21QJgcgLhxgLmxEp9pkQh7/0Shcakv
DV/q2iHaycoUE6VCmJ89NZiWiZB9FaI8nSqYCptE9CtWgNpJhwIYO0PUXrCNrtkGb491NrhTq2aT
eVxRLqxTNEHDxufdi3R89O9/vy/IZ43nMPSPtBKEkVzk8xrzwGC4s07zdylMoD29Sty0OMT5GpLr
EzZddEL6xlJ1hvGgbespz19NmDHhod6LrZGRqVvt7WwMby5oUNqcM3Pvrvz3cZURsje2E9Ii9R2b
I7Zruwt4mHNC47GY0FLzpmI9/7JKxXxsNgOTEPdgwro8XS7MCHiTppaOIwnNcqwN7XS+tNSTwYbM
H1f2T1+YSojqsLoWvEFSa40naizILVquqE1Tcs05D7p3WUFglPimCYILGPNjnfCTF4YgVlEOGygK
UKKFH+xgshyZsOQbUEhxS6ynbkeq58r2Ysd5OGrvaLwEdVuQtbgxoUIYsvdbgEFcVJBrTbL4/XSd
OKkD6USLW3RisJNP2ikrcPT9ik4+5KHt8mp3P7ferlDbkf0m3jjLmmmFBjP/1fsFOeUdxh2nTVPE
k6P6HWmT5KgSzd/ZhwWdPJfooSzMCS97V6SWx/vcFZdHSPvIut3qD2BYppDW9DyNMPOxzMI2cu1j
9SgeyruzUPmFXe3DwMUP/6aoej09xP0fpnYymUuBVpvet+bToAwbQ/9cm5SqQqJIpRGxWu4NwMjc
OwD9aPLobqMXUUPdD6QQsNV/GEOcOmQ80Hf8HxSfPKXp5QMABSiH3ep4PARTSqXNidaB6KMroXSx
t2OtQSDA8zuGvcrSgAICXP29qJ/usOsl0WHUZkCegNo2FEWi+cfnrcGLQbzj/HW8FW5kJcdb2kNO
eNw6hKQoAHfLY7yCREk1U1Ut18mpbspQhlAr6UvZI8aA9apRepRy9Xtbv9CnuppgHCZMQtxVxF4p
meKjFsGFPQ3UZZxoVT+Q7c7XdynIg1K0KI86ef09B5qpFFmp+doSJCR2ugSXPp09qaQjR6HpUX0R
TS58h7T9ZnO11saDx6HiLzGDIp6viyfpynJNukkdBiKAscndF3nhhPscnko1BryTvGCQqfN6tQVD
miwFIHBZZhrkZB6KWK1DDWe//l6ehjavc/Ykr5i2bnM2AnbS0anGGj2gsn5u1EaWRRthj+615RFs
wKbEykSALXjIzmsE7Io9M8oeVxUZ4Igd0fpN0z5wfznwqjAoYkkN321nO56CmTf5emVmv+ZK7b0v
LTCbbdi5sh2SHQgfeoVAAuIMRQf5hZMEoZ3csfpX0j0YOZ3FaH4+WY7kK0o79irKUzxyiXFWetqd
hCQndxxSAurfXFWmd5+5jQmR9z8R8EcY0ETqcKauVuwzbnLcxexp+YJGEJ7QdJl3mCkAsMeSE6Ij
pE4r2npNFJ5KgYdHXiNordjFGqk7TNFRZHS8jIWRR1IbuguWYXzHlEAjR5yTtow+WZFuSaJQv4Cw
jlK5uObQMXmtsT/S21bIWyibnTuBdrQrChXUEkC8UTsIuwMfouCU6MY6FF+iLRZBXxekWh1YewR8
qk/+IDXYhnwdPHt5cB0uIcR/KML+W6FxysODxyTPHusTyAqLLJwdrhc3OqkSKOCSqWFMmomN+P5D
0+qtpCWQN9609jH5gQobupBfLWJ/T347NOIqwia05lRg0JAL0l8reju7GgAvf/Js97pyM0xrt3UH
yl6Y2K/nbWksuYt5lZNHJA+vmTC41eE3V3FFGw3aYAuhCv7rTWgiTuY03HifcPH+BZzxbsRQCP5f
5qmVFUVWClkYFTwyYI4PHgiINnAljPLk0MrH5MVwtzY9reyNgDmS9Pz8YG/xlSaq9fqKJ4U71TMW
80AM3NDA+p4fVq8uHkrrImpsaMPd1Oyf2w4MFNRXA2v1TZF6SocupAGoECGrqLY/fvcUrkLfcC6M
gKfDmDdrj5V2QHW6wXpcZ7ruSXTw3q+ATe1qVKd1+KdFrR3pyxIWRDHFIE66ilqIw6hnLdzEOkLj
1vKI2EusVaaBrPzVgaV9JpVg3Vnn+zL3+iwzsaYXyUDSoiT2+ZhugwcFhXqNePEY6Jp6kh06SfA7
eBD1UdVi1btOS73yKrNsah2RCaUVlF2biSviTHovx56g7yD2syyUmWAYB2Qv86He7+XzWRdeLYFv
l+moxWXAKx80R4jzJyqJ5tModMyvabjktEZcRq9e8MUpQZ6XZVqNMxUXP79B20RtUnfNYxgG6xFz
QLhRojssR+mPnLL4ioq68H6v505PE7GMoEPqbWG5/nv0Ms6S74sRAjq8T5PoOfDj+ruVxWS5tyfA
uQ8jTC9MrnCIXpjaqhe3PjRooT3jb5cmPaCIQPZIzU0zmMGjcj5zse5RnjXSbYyWUrngxm4YC1qH
HaZnx5oGCZoks5EsyJqjVVC8tlBBWh+IfpHukwtcebJH3UitFeYCu4T5612fq5NDeQ4sDNQhg5vo
IHHA5mqHknodrg8ZHBxonLFcEeavzI3W6E/YGw6Q69Mb1dFOpnAjlVakE9hDo3+bbincazGUxfxb
UJ6c4CluQDZWfBrvTqq+D0b962psoa47J2gkDVGGhgf/G0qSQF/6zMvU71iC6i9EjbqAGwwlggWR
+K1AW6G4awm99Ry/JRRR9hQRKrjR3FdYnghYobBnTlDzt1Vw1T8jDdFFJ6KMrXyrtlu0ekPCu350
Q254/eGKf3vP60rxkcXW3dm6Kc9O88Vivmf25ftS7h7FT/eP2mDV5kbmVT+59vPTwI5PKehQuwkz
9R9l0FMSNi3lEgG1jwbQsq8ZJWEPdV9I41WxZKHCeUuhvlimYWhiBQUSchONt6xlFuJiI80UQK2v
scfnUEQRgUBSP2BOFgXA1O5h0zbpt6//Z+o/87s2a+7S+B3vchBbsodu56McEVUe4yYIkXJf2br5
RXPzJCWiNj741Iep192WtmW1Isy8K4Zj+nXaxs7v26jeVVIYzXkdkcxWQU0M49mFsYZrQyQWMktQ
z7FEZ8xirFGNc84Xy0Bx3ZOQflmZuyXH8F+4Y5ipDgriHWma3pBDnsIuRSl1vBcqeiKJSOEr1nI8
uhaP8DY0BKGPh3eV6qSu4HupowdNcn+uDA+b1on7BXCTlDVLUZl3sOvPScMDn7vo8UlO8raMUBxs
yxUJFd053PR9p8S1MWA9YR4i+qQExdw6NhBA9gM1MEGP0ooi1RtEYbHriYfl6R9NbKk1p8tCWzjd
LZYZIEcf2GIBfRqwDHBIbgPree6cJAWmFHd+sl5AyRvxLRVO/k7ZTqm+zvvKMwFztq2cHo+pA1mb
ZmYRZoWin556Qkk1m2JdJMsABL9XEk6P2NBUrP53K4zhm3IVC8paa09fQebxA6U7lZuN/l3swMyC
e7mztgaeKPdDLwFrUSUAqc7+xpeZZnFPtAX1HHAZZ1PQB8nQ/xbOV7Uucdc0BHMgY0z5/J0esveS
EXfvnj+RQH1cpdZSQ1nE8wVT/1ZdiKQ4AGccjzQV1aJzh2I94Mtx6KyYIBOgAiwdVIesuetWrCQR
FFzFzupX9bBpYZajDYhjxtFOuoz1Tgx4oz3pCmGE1vaAkbb7GB33U45+b3w5uWEjScdBaEJ4frpO
1lTmq5jqXtXGccgLJfycKEbFbaP5LY4cN8TLxQhHMpJ46rBqo8jhkJSmqJZth28fWiMLfz86HZGk
v0AyEnnyROETjsrOb6CciMCZfocZxb7eRrXDYbVKHBdIuXkoX6xsNv/vjUnGHfCoIFyeuAPBdyzy
tfgDngIcpzBtdYXYq9wuLFHO3/CoQpE0YNO7u0Qk4ePp1qTo94tjlzC1MUDDdHqq7r/eTT0qWh/B
ldwJ2xzQRNfEzrId0vKvyJXTSzT3iP9cQEpReaBW0yTxhkADSGElTWj8X6cpsAC4AaWdYeWuNKLs
egI5J49OqDtuBxlwz74ehK3fJ36hWvcx/cqjXQ4NjOkAqpPCqFqX0XuOQbz6Pagk2ckYJ8eHoWfg
EUxdckEm/ghT7D8nKYu7E6B7FZ9tmHc5TYkFCSUVjYmIcfLEUDrQ2V1LNiBU/X2OKOi2VXJkLUHP
1aszucvgt6QnkAfUCYeKwr13Hhn+74PHWZAXccGw+HAqwAfHPkl6PMfOpcr/PcPFaBWoalTmF0w6
p3luuNa4A8T5ACjxCaLWpaj1n4YU3SiUCVE1iZpcZ0MwimfZ0v2IM92TEy5JXrhXMh5s2tAmAsMM
pXARSvrPrY/jo3MdUZ3KDf+YaQtl/XznlqAZqrOLeGp0n+O4/yZ6R7x98WIh6WMv/RXoptH+z4oJ
Iunmft5w5t9skP0XTwUyaf7tCWo5Ru+p2j5kzxb/z2dc9k8jDkE7nV7Fi79qdMGQuLod7CXP3gOt
XMqVt2XUz5GJTvr1rVVHh6eR+XIxWscJ674G+mooRsBLxDArKExYZyWpnCAwKZdKGph3878V4oWB
/1ngrTKKwN2D77em3YEpK1WdJmK0G2o5un1f5bOb5HiYfCN8caWOkWFSa7l4xQOzWjxPZBnFBaoS
I/sYSKrAIjsg984JTW9iFTz3bXcnUtigXHjFsEvYTjf2vsmywjgzpZZkvsjJ4OOxYl1ePMV4wxJW
+98jpG8pQxfAKfFAlB4U4kzgb2CGh7FgaL5rVmezdjdn9z7zq6Q+bjYyaNlQ7k3C39LphMlFA3E3
/a1ML7ssoSxL8tycbcOIecGARl26fMWutlLx/rz3bo5FEYCxgAsmaSmDbMzRI4s/6E5dLTBJeMXr
GK/9JhQbsA8y6qf4G1eQDi4mdmdqdf4U6kH/zLUZlUQohlVpGO2RC9jQFqDRDTD3L5SYkVKwA3Zf
gIVN9hkIsEcYmZNJOB0L8GzTOGHVb6xkhkCDwWqPO7rq87y2OCpdAd6r0KzYTz1xzPcxsw+IhKIN
5NibRrTzNxi/SFZThjUG+5Mp2WyLiIQM9e1fG+3fm2RFZs69n5W+ecEqW8G5hd1HpzxJNT6bTlHW
9BwKrKfuFfZhG94UrBPAjYaFVqIo7FKiOlFAmKK8gG3B1suNubkZtUftsu/RCDV4rqU4qc4W3H+P
Kpcb00kNy9j5oquzTYjjpK+A1mroeeqjqm7V8iuT6CsZICLSRQRlG6yW+N/+X3aEGsFVzqABk/Gg
DM44ACnvA4cnSRCbQ8TWSYX7Tkx4n6bR722IcRleQekC2+HZPdeD3lluRGZQOaGIO+6ckcuWlWPV
URDIyGlUuDnPzHvuesyGkLP69g3MUbvUpBup9tGCDikLl9lsO4nLbQj2PEDhqtXwuBb52GhkjcBP
dOdf20NcSZG3Bpo7J7/ONIgEa2tOD26vg2qjswBv0VRtV8JZa+9WS8pV6NgCPiVHc0IyEDyxFocE
enB3b574yNVFsdere7VyHk5qllpkuRY4c2vTefh99ZgRe84I5arJ0sI+NG0thut1IoX4qPJgRAgT
DsAHlNHvbljuzUOacuYrpinIQkpnxaerBI6Ck/Ho6ms8tfl5pZf76pBwn5PIagDyVMoEfmUJxeds
vhjHMY0eoZPd2VHe++UInusbL8Zkx8YcWGFuyWaNCfHjM9VOwYLnhbYdy9gjd9x7u5pQVyBIg0bp
TZLA3moETQYyt160ffj/fw4uK6daEPFmOWvY9ZlkVWdDYFpaU6VW2O5htWQuvLHDcFZWnP6YcGHW
sZisOPy7/uf1nruqdZI1tmj1Aq+xoB+VnVpjFVIVW/wH7v7MjgwRHtFC2vAkWXl004LTcFN8ZdB5
MKXItsQ+Onu4ZElKN1azqpwcI/npWdpnUiZeDx9dq+Wobi5A7izI4hs1gh8e6we0F397agCfWIJK
9me8v5bIz1rYL+SjLhReehXwe9VvWz0UANp8Xomx3Gk+ut1/TctkJ/aL/rHVfTbyjQD/Z9mCU5ha
dZgG2daUHPVV99EzkZM+yzwIKWlTN1CWoh6flzMP+XZm+LmHmxRAdyNCPbiUkKQOlresHriTtdHL
mFKisTh1H1WcUiH84kBKDJaCqrsAzopr09eGxUVaDcrPdw3lRzC0bbrn49lsrM+FieSIiA0Z3jQz
UCZV+jp/GisVo4aYx/Pezrt1MofKLeJM8Sg3tOl04xhk7w4yO/7Z7G0J/CSU8OiKRNuAmnkNGlPh
CtzCc/NFF5Avdk9+O/gGLtF4oLGH8TlCYBahIUB1HwNOaQ3KCO+hHVoSMrYxBSOeoV/v+WOtmdZg
1g4cex4WwvKGPqA6H7toXnXrqzfK1dG+YC4NL3WVWQK2kW3B9HO5m9F6QqB0d51OTDClQ7Iv+Mjn
QDgNFyzwL3HfutygEe+vOKeV73ZDkSdoSxaKC1h/9ZlTmZeu/ujsR7Ec0mZuxRzu7YBMgSqyKg64
gHRsPOoFbfElYQJs+SCR1UUsoWTKd5dOLfq8rRM4srjK3gim5vPVgm4JtHkMhKspUkBVZDR5dwxj
W0ORwkpRdWNxq6A8XY0MuGtFly/UVjmY5Or9znpwZW2sV65UQmIAW4vPAf78dX1UbhEqUhOJ2TT+
mx7LCiDVo/FemRmXkbY+S3jniDd6CsMdLD8VhRl6JdvE0uFWdaqRcJcJ3MjT61RAg19xGWOH6+hz
nsXEBxKct7/3w01R9eQw4+1o7QRpRWrgdMcmWIN1ljHxdQCxqmvWAgyjtsQqg3WvgOtODL0jjC53
yy0VmqrWdoYPcSAiYgQ6qp3+9qFZoEtL8TK0XlDYG9fs5gUj0d6XyWnC1U+Ej4kD6xYV+vxoZc3g
vgQPOGUleypjPJwDbVmzLzrXb5N8RWPVy7+Q7il7AsQVzklQacGkZYpvFmGoe1rHq7ADZIibfyyj
A3p2o/unmt71cjiacodBZQghmwVqXkH5rHoylTL6i1KfhdnUsMVvLtblnJg2czp4F3zLKafR1kb1
8dcBP3nxZtbCYof0WPMQ0381l4A40mchS2/bOeqywg2ugIgmAJOVoSQWymVXTeMJh9qxyoqwUy+E
cmShGKDEJMWksMTEkXwe+MntRPGEHe/LlJNjLpCHU/c4rzcvht6+7IDyISbNQqDhtwcAMxGC2hwK
QGAal2K6M873mt8HRzPzWWCBwiOO0JKPKCgkkhus1D1YI/bT1/1Gr1hkoL2PIb+JBuQDx40z4q5L
GEWZtKy8SZj8G7V5eXB2UOA3bTAV4XRgcRYBJKQowmtZnE0pGV7QrRImsUDZCtrrsLjx+KWGH3fU
bPEJph3NkdIlospxLWu2cbVQhPLhQiqCmNE8VhPpj293xfAnxQaOmUxTieNSg4J6+k5nREhSbVLc
yEaBmYR73tDIkqVE67J5gOzU3IuZTooY8HQ6F+4XLEWH4T+26TyzTtWAj3r6aJmrXrCchNi42YfT
XTUcyE5clBOHTXXwvlQHFqpfYFLzCJXkdKEyEYKxmZU6jATNsMcaoM1fDaS8HBqLPjAcfnrF7uSa
ieqoF8ZvSfSgPnU6y8137u3UH7qQSrfD0wINjiR3LUG+oO5GzaiH3ZcbVJDGn6DTZeBdwe76XZjA
j2y06l5luAi4Vc+OPfqdSJR07DZ6Wcfi9zz7TpUtBAfgtyqIpa6OGlrYUJ3n21to7BYkN4RivD1A
3ek/KGmDIAlu+7nR2RXp0fW6zsgZSCqc3VY9N4ljREPGeJNCVijGYWGNfZ57yOb8YAJtqEcQAhSS
UyayyZ2R4XoX/QPm6uARps43iHuUbLozDzsv7BCpT6nqVgMjy17IERDX35JzS5i0lJIfw0NlAanO
WySnOblWhbyz0mGgdUPdpb9N3fdsUChjgZO7tPe2RqZjiDm6quoIBwpMTEYqwNFOhLgh3jg+MU/P
7bANo0H2/JgG1S87GggoReijo1LttEoK2ZGDy7LRTxU2fxB3unN5Jh7wh+QpSitE6k8Oh3YFUCGJ
Pr5oQij2/Z93VGHTCGvMoy8K5Sfgy0eVLO/+tlUetj0Svj8MSdAbz/eZR1KLzlBZm1FbA5Gdj8gR
WrPGYAOh1naPWouvHdziMzWiXIUZlOoS4L7RWkkPZrftMaZwOB10GGsqajW9AcCx7wwe5bKgosdS
gBJHqeHtq5aWYWHM64xGetglAwB3K0j7HQmOAk6Qppz+L4R4P/9z6MS9/wWuxp/cqAMabYsGqKSM
390yU/GHgt/xvrzD7lXnmrLg7QoH1jVAJkLCBlgAj+ReUbjYstIShBEBBcmuI2UvFPYMKsVx08nl
rlqZl0U/8DmufBUHHaBYbuh2S3bUKO2gqSg3Ecv56fMgLpy1lkGH5TVwAA41x/I9eI61rtMjl17M
MUe9/TMKw5E0ecoNFKw3F1T6E7/U3exMuClNZWjTxsHdjDe1mlLpZs/OtGYGwfAu2xuT7RdVAcYj
ktGE9oX6NvY/Dz39vtjvAK+AaANs7WpT+5DI2/1oP9UyJx1D9HL47LEZPuePFaoNUQYY6tsljMk7
4A2fgybyhnLlBJkSRB4C0h5rXZKTvd6gE9qKA39sQtBCmLppcLqGz12VNowW8x1+Jf4ZJ66eE2c1
sb1BrwoqRQF4MoTm3pE885kk64xa6DqT47xVFOy9ZRRTFFEw2Cotd9iUp4gY5xyi0GSMeIc0PsyK
6DNoHmI/rCT0I6BfroMUV05zisT2RmU3YqCTIVbSdXm0QjCugVkh2SaZUC/CFViAX98NHnbloeKm
KeoBhuzROtRelQfv5/tmVgcw1FbmnvlztzzfduWQakd/1bHjF6rTJiRGpEBxM7ni77COPNCBWHuk
xlKHp1NzKMgSPjL6l1xVNghj7mSNUyhVOy25Zd1PIqS3yCJ2lT35+yVgj8FQDxg2jQx3R0x73+8E
bKBelbdawND2aGojaiyu9crSuVRCrgq0xLur4CsdcLH3ImPgKZ6PO7rZHN2+ic4/Yrx47uov8w66
qFIQF1e7djF9E0iJzkY1EdaJ0B64UDntoCbSbfZfvjh9wILz5rMOAFAI5H0F6uPQCb/KqA4RWTJu
TARz259nXAAzTedYK8BBGxszNXCagGlboJr11V92ssRctFIx2KZlgGkCFMtQaKKXOM8pusTsNygI
Qh/Qkf+S8oFeQT36vPWIHFkw4/u1AjpdOwFRrxZQDGaMcnPnk/J0xwFI+W+bDOLQAyCH/LE1MRnL
4CPRWyAklY2pSf/7yAupKa/ZiALVFTfUhAJyhy4bD3a6j0gNF9Rp/Mqy8yUDmi8QmtjtvTb6aHzP
ESDbiuqT61a9cp+8nHanry7Wx52VDx6y7gEweHwR62RqswtNcXLvvsFLwLrkHuuCoJIKN0vG1kc4
/XiS6M86ExBG5dZWoSib5wYFhCdgv3MT4aCZZv1Rp1KqGz13m+I+z31c7swO4PS2BJSObvrruK1R
PNL8DDC68IxBcqR0aJC/qu1JVYf5SSUafNmRqGMRwbVK0P9qU+30NNMP6q1Lx7Gd6g9WsAeq4hgh
mBbbII1B6kGaiz1OKGhbm4VSwHEsI1UUesVw7pZPvaKkJxtOIeTo8WHgmegIjldV/NJZBA3zrhD9
iCXwMqvJOKosfTw2MocK9gGl0wT3uKttRkNQdQtDm4BxbvmipQqXICETbT9nrknfCdRwYdVKTDnX
N90wMwn6p48EkbBCAL61Z/PZcPD2Tx13oeH5STnDosRRiKBCG+wLrfbBp3YLSNQ+NOFxnDvjhLvG
trt7IW5delfFL5bJwjLebomOQbst5+6uKCdcN8yxEs1POsxZonlBK8vcfJ48uux1FoV7aqSXVBrh
4r+ZN1JTGqtz9A8QMVFoOl4dWWpxXDmjPH7RgMjPtkHv4DdI6eLdJNQRMEzpclMfcJ4bG1Gf0t6i
x/zpma9bAoAOFTIbhbeaUYjBCMRlmtUeyJb5JGCQmr2FzVCxfSZeWp50932MpZMhZvFTQUMkx2kl
nEiuwa1JFSVYon1GnUJYzus7JBuYHW6+kXQGnijRv1MjmrIDVUo2mNdIjyorPnMmEMeI746CQziu
6j/5JG+VlttFfocDfI87uhLZ7cYK7DpEBwNTXbx6uZFrvF/fchxxf7g4yE6J3cDT711Iqp152IGX
HHi6LbWEQYUXY+JWnjdaI5xKRfk+Lge9fEEsB2Oc/ZYhqBqkUxzsfOvRv/nnNuYZ/tf3tcQODA74
U77tlutP/tduJYNfjjqyZLOBlqD5kixpW4iGvr2H9WV0yh4UOOJZgNtJr9jYJFQLMf4P3h3KwjMS
gYsh3lyj59EeAWUyelc1QxtCBGYDwWlhlfNHgxdP1vh49PCENq28I1AYatrFTjOtkkVYUKOZbO/u
jZiJgk0a8ysGtpRIvKiWZwzyf0jsWvLco0pMXnJvB6v2y+yh8kzzN8b5EKA6eJ8JVll4MbJ4vC7M
DLdRCQ0qqBqVkpsc/ElwguuSGdPRKpr6ip8edrHbrnfQa27pySqt1jWxnXAy7b9xW82A7eFdYR5N
dwFnHpH5Uj+HY6rC3LFvWACeo1m9156S9Y6eK9YerT3WmJhQk5HtOii27HAm6cdsTAk7zJIZnFQ9
xqXof87opCGX02Fjzx6tYX87F4/PHPhlRQ7msiI53D95QYtIiv4RMSw+oFMgmkvA0TBxjCpT8PNG
9BRnIX/SxYhMSbXAGP5VbQtyV5pZTX7PamkyvhO+okR0AS4SXzgLdSDLpXrqxSexnlT+U4c5SpYB
f3mJAndS8mpKtwN91iovRrV/u1WSozlQV8VMvhfj3XrgessKwYyaUZvXCGCxqouxgPOHzHEOaT/l
gVJHr1eszuKOHTNo5uFF6DpF4k+n3VGxoFm8KDR4+Szgus+9F7huwIxm24C8s0hlAPfjajguEK1V
kmcm+bnO3xjPe84HxjK984us5mNFetcm2FaQ5zZ0xcV+DUZjS4o1V7gegZA8uPTkhB5EpVJBgSmz
9Z2y0Bp4/XyQIMLolErqhIA736v6N3jDq+oe5Ybcb/QHB7prN8dTgbNvvVKXUZyjf6jQweI/Qd73
XLmUyQbWCk6UerNv6cQZdFAE+6K2Y62mQzaoucLt5B/QJZmTMG3jv/sRVLzS5ELnREfJytJZZrfX
y6AYtS4DVgnFHq6JHCJo8/jWTu7FSZX3Cd1AXRsoTY3tnwtu81VcURsE7XlXzzhu4MoPGCyJuQm9
DsaADInsKa2DQlvDPtNWElA/LxP2W1cV0SF2Taa4JpDy3fgXBHqEmQ/+mn/eZEGsHlyXTTcEYlcj
OnU5PYIf/ttSuAuqg79k2RrMa1iFjaikHxuOd8xb5/KGbnrdEOdqngg54j39o0WnheHqc2+UJm6q
ufKbZUVatOomw8eTHwcypMyf2L9mUAKEl3xywninytDt5Rn6PtLbsI59myBz4zfn1A95M1o8DkDm
joYeMHUPIe+4C8N8ZjyseebAVRtVisyrTjAK0q662hi7WsCD+5Pki7XZWsJptg5Qx4ZfsoV7wTEN
OH0V7kh6wgrHPvTD4ZnbYZPVwrDXLAYKFu4bq7z8Xg6W3uZZRx+5AUwNknoOMsRvbHA8tDUEG/6N
HoMJXB2HLIJKz4sK/o4l+8AHZ4W9n3gu+wUxWlVzw+wFeWSSwj3EbOe2EeB8A8xjQtpwaOof1R/M
Jpie3kG+s+HJWkAPEMcH1c70qVReecQc1IaouBo4EJv6vRAED2OHxPJ3CY7OYj1kNHYd0YdK1vRB
AGk0yfcckS50MX2DxJyAvvA3+SwC6M1/rD+awXZ3oFpGzB4g8USCZQZ8Gmg3N71RqlNZckW7Gk1m
iawI5tHhKjyUlGhjyBtljgif3Wx2MMyrx6R8LOtppNidEbAKwQnMIs4+PpguR1u3ROrB8+wk2EZE
o96BU/yG+ylzxvyAjT85B7iw5pQ03ZHn5evCiZrHUKS7MKrtAzY/SH6p43kkqBTj1dpFUJ9Kjj4v
Np66r3MdmhapN2L+GOk/YSRY+bdyfK6ez7jnSwlZnulSqPktHiaRj7TEUXD4fpB94sUxChkJ3bN1
CnBd2rzpeQI3gzNdr+7TD4nPcGkGaSNoZxZkodZ8coacsHTvc/tClLTHa4tThRRTItY7xilh3aox
gEDhidfZj8TXsu6CSGi8gD9+39kIiD59RIGM01v1eBA2gahgzo5rSASc4WrTB5HQTa/7BBpwcfmo
/Uk0wXr1YAg7L6ZwsipuLvznR4lEN9yxi8bsENaxscUj3tZfgA/C0MtK8qhn2cC6J4F6fAOThRNT
9gCWBOb3JtQNWb0LpW0kTtSkiu2+O+FU/f+4+YYv+b1/KfOswQNiCMYwiwoADCtav5PnMPAoBig6
xJi/GiXHF+4+SCTMQIcNkm+E5ybHb/Nie+qhePp9L+M1zjjfcVfXIx9toLb3RtA5A+/yL3XMokNI
gpqPZifK3qWiSeUx7Zs2fac/CoIk1ARy5fjmRAgtxomskTBzRZ0olQOSec8F+/ARm0d+aP+3CAmI
TaiecxZ081N0vDeQXIqMRPGUoPNEKL7UaJu13G8cvxQsSd362pe7DJ6ZC88MKMtWXG7q66gcEDuE
cdT31D9jkgJFQrNs39UpnuwVh2KonNxgW0XPPmluPsK0T4eQwcosFm7/zxSzJ8I9cvjRXh2fAg49
nvd/yc5xVhdLP9CWcL1iM8MgnbY7Bna6QOIOwTYo/pcJOVVZjGqtNTOhq4fc4saiurj2YRjmQ12M
3YLI8VDem34qMrnw1I34zcXj+SzKAkuVDNZ66eTk+0OXOR31Q2YctqbgQq3jOb8wbyFCrRgJctl8
mUMGO0IIcErN8iAswGuyAoESE8tfrREmChGm1yU4ojI5NoOmbjJDVBVYfc6UbXFGTfcKKRU6qBt8
RpMqZM1BwKcVnxuuaiPK1OOjUOpKAp05H/I4msfbp6FprYLWZ31yNkrvTnAuNs0uq7NVFObZXi6+
28ZCq0eK/M+8UTJo/FPiY1F2A9LYo2+T5F5rJ+Z+eN5hrKu0TXnEBoBeuynYXYgQPA1CdKLGqsJh
662LNUBVPNOzfGRDYlEj1mzXNg+VflcCxL0lnTFeGgNki6m0AZLTiSNiqvTc+3aV1ri98fq1QAAt
8N8h13K8FlhGyVla+oeVu77ehfH9IjF/5hyBfbU4spYL2s5V4oFZQqWfo0gkZnsB4VG6cuK3SKGp
Oh8Lq4Um0BKqoW/myAk6JGl4qLEteUXcvC8YyxrzoxZX3vmsSDbVQQNaENxbwhk9fXx+KYUz29S2
HlKPRc522CiKkLxu5OKgftg5p+uaskqzkJF0apne7UhgLXmbbm47yv5nLIQEsFSozx+xIJ184Em4
RdGmErsBPx3iGzK+aLgh3E8b/5F+0AWqsR+OBS/sPTgU7odJXvugZKgtDYA0G8JFDKYDSvooX0NB
JCPlKOu0E6Z/wGYHA2MVugkzrV/KLrGU/RvWFJf6CM93DRrvvXmFb241KXvMx2PAK34eI2U+MMPM
OzfSpVRHzSAX4j1YbnuVzubL7NckAk2RyR2RW7Up8eCxnnnHOryrbLc7XAohnzjCJS8XDNi3j90k
enkLff2NTBzYdti0/dxmF9ONNIaMEww7M3+6T/jsb5l7XY3VG2dnJLd8OQjCm6h8rUU0t7CIRkU+
4GDSWPmQ7c1QXz2Q9C2i4C6r60FtynbGddfJL1uqdPXb54GDgVYC9Tta1pMaZKXoR2fkIlbK2iz1
abMWXnR3U5NHdQIUyqwO2Gt7hnX0Rsx5iEh72Tu2g7cifAEoPIp5jBwYcr6U9DuhiWzP/WQRPlM3
U2FEX+ooZpXHsA0A9mbuPyVB4uNoHFN3iKrpQnj2HfX8mQdDe5v3oMt1LIzszFOfHgsPuLC+Ft6+
Gj4Ljkq1plghLRIAX5YaZxAfxOJn+WCXcDiKYl00pbw0xs7bJiQl+0dQrkIahnUiR0X9NtCVj1E0
VZnN9uIRCDNFIQ+4Lzzrmcik8jIS1hPUirbZuxuct8YLpzfnR1KlwHf5/+a1Wgtoo4MSSLZrqkUf
odCkLnlBgCI4ZzQxk9Ipj3llCu9SCw7KytjDvscjMpGAmt3L5JMZI+ADydzBtTpQt3MonMEPT3vR
ER8y/421A8Zz+orppZevW+6AbPahpU+IYKg8hng0uipsr56GhuqHQSDQgzgnFbKl+5YHteL46yRo
8TpdNYxno4DzcBSduzBw44XgOXy0HKK69CDIqwMwgOOXWsK/tnBQhw/Z7DTGeZlcLbQBvHU/a8So
HfWlNbRA7YEkVZ9v7SNfQ/haPmmw4BuVQDggPR2IDcUaARsCLDerSu2k44jV4S1Xaz4UVRt374W3
fCmhfdWUCojQxDwPivDrG32IBIgRlP3P26W4loEfp5nrnMbOzpMlRHh3043ZKIUXyniQD7VyIUpS
/2F/56ZmOZvOEMHsuS14P+tLXURi/tvo+gpDC996Kp9IUaNgdNZoDZ27vdPCF3QW59kRDsbaeZCI
3m3lmcV9g4lP8I435QpOSJ8VClNliRT7Gpyd7pt4V7qfjzWR7YDY6pDnW2Ebxi94PLzbC2Pl28C9
BO1b/t0GZWL9CLjF8U1wxx/ZRN3b0f1TI+EbWo+nCi7LesqwhUHnXkKXfs38Yclqd0WxOClJv135
CAkAtr+roohZfu1L6zAQKklYCHWo4IygR+P+Gfp3oAnyUeOsk+2B7o6i6uWqb1IxuVi1vuhstGeQ
cMs5wYW71YSshO+WmjOQVHU6L9UL5kX2Ge+KAvXTWvm8T1jynKmXyWI54ux9ZKebSPqjyQXeyQNL
fBKBTKpEtQZn7q5cD1YFMEMdn6cw06h3iatFNrka6ceiC7RDRoycPGkMgSn4xsZyZcRgXDEjHKEn
Os/etlaVkSR+vv2CQysdrSqxxATnPGJpqFWbLcbyq8JsFQCPnfMi0OkAVBFbHgoZY4fq6EITBr/e
Rw+RbX9ETnchqbSkPops/tw6sEdDiMbxkJ9xRdpi8ZhZqDDdg1ltemLgSRczGu1NUMEOrw3KqmIO
CZaYs3SmBV+H8HX9SOb9K5t1u24fHVlldAYJW/ZQ2mMixFnDrFKPy/Ni29LU/9GW4rbi7JEfNovS
wccgLCOP25s6D8ZCcssxxuGumnrekLLgvpZXfUDWIYGpaxsHR1Qx9/l42n3zbN9Zy8Q6pf2C8V+g
fuqpUuSS36JZnTZeREj30409hBqn7Y9wBfLdt1Bnbklb1fqQhvfKyTxK+50p3m/UYJVfU9rEv+7c
AJoBwsevHArH3npgPBpCVmNrZckPbnbflY/gtT3p0biTmezmmDveVGWXUKOYYYGiXzLU3CCMXtef
Tq43KZ30x/NGaf5VoFhEHyIQNcaxMzwqgq8MZoNNVNoQvtDgdJUtetYyDyk+5C9NpZ5pyGdHcDoV
CCwDoR/FTYl/WCRnXuemU7sFwZN0zgo/3cexI3jM/DgHS5qiG//+tUbPWZAtDWp1Vou+4IjiqCOL
rFi7I5WLb6CC0foQH/FYBiYGp2/w/dmwMFsGaZh3844q3jimtPyLUWWS3wmCi3hpW/yzeJZwp5Wy
i7+gbiXxa86raZ+HhAbWZo+eHFDivqHIzgMLrkF0redrGfROXigS6RARsLuyNPR/+BaXx9wI0GZd
woCKTbA8gw5GkqJ/NFzwZQjmj3M2OmpCmv4c3szUyfS1HT35rQ7ZOT7C7r0VqFaUb/DGw2GcedfS
n9/Y47RCwmN4IfkahfqjxXK3jal9qOtxkitTJJmuegth3DRNZpNl8QyaMr6AnUk7u9WegvBEEZrj
N+m71oosKOt7iLBC9/tKB4uommuE+4xp7SBQgcD3gHSN4Bi4mnewFNNbPkO19BbkEYAXIktIhKJ2
7RLTsbwGqYe8j0aFEu4ANr88MP21Nl7gjwxCwj8eYvhjQBT6xOx5R/XYPs7eno5TDJU+uxTbRhNy
7lFS93YvwV8o2YVjoHdZrZxfT29dwS8YOXntXyFcaxtx0EHnRgP5HyEcFrW2CmzYGNjvkuwvMJtb
Jry7PNvSyKSzdgciYI0exgn7QS3BT/zqTlZ8ak+rVaUUqJ5fix9y5jHbjRAFP2gLI2e5n+c2xvA9
6pNzoIEOml+b7t2u8AFKiwkAdiFimH/LK4JGU7c3uArt43lPjrkr55/NRmLbaJJ8dstOHiJyvVQr
Xaqeb5PMH4+HK0ew9rfpXh3aMCmiPH6yco8CsjmHYVqE18d8roQSr/BSL2JaJzKn0LqgAYvUH1+7
yRMFRn+vsjM9zc6qoWRR8ymW5w9FNgQ4002WPxwpI/GLJZ361ssYQcK0BXrPLAo8GetG+TOUtLLq
000nZxOTlplVRW3+HoDtlFyBDFz7y7QGwOR26oyzsMIiWJdI9TuPJv5eVAfQV63wpL1tBnlj012o
t+dDQp7WN6tXf6Gf9wkKQEbWsGN5ZhYjv6OY4RTdNKU25PGY9yaHXGwkMPH8iK/CP1LId+D9qFcB
FlbdwOkmRs/zaZ8/+z83FOWW30IFjFykVTAt9HcXk+FG2NxFL96vYEX3u0k3BqnE2gzEWRFeuT+4
YQg8RAMnm7cOxGV7pODV3wId/YhvgpyFy8LHsDsHqndnKvaWGyAk5jZlcg8qMlHWb5wmh4eBK3Z8
AlzoGqA1xZIIHOryFfnR6RHtnHcNMf00k4pi/Y/NI00RlAAFRIVkJP52ftAvv1ACStQR82vcC57b
9WRFV+8ZZjDuXDMQyCwb2GU5o5NoPtp0rcqAR9WOczJzMz0DOG2orlg4yz0zxzWmMy3xhCk8Fvva
aguOZ8KUMcP7226A+MWKvWQ2Afx1XWMppv035MoZ9BoHluYP7Yp4CjEUSI10te6zVxWXD2QYBlSK
g9h2jUzfJkEXDtqpF1F3/+pUMwiM4v96kysN1JX+ztKKtOdxgpxSSQZ0RoBcvNGcIhCwvdjJMYll
WGhZe6/ZGqhNwkd454akB/4/MlffjOGKYy+d2g6PzM3b3WxZQ56WcYafa+RzWdXrZRn3VUN5wIpv
2E9MFAF3O8BqRw8MdOv2dcVWJE65HecM+bDSirKhTHTvaKgV/lFBe/zJjGtbEjXEKTclgym1JIGO
eveebhpWBpiUVZLSzcTSYA4XN7vLUJfcdzMoCignye89OvrfIPqBRUH3/UlSumU/BahTd1gy90Ky
Zg+hw8NHhmgznhob8iF4inYfgHqftyrJF+d6uiFfRRs39XR1244pHuwr41aaKdkcd8xTXEGsTQlz
ip1yTUNZW53t8anFV9XBcPSk7nKZ3vESWB3aE4qTUP4hHNKjG4QxRwQo221lsEE+Jj7SehxqgXO1
oUj8azM4M1nUXIEYr5+KU/mnxn/ZXaG4oXNNdKrpQgXmtzFm3kKvlTP1alrNAoRpPzN1GOQkYtNc
8FhlYCtxCM15dGk7jCZUVa4O+ZT1E/sOQAV0dDRjTjVXES/S9+URX87I61b4NMThrUvwUtYQnR6D
Fdm9EZ5zE5iKp7OzD2R0x57ubOkm0BJxr2u3wWtLIP4qXz1V1VAgFPF3t/Ic95+xXmyMT0tIz2QR
3L6ESAcan4nNMHiAcCBNE2PLWPGlbLpxAQkKUv5WSqId/4FEtinuqc3bKOLU8py4tCNMgtNNppKr
soHIua8ApCPIa7FneoUziDsevwnVfXZQtP/MleZGweiugwwa72yofDHacTzlaDnhRoloMmNeIfyq
jeKTXD1Sf11dTy0KVCbjE5vg+1JTAEJv8LBxkB0iASiH5g5blSVqz0a5LRDGBojTSaecL8A/YPmx
c7GpKdqE1WJdxaSYdneGw3PguNIkDgkqNNgfVMFHnU37YzCh2lWIj7ovBbPq/AIIHiaK7CCqLin4
+arWRNt7XrhVEAnIjJhxHwDDulUs3n9f7WrM3dCEgoAB/0+Q8uI86JtRoEcSZS1cL33OcoL/MoWK
e1sCIiiYYabEapGSufrTAGOgxq7qA4XAbxDZzZmRWFX/mPpLnv50RgqzMxQXzDPfNSBUjpdOV7zj
p0uqKwWTTmcNOXDpC/XCOKxsTH/tfn5AKw7NrzcUjDptqEQ6NNm18o/CfgrkT9hcGO9QJuENoCA+
DlzX1g3o01iTrEoutZormCSENmypsQ6PE1kIY5ZcVKO4i7odNQWUtzCWoUwIviqCYHj/VynA3e14
0mpRtoMWm6Ai9mWCNazX9MPccMP7u4525N5r/RCj+uNiYWwH7+TL+FqGhFcJz1FD5IP/W//DUW51
iZwF38c3So4DMIkG9IRg9ezvCjNsdZDK+QYYrxQdxXfYhYEGjL85Slpr706OnWAdfNRwXCcnbuMs
pJH5YFrre7gCGv/Wxgjwfxgqn7EKHjNtkLdPlrxYt/qhol+pzSU+qw1Vk2iDU1qchwVERvs8Tr38
MDIrYgwp0cZf8P3AD7u8ts8a1dPyGttE4JWGNHFAbdtybBWK5fBDup13xO0jlRvfwrwEwljXHLlx
YRD/FDmQgqrcVpZlUvd+oYLzt8Gp+cjcta5NsM1ojD8MGFeX1NNPn3lITIHTAdzEQ1Sj92MLm+tc
6BWnpqZF7jUKm1BxUZxjt1hJoJOivp6hkrDt+Xe8u+e2FW6XdA5MbDWkN4KQSWr043K4CJjgUZgY
mvza5l/CRgT92pr5+bz2sInlkVMAs9nBxS8XeKZH1VMN304gSFp/GThPlFoj0bjAEPhiIIE3uqLa
nk8OIo/TLz0Ui5IqM0d8AMUmOXqITfvUue5QG28evuEqrP2poNqINOL05c3Jddi6ddnTde2eN9yy
rND/r+xQKBOc48QmBRLi8sXaLrnwQj41HOmLHR0qBJVF/8BOHCDcS9p9bsMsBiKViqDZg0IiC8bP
ytOhCd8AR9Fu1BQI5Ue7RqPD8gXICcwfB8RogrQakyFQABNlejT4Ql49n0p+GLTYFwKnjrAloMen
NcNfinrCEkcw8awGomsQ5wiIJ6cTTIgNpJAr24KRd9FmLSPi3lTEebGZKVE6LQvToTyJA1O9UPQ/
mOfheWf6885NWzMlvnLl0XkXy+Jx5TREp/XK/swYdeCioPvGA2kX+JvQjyNb3AqxjuO6dIKOVXgv
/xFEAgHpC/2+F9H7NJWx9BtJqf6MWfXzzUWNiJcVic1o3U4pLKdTO1v0FbyJUWgDkJAtCnZBtYgz
MeZ3IPiElODKGA5+iaiipyM6s2yGcQsgLN7ywBWN2+sigFdR4mFYjbNx/X0pM2IGI/X56grQEuO+
Du/Rpi76TDPbhZgzCOVy3PX5Jua9d4sYN9vXRYsw8d7lzGYVidltMxc7bRfCFwNmjMabMNaahIsy
z+jb/RItkuJRBXkwTOPIMx8xHx5O95CAH0tF6rw3UPPgVsWgjNfTCEKqevGqtGBBR46Hbf+7oleI
0FMTlrQeUFHOq17PMr7sy/IHCxgLJO8Y0Ln+JL0ezc92HaNpaWCKpK6AjFxFp5ZFqYJecX1WZwYL
LgrtSTWdD1RXqxsOneHOD35hQZ4SSF8TFvP7t/yuneIKfxBmo/g89fHo2mywr2+X/RaKQ0noyE1h
ppNQ70dCeMrq73WQI1TktT46xMiy+UoODCUL4BwClFgXw7A5BcRa7Z9IhfRGCzoL7QdTfeAP6+9c
DlhMfqUZZlvlIO6rrAndW5LP7lygFWKuNv+ZWYympfDHsa02+/VBF8DzJv0yJv2aEGis3t2BFSfB
196/wdqGDOOBRD55RWdruOY1vb8Z7+wYTpghHD2r952lW/thvRTvsZhsXI6waKHcRBS2TOPqdDHm
7baZfaSGRfht3Z8hOXBPcLmD5qMCLwBDnUJdgtQXL2V6JYmYIBsU54v1ltcux8mOy8hmyp/vicAR
8rLmRmozNd8XsExxrr+Acf/duYhXOGOXp4EFmCiV48zvkhKqrITPeU6Ni0ha1bYKLMTz3uZBgsFO
yXEuVKmV1bZZ080u3zlLznkFrYZuNINYNwoty1/Bc6TPXfDFCI7gJwxg3Ad1V5pJD0oO/fIgrnI8
KRscHitcruwGdVA1H2WGVNRBANUtUtu0WkjS0hHR63tiWSuqS2ua9MBcruSDbZmPC3h9WnKQoYcP
pAtdT61HB9XOAme62lsqcL3nAZ5w2cUrPZooXdv+YLWuxHZ+BrmaTLo+zH/EiwvKJZ9uvYi3ttcW
uixQnWWbEjCkUe+ag6cQqW1xx97x/jET/yUtip4ty8cdPyenFctjKcsl0nun3NFUbY9aKsbmbQrw
XzcxEg9cqa6QUZp3mro1uwOF98CArHy89KJ9mVarwXIWXWFTQnwVGNvC9CY3YyIyTF4IeC77LZWJ
xcpZNVi9N6pdayrLdJhxNQo9e6H/uTUd4my9hESMPGZXv3ccehS6YP1k4wRPbSddfQd6WN9i0T0W
0fMUjbvhNEwm+uNDw8uoupQcsyXu0W+E3MigoMlP7KQKKfqvVbdtdJBRS8VhQd0y3rAYAH6Ilru0
KdYiRpsBk6mELMtaSmmQQp/FFanZPbpfCQg2fgGNFyW3vXWvYX+p+Pv4tVrihGT+Vj4AilQfFq0D
OiVvfM3h5MPhr3Die0+vsG/mYYi2KCde85iTqx6wmWMq9wSvDsZT1MWwZMCV3kD6dzbbd23UA+cY
udoE0IDSQYNU22J4ET5C31kqlcI3P7KaPR9n9sl6OvoBCT5YW13tw+e+Lrdvt1zvqDqp+UfPNIud
NTROnIp/ErkGb8eIFLHBwtGOqNajDojTFMfMEh50u+pi6lw2QuNXMMQt6Gd3nM3kMwhU4m0g3ADr
L4TynP8M2Rm1dUHDgwdRz6B3NrCRryp7s5gYDpg3Mby/tuVmJlGkNyZ6pcWOglQaq9I8BMKUIrCL
rkEBGc8ci7YNMUT9cPS/334QrJW14m2xIGNkhV3uJmsmrwgKD9bcfKSFtBzW3ctSsm1H1g2KPJKH
KXX1OVcaqOCM/1PUSmPx6qIO83+pz7uFT0iXlkysyFPEM9WqZWamA1LBT7rre7HTRekRdYo72S7h
/ZKIJXV+2izH2jv2zGxUqe0K5IjmB+pkQWzm8LprfuMVNyfkWb2GlUF+aAqFN/tjyHO4ixGGFcdo
hhCtBJhdTTCKjQc2JZ3as/aqLhkvFC5m/LvCvZN1aL2SiQoancsJ68AcAtXn68QfqaNvbLsOnJNR
HUGrOKwT8hZQ0nTrtmWHk5Y1bYx6s5tbpwp6UAwnemqVxBzy2zFDuGvHtR7hbgWEI1m2XFi21ZUo
JNoRpiNP6GyR9Hx/d4mYqn/KbKw+wDbZvIHSDYJj/S1OHVVmmp8ngBsGCkWAJxwsQEs85t1wiiMn
ZlL/Xyy7cmb8dPp40+QM8vC543+dENAxiiLkY8/WSEcYqAhPHKhPyPR7cvP5MnOE75ei6BpdrvpD
bVpnjwIxDlFTNiMOVkXFcIYBXC1sColCC/y/FGUh1VGajkcC4vfEJP2/K7L4VwPQqvoKSvEIXXXT
nudaZ+SNpSxAEsCQbw8oEmVNZ/bAftUr5C28aXiPECZGeHAbnvBryI/mP2ZHxxRUMuVGN6vCj3TB
n7LREjSjRfZ7bmxG9ONuJEdrTl41CcG153LTTbTb7iahJqLxPh8DHVan/2r1MXluAwTvu3uYrhQF
bZY2kayCyG0ccecAh7Y+1p3EwD9nYLBJPM+kch3m479Cp6Gx7Zu18hKY0yQeAEMCCKZSY/PYgZEK
SWdYmBkGJN1MrGOyDtshYxgnziaESy2GzFYZt7LOQ70c1hgpHDGmnC7NTFr2EusNhBoqnDZCfz9o
nQZHycolYeSQ2Y0PsOw9+a6c/fSdd5aOjIfx3cW89UKi8xBTOJgaiNCqtxuhgBBWAlBcb4gdIABT
T9hpkeAIvhYKBkSHab8UaESQDqp4ix6tzekLsvc8ZW4vDitCrW57ci5bfmDXiZ0+u+vXUY9fy0YV
rfbXixPsAfUFuZAlpyiIrVwQzcW4oRCl8nO7Wi4l1VhFcl7zdZ18Z4GBS54zi5AR+6tuMRpwluWE
3A9r8oLN8IOl2jtI5Njr1Drk19x8C/j1Ry/1fKpjcHfXgBh/Biq1n8cCDdoqPY7h+nHwRI1I4vR4
RGd2BRRikt4su3BFRQJHLJFJYLANo4f9lYjFcQbEXWMiwqKpIaiTvt7xMskC3PD4vrT0lL+TNtFG
HLfoMb6fudA/ZuFWcINrfJX0kax0/Ov1GJgS6g70SqLGgFEdo8YmUeQaupWs5p7a+mGUFJllO0fu
FiB9rsGmsJNSxDNVkOumOmuC/gWixY+D7W7UObstFX/tq3Vpyxdn9+sRPgW6W6tiIS4E0VFH/Pi0
znT9JQInVwYELOa3iAf5NUNluJhELdduYevFewTpUnF2ZTC4udgc4yLkANDcwKf2kesD5HnKD46/
MbUAyWmPr03LqIEcgU8o9Z6Rz409MPamT5ZIQ+E5yb3az/CnCVS0r+2XojT2LGVzxPaFCd+GQHFO
cA0eaWVubHD4IjeCnvcOrdAjTDSIUdWxgnPTBrPfH8fOjUMPUZxc4GQQUy8LTaHuUln24sTLGf2Y
pzibcS20ZKbuWfPBnOTyhbOHToo+IwPN+D1h494yW9lX9g7RwHKTpyhzVvPFBikyyPtP/h6CT46j
Ax87BcDtGA+oPcx9apuwlNRrsynvXngWTXsnHH9lFvfKg14JrmfTFqXSpVT1Jx0fzOOac9mug7QS
Sr6r2aEotdnpii6wT2cnXwSdQ8JoMGS23wUv1fHZmIUI+2geTO55CtXH6hCOgpbXFzwfyioQX7E8
onXoPHZVzysS26rkNooiOxrM1oQAflIZ7MdX3EvC3WQZHfqaUusuNeqeeOEf5rNH5kUaz9T92i9O
v+R2ADJoLd1oBubRZHZhTqqtwM0sgM8tYOnuFfnhL4z5xy9kSgZzciKrHZ2HifIKAd0zO2TZTcxE
7sV2pgiIK78jBulMs1ij76zgnErMKphqqYAPzZpxPfuBNXRKpICNRKLHESJubAKRLh/xQhdrPjZH
WXX3k2yy9jcDdVb1o1yXW3doTAsheJ6M6ilSyItKi575j4CA/z4TJ020xhRuBSDwXr3WuJ0kY2vk
LbnouVGVKtljfYovp1790N/sOAGTA75J2L5hN+2UixfCW2rdc+cwpFvlbH64sxC3Ne/WiBIZACMR
/ryqykp+0/z+t3pAUEAy7tXaLafT3S5IEIUJc+LiU3V4iGKEL4WSeIe/UYLl5CFtbSQrG0bzOz1V
sohW0okbTC4C/qE4z9kyHspaZ2CeRnP6NtYg7DKPvKh1uWni9MufHqtCHPKD7yei9UU2m5LtbbRS
sZpfaULZLVLpMXjGztLPXVaCQeP5d0LXcuFrrxdwzt9IkamIF+Us+07dr8Ga+28/hWk/2IScWUfM
uvxnRe9R8Ud6OUIq3mmBB6f3WiVwT4ocMpz05ygEkG4/GPTnU3Lt0D0HzwPLir5rP0I46NFbpxvt
tfxFAtpOIiL3uqGhk/romqDKlIh8pD4MycJCIvPZKjjGzcluNgqHrJbt8/YS5qEn12h6ksOFkISY
ga/JSho59MY2TBaiR6m+cWlvynEsWQ4AD+DJT/DzSa81u+mQ2+SkcsvoELsQYxJ6WCJCGyqlQwxf
P8DiSFF4VAz8JbCDSNqeHLnxRhGIncIxDzGRr8q5uIxFLIFaOI8P6Wy/PaYnnJuwLTCWY0D1R/l8
/YDdAQEpL1zEQwSkylnwDVNFXYFS82mUAU3KHFhr/AsFZCbkXscZYE479N+eDtnLVzaekTvg7zPG
E/34OWWOokFFeH56l8OngdHx3kA4t/Kgd/lR8zSmJON38nH9XXSsjqW7Dlflj+FC9wV2qjmxjQ8V
UBbKrxsiWqOPeseW2Y3Aqny6hP+EdhXRo52JIKOIA6+gW2Ifa2XWRYs3yy9derXe2QZUpCdX1DLS
KZow0nkbxiwJdz1lw3PDDrQb6VYFcn9+uArT45Rf16+YF8OfbLvYHgRX/2vuDWWDbfruvBZSyh/g
cOLyei53qMzIrtFJNKrGsiNc8tLSkyGQb8qv6jr7zaAZesvaQlb4bbFmcECq+gJ19J+0CXOtv+mY
Ww08tAdXjHPt50Y40pqaeef+Wv6qWLasE6pqw5EImYzEujycCNJFjBNe3oZgLC3uM7hKpaz6fc5q
LtZCQh0K71mzsxtm9Yp6MHYsc81sff/OZBWOcbAmYjzFJ2G1AS3TJVKF3QuwSNyAmTKO0uVusMEg
OvJM7WPecjPhMAMWNlFHojCP/DWKDrBAbcEL6RgW8CFxGf72lvXtgkvnJkAfebzvEmGxGAe3hDZP
2NezoEke7jJkSIv4teeLVq9U9KbOmPZ65U78JJ8qJtRm013bXUNrqzllIwWU4JU+muffLdCbmHzH
UC0mxU7YfqQe7kcX6v+1ZNAgVvfNaApKBDOUSjO9Lqbt+1ANFmMqYYo7kJu53Nwvt9lGBmeetflS
7MgdK+n5+U1lTDJE0lPPVoJDggw1c2H97sb6kbaEDCtyt5JTiqTh0/Yy1TNPUL2R6EebMpWyOCas
3Y1+7wU9JNqD40M6fGtAUrGNkrxpIZHVy1XqIintVZXVIwMDZ4RRm/iKleWOPZqwPL7hxym3Qdvr
5SUZtNSkkcLD42WD/LRDQckuK9rl1pgqnf4Vneqj/HK1DuhTmh6yzCutxTk5GldOC0NZSFTNfrCg
IH8RcOODpuXh24o7WG9PKL1iksXKPcVKV4G/Y2gFnqfG5j+qzEeT+RZKBtFviS847o5CrSV0loNb
sJGKOoMqWXwJgn3KdMgPgBLIyutRrKlvaiOSvLyaUtc+Fsup7DTggc2DBq63sg/O45VotcIpSN/g
rPKYcf5OdckHIaxM+s4yDH+bFI1cxFn5GYs6X4C8JLvXQ88eq+sDwXpZFHd3/hO51R8fmsDrf0K9
d7I0bRIudFKX1dK7Ujs9TVEyvD0WR1ug5Xci2ZjBpIS8HrOQAZ8rhJOu2l9Qy2VYjz2cIkFSvd7n
S2LTAP0MYU28Bp937b/7di985ksU54MjxtIevgsjpM0+NXxDsaoIqZOsBpmruX6TEcvlBspLJdDx
bMiTTwwmsuWtR3f1b4Ks26pdCe93DpQAxsPGbCiDvDb0FKJHYtLiJmlK5oukSfpcUsYFg324t0/u
x82/v0M0LfZ/7iVJiASZ8n2Kv8AUeX9yy12mWqZLWJTJtDafjRIm6q5dYtgm4gvWnAFSXavpTrMT
MHN7PFHyt9BoAjUZpqcdA2QtMiDGiA/PRFWRTSDfhVxxmb5+gsqYzPGedU1WLClpLzi1LSX6LFG6
icK85HnqzJXDkhedF0WZ5mdalDVbPE1UFd068OXkq/QZC+vtRxTqcTeNfUo5GYQ4K08Akpfgq8RF
epezqr5GRnPDeMTZzRaRQwiUSi9N2Th5HHPJyrN89728WNjSVdXCd7+5JWIbyyFMyHlcYvxNjnNe
ayzArsdPEeEE2cswGHbLRVgHmNGrVTJhiEOaCC8Ovt17IeRpO4WZU3lZyqFfo0ZU6bfntYrnQTC/
kQ4p+W9TJCasmUZ/8/j5VlfYQB6799bDRl4sFpddwls/MiqWo6KX3bs9K5GE3w/8eSbfFGM4eIbU
0EmOTKLLpKAzdmqQXgoL5+VBAsSRFNrbSFGcGiaKmrZbAHqJCf+9NpCNpkN9qgXyTII3g+sMaxqF
wIbyTs647i4IjVPAFkQb2AGe1P09ivkZD76sf0pI0kCzTJD2duo9w0y9qyd4cqVypIydrXaqunqN
tapLRg5zFd/WVCp4aAILLtiawaEwmaHWwftNL+eLwHIkC5L86lEnL0QAC+H01FwetrHW24wuJrKw
vLmGuilA9LzqBJYOtoK+hO3lzpCIbncQugVDW+HVnDv2LXcAP9xjw4TmV5Bib08fTlm1cOQrf/AI
Ap9H9LW25rcyIb2Q37CbWo65raph0n0qB4DePnhOJ5hsa0XdsxYTuDtN2+X5DVMTlhfMuozE9lm4
mC0VuxuzObFT1cbTQWwohUvmwHwFhFxnXYr2KQN1QDxzJ4gaU7MMPAQx0M0TWsR8IIMfePPeAAOO
XPfJCGM93Y62HO9bGr/7hxOHFLb1mIcIVLylsEGEu9qd2yDMC/u+CrBdu1bXM6n+L+anbONFpVqw
DLJ6FqVtyHVq1dj4sHc+P7/DAMVu8m54u2nONbsHNffWKYeMTIQFokOakGk3qKjDyK9mS2toZEXX
+IeoS2KaD7+TVCRSUmyo8L48whwZhWUq78jEMVH+ikirONG5EGfvg6Luj514EF8hsZHfsvka5sgp
sGLjzBgVk0OQqvtSailJvlaRIjBp2ZtUs7l/YzI2WJqXa7pBh0PipOgb3rFhbx96SLMRWMhfeMcv
TrlkE7fUOpUW8tZVRngdEFTXA1wAhwM78W6RE9g4owwMz3qcetTV6Dz7jXg3FsAX7NiTy2mpgQ41
VikzQQwFNADGq7AGTlFedjyFm2Ad11D1RvRdyJTLXISwgMaC8EViVkGjUJOStM24r7cebgC4NlMx
3IV7Qp00TI0ttpFI6B4bjvrDCEppShqNm+RK4qVnB0r0Qy0irWhR2BX0R7TWujKL6tQ4gqDliCHC
MMIJr2oPn9yXvUpviWbYzRa/SaY/hC9bozAyMP1uPKze9lXzdRZsHnxL8wRTAXaV4fbTdWZdl4DB
burBKrxVN7VjuZgvfZISN4MzLPfM7KFFe8bYVMVsDlMNsaj0/6/jUndkmaJoQtMAe86C7a8AxFeW
Zc5XTOOqRLB56Y0F1Z/pD/LYkOEYB7NVrgToNVPPzTvQhGB00LEqwOwxKYwyBWWZUiznVFTlP3Fr
MCvqNgJ9ksihjOz7Ah5j4FjsEc+3s3x5Plv6FK8kvoKnl94nBqWDZFQTs0HA9hMOqbSiQOdTJsJu
I8V6nLV5Jfno8ymviOOWkKC+MW9c9JwuXzaPfsWznAKIEfTJnHl/xM1iScNBN0On44CCd543ohbQ
28GJ3HD5fwczxmr8obgmIRhY1CrMotGa9PBTb1z0VFKKKSgMY77rtFPefSI3Dn05AT8S91r+fG3Y
0/3NqvJzNUF1ykURLZKaBXiHzx20PbpnDPCW7mly7hZS1dqwN+xsuHeQqH4SOk1lKec+G8bvMfxc
Fv6NkLfNyo03R4tZO0vyc/3dwRXV9+2gop1t1ueHs6r0RosgeYlYR2dKbd+LogXyiUmiUISCOuAH
TdkCetG8jnO7Tz3zbU/La3lBWnV6cgNjeHLVR4gJARA/HjxXtpdKPccA80LHamV79sMWqCI3KdQZ
ov/t52XAyq7n3ORGft5XXSu3iLrpsBB819J00M9XS2uPHh4ebNVPU1U5Fq6xFlmRyeHAmC/kRPC+
4sKzEPqWJ+WNOSxJp5DUWgQjDCjiAD6fpw2ltlDFC0venr8E4HLV/327r4B/fuRlQ6xQ238tUKch
67/7JFuFaI/HyrmPkC1ENl3jDCZVbJu8ZfbxxzCXo/DeGxwDNSlU5cu1m0sWhvvORtk2HNEkwFqa
SYhpj/GJ30GCLUpzTEkjSeDf8AdOBBvZ7sbtMwxvCdf1nrbc2Y+R0rEp8xM3fn2YC5wwSVUeNRnJ
paLzwOqbL2QvF8jmijvSvV+Mlv4u5W77tmgs5qKPx30CDp0+nUxvXRMKl6JSmijz3PEW6P7PEWQc
zWe/O7vjNOEHvsogH3qdGJcbWlPxf89e8sgliQshiH3sbeZqWX5/79wXAxhxZ//U2wk9Plu5WFyN
Nd6RNPz1f9sPT0Kq+pvuznMy/ya3emd9dm20Bga+qnAVGb5iP04MDGYqW9egtbLrehfzaFehV6ov
we9aaoJj75fKVQNE1XB+gLed36wU8TIfaVbVRFEHTOMpUSxIJa2QO0yaCPKsOuX+efy5IC2AcVC0
pQnp4x5lT4KNfSTnQJRStJGlc1keISu3zoFyo7D4ciUh+er+qkZbIYzSVEKSGnUvNcDjMW0q0sMJ
sG4BZCxa8nVOE87StAUFUC/VzT7/w2GRwAvGfhjjZIVtgdW3QplJVs3alDVWIDg99ZwYjoDkpghl
mpF2/Z+l5j1pD1y8Os1OFt3fD0VP+nDdDTHpS4UqfZCSZpZuUWyEexSeUqOkfTRyjNzp6GJ53Jc0
jYVM5jr9Uyx1Y1LrfDfcO8K8dN/nl23ZReRP0diGCFXeRnPw4/8gyOMcIJsVCV3CL2OYV31RYQCb
7sCbvgSOovNVQjlgIkQYKpoUFR0LEkGtwsA86nYq8Yh/DZVxRgs7xtyHxeFXFvVtihEPcYidGmX6
g/JhPDRirWV4JSWUrxyNLHVdNRej0F6CTGdQygkRyEHvwADhSxIPiExZZ3ILp6EvrWclh9Adu85v
+TNlMpZAzYva7HUpVgQvDvs2Y7RtjqksBQAGj8MpcPOpsrC1SF2VhB14aRbq4XPg25aMoomxx1Nd
7QK411o7AwpE5PwHpfOU14HboKdKvjE4KoVNouRDT+nD1XFLjFzZ9XNn3bmFW0ZEoc8meqo3PeNm
C4/xtBh/H8zinkGfs+zyL6BuKKeLlivK9MpHmTdE9pIqgBn9QosIdDEXZj/ZNpL0Py4Soyk1gVUg
8BfViPyTT3Uo4OIdOrqwCb9FnJos1cFL+mX4EMhOVE9V8p45GCGez7rzsVxN9U2sSvDVUfCQVVOH
oY8IRn5JFC6OBgdYMozoBY/dqmOkDVN8f3Wwl6weGqgTP9Aeb+kNNuGtMikNHsGvs5A/F9XkWvBD
526RkztHvGOIWNFYRQr7EePAJ9DMSBgWMj/9CCz7BBWzxWPAt1qnt1BEmqhE841pTFfbBzZqsyiL
87RQH4Zmm5FPCk515y7jpadEjnXKDEo8XrERWlqMkZzQsBMa7tPCMZSshDgsdqQ8Gu5g4ANzKzt5
k3FXMYB3reb/EKPYP/B6fvXvCzU+cBVIHCfvQ7ZmYzMDDqnrKNKMiPmD6wZ6mW8Soo89R6O2YL2v
jBv+xNlI1bSqA0/P2EchOZaBuHIzrJs2IkeruLT3BReS2P02VrmUJkUhTKVAxy78kvvJ1xdOvhp9
6LIFufnFhTfSpMXz0pHdfMPXWo0ooAa3HwBn/dHwV1aTOmX87jT3+3Mq5kscP/A0PQCs5DZYgiNZ
qhvCowgLDP8ScesISYSi3nhrOiaxylJmaRmh0VqeaGZ3iUuCRlHcrYBVCRTp/7lgtmQTdZvDBz33
rY/3asdPltcMxBU0NdN1chQpBjxLtHaiXLxhsS82xg9vScs4IfWNrnIS8O+x+K+hawrIhx+JcAs9
czcdjhWRnnEfvr8zmGwP+aOXDBddBKP1vHtVQQmB2QheMY621de/8EgO8nrHzx1q99quN6XjPjEZ
lguj5sbna3m971iaQa2f2w1jX91Ynmrj0KMtNFZfaKYm8fjgSEkZvmgktGiUCQKQ+xwNznt4wSam
PnEv9TS8icrx2IbPT4+Rekltulz+VHX1Bttzc1YpiMJjGibsPCFLTiHT8yiqE7Q9VZDZDz5w+ItL
4n3iwwHtD5iHeAb+M2a2F3IInE3JmrNTbT3GD+yRwXb1+uh1jDmEhsPGnPhwEBs8Dk7m9UC1roXy
hh4/rfflby3VrSXSXNbCrJ5FCOI4Wv/j2FwBTskbVZoKnCsZC5zewoH4V5YARHohSKOxfiV4DQ5x
RPErZ3HEFNFDd5NWmApVUvW25E1kfQ7aZTfDCJ6LUen9vrHxSDGMkNBDSf8lKnUJHKIwQxUEU19v
PCNsORCKXjhsi0OGYA60bo/E90qYF4Z/yHXzFKefmYrqMcnTGU7Lo/4aNMNY+CI5nOvkdD47M5pf
iE0sLnZxR6T5s+1BXYunCEG7m/vqlZCjf92aLtkAooyhWOIfTAm0zYRGurEx9CokUDDMqwBRhqo2
6pBJM596Ojz7tmeLpvhU/17mAJZOssUN+4C7YxCl3QmvSCvfFBoSJga8jJBESxn3e1j8CtOPYHRX
AtT6BTqIwVC9P4lpwFNB/ycMieBl5FhFPKxDb36Vn3S0mPejvd+erW6qZ9sA2Ob4B1IRn7cYSaB/
l68A7fPBZNlp7ReYcN/qVC2H6VCR1SgNM8IYvU85ssaD6DuydS9rskUW7hrDM/yR+yokidMDPRzX
rzJs+1YbG+n0eXgaMwEka18BwntjNqjblF7rAa7fu1RqcTkvxZeFC7s9RiWmFhwzdKeRHJHHxVT4
GIrB2Sc4O3RG22ImNjA2aHxbjTqEiS77OoJUrP9BC8fTsGRirhDV4JNixiIYc2P/6pPNLH7a7u+L
ef6+WY1u4P3bRaXlkxqeokAgXS7rNOIvMQa54E5PuhKOsWfIyMNnVGlyzzhvhtQdSyw9UjwIJQWU
U3r9WUDwwuFiyywp207Bt+MbmgM0E6gw6ZEecL/Xy2TQi8ow3BZwslPiNpFkhouSpAdWX4lgy8r8
rQHySo3L7HqF9XfctYO403o0UCyGcrr5TWt7Y5Vn5aikaZVop+WroOe7QbVVsUPakyK0J0fR2TOz
LNzZ4+UeTE2cQw11n5j2EapyjMYBvpctY8jhGO5bA9E6kedkMtIFUTDffbIGnbLrtj3zr0nRVla5
VH8sAwZ0rZCPtt6Y6QfcdQ4Xthu2YqQYrtTw/WtuTgc6qM4MPC7kZfvOicrwWCQZqkNy8BGFUhar
nWzFZQA6wQ6ssV9LPsdmB212M7/u0ezrr/9y3Lh2AWhdfi7h6ReKg0CwWiCzwvbbbFCHXZ8oK2G6
wYfA9VhPp5SrQLVPkBTxEjiCQahPL2Z2e6CeRalzyXsGDU/Ox+3yYMzhUOHfBw+mY/QjZ30Y1k/9
g1NSrIRgP6Qol7dUGUTGUlfIrbFhntF0zMKurx+0ROmfv+09Jl7OlGitR04WUPpmdl5zIdc04Xe3
E1HznTGmzUi3HCVWIs48mHKLzziNKMzsjbb2QhgLObawbhkO4UcXDV9jsDIUofrr639GX27NGn2q
f5322H0aXyJmVAfpYGbShGdVJ2kmz9qv64dFXnKw6UNIQNPhj/Ll0KmUFmJ+VKD3o3vEbiVWql8S
0yPD1gV6IWD0MHf9531y+Wlb+5GXVi/qAxmuFn3ojBExd9xVxeWEkyAOUjwlxHB7Bel9nofW1NEH
wL+kQtyDCDdC9avIzWFXxUBZD/AYos6ChX0Djo9+DhCRTRNn8wXR5fAmBRbXX9s5ywIqi8IihF9b
9EZG8ccylyLuXW9tUOFRVS3IbVhiXw4+zpsqXdS6qKnSiwYb4IMQH476JUUQN96hnPkslcM+uUX1
1Z0woRCXXWehOuFPkioRkAzHYweNTpXjoUAKp3IvDqnq/tyTYROyzSLOg0pQsEn04u3n4b4k9cac
lYjN4svHaoS5oMbvpirzi4aPoU8htLLd1BchrXuRcubZXVRW8Bv8AkQXh/uWqtziacz0F9d2rOW0
Dm6PgpzmDFbzQ1B0m+hCH0btsngXCzXza7YlVSJZ5/oIpGUEDCYNWc4czElkxXCKybKLLgpJY/Yy
UUYROnG0Y8rwX9nWRyE21Gximfsb3k21bMde0vYy9Gswdwde/So6dEgQgn/Z5H7yXgD3f2c9R4pN
barXsRP4NhHe1COSGXmYAQxhoD+zEulA2pdm8u7SGuJXQnklcFWwGZ+pr6+EZ7c1s75rPyteB+0D
bQdVH6affxdF/VpiV/Ha+bnwVzYzc7KB22Gs8jCoEwQskvHtCksVGRVqmnz8tEJWi3/hbut1+4re
Nrpg8GF/U/DrgZCoOtajnGzlEOcSJiXPaL34Dri68tYvw7qU4LrxFjjcxGUR8suB6UfxAALEw97b
ujQT1171O8tuwN+mnCcLlpd1cK9tnOlSbJ4Dfytx1OQETaISB32kD+oPgwo8IhuBMV+p+FxLvJbq
6Tr9UF0n40DE3pn8FNHb/domGZWGxaGzAJKQjfGRsz43HF50iCLS1Nd5sQkxp3uAaeJfKRLMp3/a
aw/YE+13FR8q/1TxaNxsd3zom3EtN5OiFRliSOJSMWJqsNh+ISuntxGetYm5jSrlC4al+YP9wTMc
+sfTgv7r6sfnvvDeGgPNQR5sb5hv0u/YJfjXI4LGHHs4BxLj7FmvzUT/S+gC/Vx/L5TXJDif3ewU
1i/Pga41dLaLKU4mnhHYtx/4/e2DzuA+aEcMZANxtqO5SvvItQMZWUxE+5bqRE5SBlhJFtDBiP8s
F48h3E+Or2+tnc1wtQaXU+8L1DnIpPRjxv//vLHpu/qiuY9lPVb/q8sB5TqxraBu88Elc2TE3NXq
AWRhlF3ZRO6V9P1LK42JRLP3m0jzHETqaFk0zzOgfDQ4we1K4WzuQR2dV/msK9NpScMAMPQoE9jw
yV1gV26wHIN/z0OuI8N56RQvNOuVw51aDz2F6qh2R0oCiTtJYPz6RsSNNYYGUbGIhibFLmr6T277
P2ERFSJ7/XUP4BWy27K51s+pdsVZoqIjk8UEy0yTul3Q/krj1KBWTSpXr+2qxj19oWDZ19IEa+I5
OannHSyDP5dKJbP9kIGWOS96NzxbpsCqZf2FOza0SIvMHkmLDvsDberZADLeD7TrdiZ3qvYXbphI
OY79ctJqXo2hR7ymD97JUt1ciNeI+B6emmJTL+RVciLgWU1BgjTxRDiyPoSu1wu1Cy+iIIsAt0vo
A/YZsSITvhD3W/zdnk8336N8eB0CYRIpkDgxgPjvin3dX+IUlGETQF+mGeKVGh5XP3HAYuVXzmsX
kv4WUPTmT3vUfUpyU6Pq939isO1rFA6akF2P0+rN2kzpq18g5bh8bD9UM5wLmlIlK+VEq51OdxFn
nnN/ptmSc5fFfxYYzI8wcwKB6O/DTVAGn70sYW5iyZ/TpYXUJf4HaFHXzDHyICnb0uNvgaCD+PKn
1I6FAkStRpi5a/V1+HiKQsleP5BF+9+UL569e8UqKvjEUKRs+yZl/iAZ5n6CtTsY06qt3vnbpdmq
p+MSF32TATrnUpO1ZBAhYB2SmL8O1KquCLa/DYxrg/mEAKlO4BoMpdgCtKpWqMQwSp0vsUlMza0s
7sEnAWqxhtJGa6czYlSf9CNAkFbhHvllKP865303jxYy7SW16bExrZWsCkte/oPgopU5BmE8qjSq
YZClw/jvBeThqeIrkJIuCae9lqEf0A849VjinxaGFjBc+ALYmnbAOLrS8l633nzM5+9rPb39elbm
cXcfaAGg7IGPhVUstWo/vgRObMFZfLoScub3s6uLB0H6ZioVa3MMi7b/RjYpgwBMGTNt2aK1BrGp
qVZ/1CYTacFiD0ME5bkMbOv3K1kQBzPSUrSDT1C7p/3mOz06vOsyTUJK+7ykOfoqYA8yw+Nn+0jR
QLqbsngARAbDbSQ+wX6aSX1gkCOa/3+p+2mQxa9V6LU+8fGn8l1pNzAwiqAiFygKsqvBj9YniOcI
VwKqwpLvHiUHUKSJFbOQOYaepANMJNiscXsjO5NF7frMv1axNSW+xHUsfiTF7mYI0xIA16o3mpEk
uMGCYrUaHgH9aBg+lm90y5XaUUXjFBynhzSo+QWln75OzTvXAoC2dyfdvVIv+P7hikItHbR+g6UD
7HgLULsQg01Yg6ihpT4STxnh66XFfF1YSskGzmBXw3/Z/7VEPzSLblibqY8337qAACHQhpykxP4M
4QSpTzZE+0liJTXGyNb3idKdl6QMh4b1+1YYFUIwJQR6AMTD4KmvtZIanqbKISb5ABjGC6H/IMKK
FjgdRPOviV6EXxrM6t+wTiG42cu7bbZe3U11HCP6tk8OMV2svDsKLkrYY5hveziSac3c0+8MkBIG
Vy1WBLHZD0n3U0DrAqmP0BMUvZIt1wFEmcNmlFfsscuV8AnKogcMHgM1NcirDcXJTFVlWCABpFSm
VLhIH6IW6QCf/r6WSh4KH+mgDsg4GZDZ35Azl/NRbm3Y/4ZynEI5+y6rw20lW7D8jP9hOI7cScdj
CCo4ScjKsBdAV5gvMt5qhEwW2Sj0KDgTSOGmteYbiJJX8/Oh6G97LZpSdehoq9AZuIWCNVcdTd7P
tXVSXG7wI02hsauS6lkrA3vqUqA/5cYiias0qnhX9+Sg3R6IBNuHXDqGMS4oWVLVPDWaupBPtmFu
noy3brdmSUreKWOIcz+rFHTKhDS9EwDxrUQC9hXLO0LipYOZz7Uxmm3gn4gIGgAqeiI/qSTY/0JL
fESfpPwUY5aC9Ja1QlCguaaCdf4/i7ltwvqvDbHySwzzXCGyKTxQNcoDKwgkPyOVIgPfHZ7bTybX
FKvM2cZ76hUxZt9vGkHB/kibbRGaMNPph5D70R0hjVKBoywwv4s+/l6iBRkDnW9vojZxo4nayQ93
8hvndhvtb/7TDLtHcr1SM5eZ0HZvXiaAQiGLb+QQcp72A/YYZtGdrWn4CXD7hlLTKaAB6qWaSML4
vtoFq3pnondaGpxoFhAc12ogr5uqvR0SoTUefWYh92U78KPLIrA+jtV0pIYg4I0fb9fGu/G+GZX3
hEWqRocD4hsGZiVPw2f9TTK/Mqu+HrKkc15Ob8HjikdJynE4cQxO4rbitVwVOj/HaIDd4KZyefoj
xnBxVJb/kF/yU9DNXRoJPheHnRhD76izGd+zObY+0w9QmPSJSrUElKAkj7apFg+OMS7i/BWHjcsX
1hDIVHjjRX3WBb9aJgIi+hvNLHdC+SIv0+dihj5ZqrByHcVP6DdFpEOJclNNqByYou/ePd7b8c7q
UyHdJd6+YJsI37uoE3cQ4n94X58SY2M3RYDzwDk8DnYwkGZETp60gBz5B1N/5/f/yNDAiihs7rz7
ReblfoLBY15FVOX6lcRuD11snFu7ZDB47aHztexA10uwerPydGbQBjLZsOgakjA9Rlon5NI2rToL
kDO7XRr0zk+ejypZ/Dnoc5cWiJBnYJ0I7vqvcO4Oq4KjTxKL2PgLz6kpzX4c85cpZi80do9L69Xt
Q3OX37Flj4kEZ3K0XMfncNrOW9g1sqloUCZww2niIaGCZWXEnY6u8+ms0EFaZaHYQcEWGNeyM1wf
XbSXRnyJRApjaX3p6gZauIz/M694U+rBS3LrtmWNSsWklkpblF5sd6c+LD5//4skagTsSMpn8Ndv
0Wxq3pqXx6akndH6dc3IAGaGJeGwzaY3VCIYS9GMUBGKv0mJzpdOy5Kz/8+TD/3H0TAvwdRyvg/5
BX2f3+mrSmIrmend8MxMIzIFFeE9s2wtoACDF32OGmwOXLzDIoxcx14BSVmGl86YhZxf7k/EZl5t
WN3g/SL9j0ct+7mv0yd+WzwggBX55lg1OJAiRb/FACSj00GLw9js748wwjuH68Oznt7TfnaB253O
ziIOem2tQTO+3v1TkZbBSbfuSc0mWlonS0t+sVe+RmqKdFBdmsdWZzER+ryjqnfQPJh57DgHgZFn
hw+xMdWWGC3NLI+LxkKNjJHwJyN93z1mRBmaSE7UcRt7LUlUuOUsSEgYvDSjS/okBhccGfaO5dsJ
i3NhX51iund0YsfUQFLYM6HZwX9gf1OR+bxYljNhs3jd726WZBvo4OJiIGyh2+P900X0nvc+/HAE
MJ/YjtUtnZSg8k12weQ0E/j7LS8kAAxJRUXblSgluPkQpxhhr+bQeBS1RYOUAjornMgSkGBDrLJg
puZQD5NOPnQpiehedCVDRxH6Qzgk5/lvnnGxq7oEY4Mgq29OkHmLFIFRBaQD9k6mP6DIEoZhE3RQ
YqIDKtHTMa4kutRnDtEjAdWccqGQvYgbY/sXGAw+d8hMvWi9wr2RqVJvr7dRxqtSUceLGyFKMN+i
48mNz3uGbi2PkwmwrwIiph9E1mrDzhUwD1q5zuo4j0vAbHdkvK5iBEut72ZlV4/7gUkku5mTNu1I
qMnwEdgZxCCPs3PiCHLZwjvTDdCfy8NIG7YaI/e13HgzNCQMYa9vnnuiwK+5hLZK1nyVFSQ6Uwfh
K2Qo8s/adSqaFyylhiAgblru3e8ypQuzhbfZX9pGydwDYgoYyg9nc5n9Yv+g7qctvPlzgEczP5h4
pfI9NlW7loTwyk+oP7cRAaH+G7oklf0NBeCvYUrvmGAG6NyifDsWpEtDSGmiM+zUSlakuZfTjL4e
ICRC15gQdQtQ+w+SnE8q/uJPM85749qioSQIIBD2gFHq5McMpbRuKD2I6PhiHxBG2VMhtqfsVoqQ
6Vh3FLLnzEMWdMnnltax4+toYAhkVJhy80JxK7BjjALFlq4pQhSix6q8yn6ed0cUvwAmiFU96ZfH
4PHgREz3vdsKt/d1nmCTaRqqLnDmU5PG1tt7kIRCnd1PyNAY9QcGxT74IzZurqomCTeQmKwyZPaw
B0JAFM3Aj7fryfQe2WxZ7XqiBa0eOpet1B2dj5hkNj0nwF+ckMAxVdzXCSqtzXhTV8wdfK0BX0aG
RrqYWscDc0RYXkQrbnkNiRkFi/DG6N9sHn4qp81gcKSpjmKYR9/FHHr4AJdP0O5yv7qYFEYnjSDR
8ycH0BOLEOz30snFb+JIaDgpVYSSBjSozbMmAsnNw7vuUC8176yaqeAndd6nxyR38RuJRiJCKpsD
uIPiTgaEpAT5uEEncaxPw55Pxe+WSDdWG6EfatKdSxlvXy4VagRdRghovNzIk21Co7IAUxzeLrFE
hRV94PEklKVM9yA4MutlhhyScduYGJ0myIB5TVilsuudaYDxvGniRITKexjSELFqtwJTL+ok17EK
PiGDmkL0IFPI9gEUX4wQvgl7MIvwZhr6Bq/1QzjxY0r0+3YICLctwiJT55iDnIEq7Vxo1Ue16B/K
OHOze6aEPs3ki0EfPxJADQFeu4oSuAMWyRVzcHVbYT9vl05A13XZxYPlTTyKZ3ZfhE4mw2VT+XHH
idnapaowPoCwp+MSbRU+ZP0wY5zzoxvOSF1LJRLHhE7LgCOXHCgH3+rptuAByBQ7/JZG42WIqzvh
VVpEXLLUanoIMShlmiZss8rfTuYNtXQ86tUoWpHRcbJMlxc5iCRfEyGSfm1cLrVxZictqw4gfmus
7SamuyGzVRCj1eZUScP4Izr9/7Lvk6zXSlZ7MLM7YaeJ+y5EHczL1L9o7SAfS1bSiufywVqoruye
DfiHyS6Fx29IwOioKoUEnrL/Wy7nGYhiAdcYzMLEbERMdua9uctCQccWYXoxID4QD8LX9RoYdQjT
Vcmk6OqCEUJv/RqcwUeAXn9iPZXV5oPSms71nlLk6dBCcVSP2iQOwh8WULnd58y9X9Ay/zHRXESE
h3Uh/gEO8gyReOEfHk9IKH2U64UF+lrVrVGND+rzdO2kPpF7s2cvzfe5k/buwn03xRZA6TknIm8m
+5VNmh0SkQxngQ0NymEKeB5WHEdmFuqu7TZZRtBqniepm5MxJNpnI9rfK3BwhEojXcA+d3s4LBbO
7TOIctvH8v15egjZmRoub3wViNyZYG8xqmWCVG71swh0cCWfCEyOG0MPZCw66RGCrs02kH9+MRgG
EJFF0i7bF0SRQj3CBi4aQ+o/6FycvZFKk1KNeiZTTPOIGsV1Py3DUkl7p8psTA4ASSO9+Pc8rxv4
NbfeKfgSS/h9BH9M+eOO7mAgOtppgIQt58kC/Wrbzl0SMqiUdN5OJTYQLzz5Cq1Ni7TeNUI+vzJl
r2d/8AHVZZyLrky8otdZX2gTYxp0zn17NYE8Hf6ISCQXH1sURhSwWCB+UB82L4GVeMyIOCUif1Xh
0rizvKLppEsZ32LevaIB9uWwNlKY+C2ZDTHkO5Uokewqe6F9IZ/7w/nJaZUz3l6NLrI8WcaSkebN
ekN6MnEi2+sy4HTDKyKMJx12TWiFiRrATZGiE22vu13vt7eBzW9rXxGnyAtfNNhQgwYqBAJdUbmS
I0xQenMYrtPsnXkDTTPAIwXo2qepyGoQ858NfGEGJ2vIT+bR+0H8TV4T3uSAR6mconGNCnJr5pJV
WIYUWw/IaJFsEAn6hdRyYmGfAQzDZfAx0BS9MXeg97n5OLwCLoKUN7XeptM8oOa0nUQXnyDPIakR
TKEXG81aSvsEgTQQ/+BQVe/Vt3XsY/5e50rUEmLspcDa5uSSZjK2fizkx70Do9qHZoWHJtRlX+/O
+FKKKKlI9FLLg/EL2i2hRWDpwb0dR73oaJeODEY3au2rye74BP1EP4+82b5FYUxRsi4Z2HVGLTrK
jlDCyKZWGl/bse3Y9CxATUPzsR6j9DYZS+YdgvRt7jg0bJGwJpaRSvQ4K/fdQHfz1mgEz1vNwSNI
8o24ud+q+rZJE7bOYluQZC+fuPaaHXjJ0YfAW6S1ojcoG2KnJFCrV7UAj7EY7h7Xg7FBHCFKIh4e
TIF3gqjfF31Q3dcajEC/gM1xsXQfb/bzlM3h0uMgPq3ZmtaWtn76dmGf/JM2o+DthE0kszqUaT7H
Tz2FDSSBW4AaqdS/1ADcAQACTTb3fRjc70MriPP+XsSlh6iTLMsn+Z0v/jUitLD3Q7P6csZBF4bn
ZCC30EtWO0aZWT0J+WAYfNmdOCiBtUkobyndPIMisLkXWr2P+7SHbBz2R0/Xr8vNSNvY16ejqwoN
3TVOuXlJtPeNWU+IJdHRAICGFbeTY8+e3AOJncfO+u+o4HAVhvTtUGGnUor3aKPG/QpGCOVTgVhB
t7mUdvhYh0j3pfJgGnqCF+d7RC/CHYj/YFdvxADOPnDMDpp8UToIQjB2Oh9+c95qTzQhCpw+Fg5D
E7sMXET2p2020V4FA25u+tJBhWqe5+avbcw0mTcX+ZpRDxJLIaVFFUBgrRfXVo/bkUC/XHCwZJab
JcvNEGJ7wQCw925+owZMgBWI/LJ+FUVOGmL58yUvA2EN9mugY6Zd4Om3+C+Tj9K7Vemy6dJKRV6E
OZs6JqqbPgn8H4qaJrmwT2mMauYtXON0CErrZM+HiAO3SE+kqOvtIad74b1ntEruf0n8oPpjesUt
NdFgD9gTxd133e57cI7CI22cdbaVAzVBG9EgydwcrU9gRBkTEbECTRDdZyRHU9FX36XL0Eh0Ww8Y
ERlxWr7HMHt3ZrxZgkdhLt1C1GHWI7YZI8eydgUFvipzIUNPwTM1xTgjNvLuXDfUXIn0NJGWi/MI
PZVFwLTsPMBUF4mtPas2OHyr0xsGuiftKgj6WHz6ECXec0JNp9+vAectow7vuqfbSsfKCnXGv6Q8
UeV2Jrniq4zK7KlhM7IyW8LJR4tQD31XUVh3qUv0+nRb5pj428Df8rkFzEhKASMO/aqaPxurnTle
UoviW6cSuHsnQLoRdxIs/BlR0S0li3UaCszS+2+JpJF8c9TKyW3FxuL0nD5198taoFOgIU20qgQ3
3DkW8d1AB9EDS2nNxoycmRdF4nW04eWjFLU9w6dPae1OuGTjDpwd7XlbZ1zU2n6xBetGOOgkanxs
spGSRLHLDenJgVc6oUlqV9ipYCtfUPZq8LMUzuy9EDQiyOaQ4SethF3Pq3h0saRLluy1Qnx6FwMx
HE3yU9/8ER8LUe5DWtg4NbMIKL9inahhEDhqHbkENSkWczDZ9Ef/BfhFf43D/2aguhGpZTuSc0lp
ZPLrco3NstxlUPPYF7xZhm9GzbQ8wYeV1yVjSYyUUaNJi+SWcnK57vbJStuFNytcDatAFLrb74bS
PVCw/vjU7hdDq1Gs9AZCvI5LO9DBJebVsvLNqSbyo3A9xvVfVHZ6PUwERUXW3tJIfv11optcBuhT
KhynqjNw4Eu7H06Mf/1TJ3lEibXBiSNV01MgRDffoL2PGZJS9cABtbK0jdCdFb5jv+TjnWTv2mhN
9HaTf/U+3FiNy4NMzI1tcVTeOeSOA4Dr0VWc9XFqnUJjkugOOqr2c+LiljZiguIlu6krrBH/DEUk
KSm5u2QHbrPAO6X/SvlOxpicLfqzbyXVKpPsRUlOxSLqYQhYbwOfhbVn8f3/EzlHG9ahSzaoDSG9
lMx3ISFMho5D4Hs8FWZdw641LWD4MI2/bRDObd1hYcJ2L4Zj+zXu1PtXkhgjOO2CRkmTpKkFR2Pi
kqw9Bd35nMc84C17vkCcGtKMWrDmb/TPw5/nmP+EJ+S0Y2VYOgcHhJDp2epitvTsijTB227ZHcLw
oLw7UedahRviMVmQeuIzM6vrt1wlSxsblJN7fpOXmSTSWPGPEILTGKi3fpYM/w0umihL9PSVJqks
O3afEVV/5Af+B7sx6c02KHXJww0cIHyTV5vaa+HsWx2ZzzTfUmpdQtl0gZqLWmtERiyKv6z4k6hG
28qPgqIlyeMn5vrI0XpVNuZq5rvlFkJgr5Y/Og0+TZ6qBMgQ6zSwPLZ8xEvN6SWUKB0zFS8Q11JJ
SqluxlsthlOou+ApbIP1wxzeeS6szJw17iqAwptgtinCweiN+PkFUW5P0g5Lbs3VKFxZ0NufIajy
5WuNmDFDl7o5grmYq57JakQT1XuN4a1h/7Dv5vRJpFZ5RwYTZVMF90BEBcMvz+F7E5PljLZPR3Sm
7mHBQwcruvp5eZhNVTlxELA3UhT8hXGu3a/Cd0hlS2xQd2ursJPkryNjlbGrxDQd4REIttsl/u/H
891qcO8O4LQ4hwnUITEvgloGZAdyQqf+q4kVsgYv4/r/bnOtwwnALiXwJnBQakTsGraIt+9NyUu+
T1mYXmUDm/AupXCKMSWy8brpZ0agdxqm9+3IQm8OV8kssZhAOOIzBorH1fNpXlPB1BhFN6yx7Pfb
LJ/1ZfDPeO5p3MkB0fcLCegqwDST7sIGVrSKHhQ15MMqKt6+ehurBz28whOqauDwTwhyhUeRrYui
DPacRn8oo3mdQSHdO8wJ9pfQ/SXOcGXN4Z1W6cd3GNRf3nL4spQ7Jmb1cuXPVOJE3I6mElRjidDB
1NY/FPB/WlQO4+Fwy1fBTJnQMwuttJbWd6mmLnUuGxoDtJxVqgUaLqJHSHV0aNIEQoZjLkbCKafw
cF7uE2o2bw63l3E5RkAjniB2DR7qdvJtG4J7MWkDnOHvLjpHAR8TCnvCtd0W22gWTSDdOdJq5m4t
BCC0wou6qhNVrWqvOwse8gppwR9TjALbMj9RUa8eUqN4wHeSaomI1DTZMdtEI9FYK2zUFw/iQMfN
pG3WhC32xl2Oq3IsrYSe+F9tzde6zrj6Fpz9qoTspEBRBIEDtDHeq+mBFx+QivtCA3hJ6cdgbDEe
Vv2FqA0EK/lgAsuf3930YaBnHpBp2mKMUMq2fh782n11HYF3Lrg+Xid82aOnAWILhfx3iNaXP4sf
h2cY1QzKhqZvu7jqHJcm3T+4+Dzb3YybPhL6dqAUsKUmKPCTcsBifnuF6N3Q57kUuL5+T/IaMSq+
yiR8O4O9RYtvllPV2VfLUZjJomSQ/osAmonrElXAOLRQtP1etOClE8+9hTVLJYlfRTSA2KiwvRLA
92uKTnbLECQYfkrYvWFJ/AjYJnVjrX4iWu6CsZVMr1Hu6D3Fn023Yw4ACZvFhHlV7G9E5WD/p8F1
0bsf8sMVfDRZHleM9zkTgIhSqsbXQkUpFdtCdLYrardUf+dLg+P6I2NYR3qdyxnQm34GAna9kkjb
+1Dga2BE9pgjar1NYenZdGazV8bI0E0mu7YPR0to71S4OsC8bsUu1QyfiN4mV699kgrktGEqkLIy
TI4mFCzUfnX3rW8hB9gzufdE1Trcv1Dcxhs8xT6MNfRRct71UzVXxJCTEtl7sDaHQ+2lGdMeHWnY
y/VfynTdZlEaWS/tda4Hz9EuSlWrUFQljy1LsrGGNSTa04eFFV9db7V+LE/IabvGXhz0Ap4gSlOY
usSznAVSCuUQpJCPKkScwBiCw7ddvi0Bg2PdcLVhPYkL9UVYvNCL8025K9VwTksq9ED/yMlVWZ4G
+OyyliYb82Ig2qYLMztn35NVysCN9/Zjgl76bjENVZMSRrhkSUyU14wyEiid6IrEdRAjLZYvwKrp
qayP2A2d/mzzFKtzn/1+0CS608i4JoCCsaGpDhzMrviykXLeEFva+2v4yilTD3YVlJjEjyreYOX9
eVXvlCyC7LMwlK3Aa5YJfFYYwFxgz+0WZDPqKVDXfKEZaES71K/iaLusSaAgeeiQLA6uVq7j5u3H
3uzxt9cg5BW6BoAY0nbqOPC0sYojeC8859KtCE5Pty4MPZ9dlcwPoOydvULljUbcPfSMS4LLV19S
LuXNuF45DWymWfY2ZhY+LAwqSDDy4EIQcdWaAL2JKIfwIxLKuCssJdqPadNSSFult6vZEK5uyhdV
omP+zu9l76ymSoZYjuw0SkBBDlmVNvGp+SjdU3w/NtQVRP21svdmCyKt7Y0DfJW3ebIoI1eUPiFO
RlRruw+LHj0tvuZC0vL+Rvpsuc3I+Lp7CDg+3+3PtfmCrUX3KCoBCzIPRIs4dRJOv3mkuNThhVbT
G3cXHe1JPDaDkqPnv5KUa6F6ZkqMkkzHvEyB6At+RyPwImGWBQNX5Srr2AwCP3bY/YLq50fKSCan
KuCfOR2v98Hl+D9R2h6YRJcDQOuWUI/o3/b8f+ZeL6LzSIQw8BxVOZPQWyV0dbp2QU2RJ97zfzAh
fMmiw29lJhifV/u2i0/gYuyENn7vKLIi/1PukerHYmW6MTkZG/54EiGaE1wfiRiyung8udY4C20U
Wu8D1+kt2sBbLsj3n5qCcJ8NAFJou5u2gn7zNmcFF18M2gBbG+MN2Q+jOZqGKJNamH9ixLNkNvHw
tf9q2J6OwoYckBh02eunpch68PSZy9KnhfUOKHVyZX8ijZ7oYYJsBwtM3dHnwKS2TpsQ3YQyUoiu
/Es4kKPl73duyZfkR9J8AshiOR8wToykxTyYAHpQtgdZo0ppllHvO9U4z0vDbqg3rIzqmaugcFML
Z0fTV/As2EXvYNTw24Hy8HVOXxkqnz0MZZQugwNGlDE7IuwP4B3HPvFTDViOxJZ/axLcyHWEkA8L
nyT/Xx6CDrGezvq47JFVX5iCWnkaQNmceqAKVwMVHR8e163/dDiboh1QMyfTghCVwT1yvfowmNrm
BcccMyhwIvntsND8OBTCtIXW3THotwufiyrouX/Uv/52w29Ss3m/FZ+SYtC1AYP9d7CrUkJ+z6SQ
ivqnyk+0kfEcQc2iSqvT3rS4w/eQla57aijl7cYh6zPy5pkneqm0g/vY6OF9s68t7DwoWzz3Ery0
t8EUyHpWgID45uDBduqnTQ6dwfET52FdwIPsWfYxQfojJlb/lr1mU/CLf4Bo0mcqxuiakCnvK4f0
/16uxSwVtV15eljDS6AjjtgvTC/rHK/gIukN84y6NSGbatEWSCLulqWyxOaRc5mfcFNUxFin9kdl
+km8s8ukRglYQwuYl7RbhSq9TH4eXk9RXuriWGq0IsbFbZl3K5tk3MuMwS/w8bSyW+nb47UvNivj
fmegYN5rvIWrT38FalG051R2/LkAqvzmKl11x+2+kQnOV8L+4iJ8/uNZe4GLjunWEeJgZeIIZDjd
L6YgqXOT0mayZEKWrgAIMRF0SlzYrwo2rARNNFSHFsXPXrKnml/1R1AI06ZKHc8aM7frk34r/kTd
tnFCgM0/0/HVS8n5SFMNj70VkiaOU/hM9F2eWlPTUs1ehD2G3T3lCaTPF8ovimSQbMLFmgPF53zH
ZmHr6yHYo4tiKwprfqclif0P8SJn0JQz+7j13JP4N9+nNej1aPPzm4I/gk3s27VPNK6StAcTxRwm
ESWEnMtDwU7CtRrTiVflm0SYVtASXGO9rcYI+PSOePDOXUjQGNpSxu9rH4hB8ZJjKON2Nxv+rX84
m1W6e2EDyo0ihOSygwACCOpHlwUzuH3XiyIspJP/p8GJOifhdYhM1flCCAQVfa6v3nRBtExqQxXH
S1Km0r9+bhssCCQImuECKDWB2NVQdi0TM7UXQiVTR9mcDhdZxuDEBWxzPTYz9Gwb37+OeV0l8Qgf
LYvq0QzBVzSxhdjfHPtjnKMmbkuh81Vv+TNAh6M51YVh0kfdvBApBT3Rq4Tkmb34MQbUUiy0VUsN
U0kT7cvHsMNHWVTT8FVkSuo4VmBmuxOArN+pM63LAcYJvlFqsmCLTvpmUd05k/QksLsa879pBKdg
78YU0PMuYJg6f82F9pIw7wy+g7iBCrLgY+y6C8NaxYT1gdOZqCEWgXgd7iTb2vTCRYNLN9LiStmE
nm4jxt7jBfAuE2auyXG3K9c01F/Wr5Yy/7h0IbbieqgUd0njUDL0k/lCcGe8PSNDMk+qsktrhWO/
JWmo33CELGQKDolEdy0xNu+W8sAxVrfwCbkWDSQpSCQNb2BfxSMYvDRA5RUaSAeKrl7kHeTvGbd7
cPSW28E3p4WEXIGVu6fNhVjvs5D5ROIuxQnqY/pFjNdWW1/514DnYv0kpCWI52fCxg3XqbjpQFuQ
0ZjawsEPFHNe5T8N5tn3XSlvRI48CnIg1CbDHPISLm66Z32bnplFD73Rf1Ck/d3XN4Iv4Qjjzk/e
UHMPrVFSGuMnH6bPj54SIWnzPz9A6SQQ3xAuA5e3VUbKskQqdv5Uh6VvtjPCh++zPamssVqWptRP
OcrCa3y0Ny/MuqfS/MTBXd7YISQZpzbJLn6Y9YZCEK9qhbsBRC41iTJj6WX9fUmEzzMeQaWoEE9b
hYvaDsr2YpOwyxxkPCx5CuuDENlWrTIlBcUzTPvW0eKdon0crVNpt/dcROIHQD0963w0CztJL6WC
2GCf4h0FS/onOk8rj+Jq45rkNpUCVI4A0Yg3hZq+LEhgHPqVxcCqnh2dMySe0HDxJfif2SqrS4J5
i+XJ0T6vdXt6fQJBIn6UxJvN9caxzyHeUXR+MKSSTwVLt8X8H8YRhMx52uNMXERz0vLeX/RagoRR
IWTNMP9+RzEzIk0C1tUHABZIfwGC36JPTVf7RtClTr47T+NRwTROMJ2cQ1h8XKfQSmxgQmPqhyrQ
0Qo3dErXmY07DRyjGOLeoNTUYQDHZ+fDhzMEkhGdUvp6QdWJhwnE58s3M/YaLdZbT6lvytWXLFmC
RktBEFBbYZg4N0JJbN0EPeR8x5AYpWPEy7ax1oCYtYAmmlUKsPsClkkVVvpPhm/HDK4IsE80X41U
9tf+tMK98XXwpxKgEiawwA3Iu/dhTaQIPBfOiGWNzDxevukrXP9Sw7aqij6s5LzM2zhnAofialAp
O4XuQutkSiGJZQW76qCI7ZydIpS66rwburkbG16vUR41at4ws/FxUYu3nhoCBIqmOD9+zP67ZDjq
Sf2i5xtyWRHfHwvoS/U23fs2SfdYoN3+WaFvQBJtR27CyejrrxDSuV1wzH3XjhcKLvD5Majb5Hjn
rklp5UmQ1KBhlBOBgkTCAipKA8vIfM9DwxtYKHhjeNrXGJklbD04UO8OrMSLxEM/N7V7f7CeBiUI
7jCnyKOSa2xtE/OvgyV/JP/TyopWAE65/qSgUFoTPfeuqwNdbt3pZm8fnAEU/1w2Wr3eC7d0bRRC
ixSwAY2kJlFu6b3s/ZOcutYM7bgqC1l2zj10j1+ez8hLv7UYsnBjgWzzjeYmdSfWd2puCav2pJJo
97EJv+zY+otUM8ClInxmRGQhMMaDA7GES8L/qSWF74AnfPWNn1+n2nD+6Y2zwtBMKHIX006bPUr9
JW4DXtxdU4P3/QOWiVkB1zJF8/6Mz/WSLd+G6uLIZrzPWjfHQiN5cbgKwehwHJv5gpVpjiffGSoK
PDaIvQkFHH3SDoyIhAb/9L+VrZk9RmiuYZaW88/vyoPHEMs6Q9hzF3iZslgc2Zkd//fGb3fFZ9Na
O/onceTjuoQpzcWnamj9uJdees0jzplq5/i2G063tP/wgea+H/FTeTezzB67XgSmCROyzVrzDs0L
ayhKkSgAYCKmnkGERId+SGEIpu1Gyb+5uYS4XNj/sYtxapCP6OpeeHuyh+GYWqOOXyXnCzVcMMEy
CYcwLzwePw6d4ZW6/2ZfD/1uXTc8pXecN8Xw6BGqKTBOMRUnxtAcz0YZcsrEtdUhWQkfvHgK38cj
+wUhq60jGQugB+Z1mgEJoqkPbRjc0/uBIO0kPsiRNhEhg47326neizVO9ElhnlytW4qMHv9e6r5g
p9nYPquChHOVUui3O5KLyrSHC4RNgXWzG2mKI9ArhoTgWtoKhvob59ebV73jV0Lhn2hl0yoriULs
LMOm9cuDTyzcNr17l618heBJTldT02Y+lIemcZtR56NIFU0Jh6XbZsBE8xAzCYj/JWm0VovaLniv
sQ5ljhWOZqGXRO0e2naML4E2J976in2Y0EjNJENE2c0CUS5DjAlJQUV8QxsGl2iBb8owYamFycDr
0AxKUvH0BP9k93tGP/7eCjw2Cykjl85EAOzwraKtT5nl0lKn9082xD5jfuLB8z7deuWKZrR47Doz
v7PyobusGuVyv+NXK1y24wjp+4Hjfzzr4qHJDf+RMlHYWEIaRddjXgWSijEDxF/f4+v2tsXKPAIC
MHL7/WBXxkFkdGd3cP8qxxHn3DVFgc7c5vHqcSzal5e6WzXavahRq6wXH4PLoJb56vBWMFfI+0tV
IwNsFJzky3OAfk3Dd2OTX7dh7uFFXHjAiMQFK95vFZ5hO8S8tE/0SYE/LFTaTx0yDlSjCXz70VtM
ujR3Aq34zNnzDy+JSao8LmBVNz/I5ThOPTXQfoyu3tR+X0mU1OrNnMVH9sHr0qJf4e++zN+xEGqR
00leb9+7KfeU7NC+i6s6SmnSXiFFTzelYXw0pCNLEbGzLXzdxr+Y3YDj/cClXBqkCZJ6lLrS2K+U
JmGSq2ZtKZS34GTedGJIfRlDuLOxEw+uvasZPg2JfTPmI6k5Mjy/GFSzrU0a9ZyEXBO+VjUi49gr
GgUJGIx4jw9GPginSzpMvr7tYka90wo++xoKnTQAnpLNTlyu9dozgFlAIZouKA9pynxmGRBt3TQ0
ZjRyYcVp/K/55/X3aKprMIEWxy6KxO3uHNW7SGSSOh/BEA/TqG30CjDSuvK0VncNJ/P1S92JVo45
sDlRbx15PEVjhusGTtNWuj6S89cudAQ10h52Elm2MMS/8dhQgxL/fJwZj/bVnye6INaNG7Pjfn4S
0cHedCRIyDQsN7Y/AaTBpHq5HBegh+NA2yu/9HaoFLL2AFW1aJfaAzpcFE3cGdrZbBAQlTWTMtjc
P1JX4fZd7fzBGYVyIxHRBuAUUlEXmZ9MXRWMqOm8RWq42BCkRAY0R6TmvIuXsCWRk9fToqnWreSb
Be8FRc4Xlp6NF48A5MhXho8qFsqO76b0TJRB1jvIbkQgZoigb9ykInu9qZ6SY+ZldojpFOQboC2S
rxs9uc+krx33+WXueGs3RLBo3RF6EavavnHNiFr/5Jma2wBTAxzbF9RWx5IjH5hXX96+y5LzlUpt
vu3C/MDGTWxVGBOm698EcdADijx/YhtfwX7Tn9KKzd04A6Qg2udEdDTbr/sFa4uyehigXg+VgQdf
ubJadczlmAX/ZAURqQOg/eyH1LEE+0bEmmVij32mGywKnRb6D38aT3YxInD/MHZmnN38QaBzhdte
N4xPwzseOxUbRiH5fbZVQT194RAiPo1+lZhbvuOxEwTg6foNnRw8se/AEl9Zb4E1sLq5xKFh/6dW
Oajp5rhOo1Wkpmrze5Ur36twNx+uw8uVm6IGdFd9kVPPO6pQ4FZDwb1a003ChpVFujGkAnaulsS5
nPiEVYYMS7I+ss6dkVsHd1MndvckyxrXCKjmuPU9bpEH9OI5KRlgo2jNuRTPJe+3wQsfEDJSq0a8
lA0SYQhe+YTCAwHhvDMIEzAe0rjv/NOSOL/lry81XGU6vPS75hIwBljqhpOcQn/VWn8jHtPQjwg9
97ZKewk+NGSZsWUAqFQHUZVdRCDExqZpPTBdqa5bLubDdfiVrAwerhVhcW5zNcAI/3drtKUy/KAB
7OykSffQVye23w/1qM9Apwani7Mj+jKxD9es0E9HRbg1nKZJPN8vwUbE4GbGzdT/ioxHjC0gvspz
jFQliKgrMIMKBEzTj6ZafsPdBoinlv/9WZ/S5NEXjL++iB1E35tmobybVWmuqK23Jv4VFB5j3/4f
e5WH7wMiyyjrhm2jixabiqxQrG23NwvjO7pfUKxnUjjvyQgJg/2VkoCMX/B5055O4aVMtlqzSR1r
3wSA38tZprPTxLqLwLXuLf1vvGOApi4KRRSVgfnAgqmSxUHb95cTeICv4uBBrpbLDOVccuJ76M9T
tsa5/loePNWU6/SKnOoW+8FPW5ZvTj+CJheCJXKBgj2r2Zd7UzdSyHMtXG17P+Sgr5urxlrL80td
rP9D8PVBoqCGb1fKkiCFZAaAlBvZ56WkMCQuIsAYIe6kfPBhUGCcw1K8D5tGFRNwVl5/5My29N46
jJswH9e6axHdYZHimDTJ2NFWxIIB+ULlZSfxBzU+Xi/UH9kX1jG5XLNSt7TS+lputPn7p75G24Bb
tNWQg0gjDNjCt384SPgy5HRt8lI0GjFth4NYFzZjyxCOYC/mFyIb+zdkCV1dKx9OHdA3XhrNq3Xe
ggDJKmnQEwAfqsnmncMSfl6d7gPSpCnigvFFn3SKp3o14OMPxGhKKEN7LiCtYTe34Q/0P5eYPsnz
pzA8YauUudXX5KiuNJm5uFTtfrE3mmQlWOOpfc2jG/AjhyCDJfYcqNEjW3iIFp3YHhLbwtIoz9In
Gq2yQW/G6NVS5DaVjVAVt2nJQ7z/N6vMIRJagw59bHUZbSZh5vdP4D0HdqPzGOIj7jmN6c2mJHGT
an5X/scJNML+v4PXSRqc8yN7diodKsry3AXeufOib/Qw6gq5MfPOeMsqhUD/EmDxHTdYhBHG35lT
TKCY4DBHnfmSimgnswL2UPzcJi2Cdh15gTHI/HI1DNDgIg7idA5c8LGX2DgFI5uw3qOHYf0PtQ/Z
fI0IHsz7SnpZgWxkHxEXG8mG+Vszx12M8T6zlCdaaSiR4pDhuazm9P19cE2f+qqtzjdsUj5XiCuT
oZ/rNvJDpGkU+yOWRBaJ+WEG9q9VKch2L8lrqdXnLh+0dOH8mopgRoNkJbW62TBbXEjc18kf1DNR
hKCiTjuo2pl4vt2Nzf0Q3RV6lXnLBjbboWiDIQsRX3CF3L7suWn8ie8oW9eblawMULQ4vbblMJBq
kcn0+rEiTxau8zMgCaCKbVPDOfM+Rwv3I/U/rD92Mt27iQGOz7ais5gWC/eUGAScpeewXRM5NtkS
3Th9+D2+VZCioLxSa5y6ibEl6qxMzl/fPtbnYG3boVzHHghrBTXY4TYRS0Frb2nBD7GiTKbKTe1C
uDXqj7+GVDiWdeHqF46fZ+Ob6/pwjWsY66aAeWeMEMS+jv20jVRLI5lsurfAkNiWYBgUjrpFI9FL
hthgsxftJCytH/MXtB00xJQY1HXCcvYa0vOvYxH1D/CxrBgG229BiqsJI6D+6KCTKKapctQjT8tB
LdyVmmx9maS8gQISvcnzYNxStwxzYydMpCXTl+a9V/EUd8AjlDoOSFNkt2gLyr5rIgc2Nu5VOH6d
qUnwtVzF6vtB1sjVPYUSfv1lmS5ts3jTjvgOKeNmjn4AlFedeiVl/pi+daeWUmSIQol1R3HjLdxz
FcuodRqZllFHZ+XzExsPFxRNPRGAj/+tkA553aC00eqhSKhdJADfUGmOEmMtzdG9dH79yvapm9xa
2YZzLPinpm9bmixMeWfrS6v50WTCf9rcXvf9RMnP+SXT/hIBFKVwx/6TLgcVgASmbL/IyMSUS8nO
FkY/FSe2RjBuK7j6nZb/NgckfBla06llaYuwCvdHChsbFfBHFZe6+tWLrd4o/98Owlwii0m3aEzF
sN9MeSt/tdilgWEnAYRShK3ZpR3l+vyocRBG7/SeahB2yQ87Yc3uFXEn+QFHpNvd//gagf4Q9Men
+5lf+vCv3Negr/m8Dqp133iVM5/BSdrGOzAHvc4V9OOcaAeaIywxVqdU2Db0y07P/3uHJjkYS9Cp
NMFrNQ8HM/R1uWYEj9mS0dVaAXGnlhVCo78SqzuAJG4HcMiN2LavuDvaW/V5QIUvS1pVeT+S86qR
aQSMSNFIWSu7BcxoU+G3RAZVKOYEq1GA0OYWJhgKYOgyl4ZE4L4Y++1wSqLNVrX3+faNQiTnDDhK
FNmFO289OqRVE0kl2yXsuqgK/adLhtwnO5dAZ7zbzMaKXw9U3s/TdgBzokAvt8UZjpRd4O/qT05Z
P9EIRr4m9lo9R8YZ+MmjbQVyFkyh5ASDdLPiJDuQC7OJCfahx2WMER9Q8e3LP+cDKMFZEQcxy3a5
Ya3YqKrQYzATG79pqpQ4T0sQgmWpTSRUiJkRInKsuSNVJPXfcalrH6+QoRhhA0eOA+sa+ONtjakb
0l+VKy5Bd5Q63lncWxl0LEG+JuyT2cvANyhJutz56klQ2LMFuH/nf5IhaGKDkmkfCU378ulY3sXn
cLbJ7awfzFac8jwXJDCslB8Ev3DraWIqP7Zo1XR/tuMGfqIRZFDE15QaHU35qbs+zzdOs2hT1LIM
IdKl8XxREKUzy3aLjlS7N97BRhKUc0BZvuWNYbAjyigfTSpJ/7xOO4hsMTIDFk+r4gCQIHPF/W89
WKwvqSBw1uognCHXQF5b7xm9a+NcWZ6FY1MElWbKROmeWcqHDxPLfdSZhaHMtcjIDK87dU8ra79A
ENnPGF3j8FR4IZPB4ln29G2GQ4cu113PRN+hdqfplp13rVuvavvKMiz4Czuud5W3s8N76xd4e4Q7
oCGVRaU7PrnNOyEb2UjFSLL5T0NgrJdyZnjQTXVqNU4RdkShiEUKn/UOXP8tUD0x6lzEnLkCADWZ
Is8n2S12pxeljR3QjRCWWEOLtqjYKfIgah6p3YtTK2ApotLn/e/trblJshEUyvQ+im2Dnma4+gX6
9Rh0JbVumVRbN/sL/6qvGLdBsFlBVXXeKGR6QTkFZ3p6yfydMCQ3bTgdiBF7y3b/JG/AXNOKewCI
3VO/skR/utmDz+EvhmtTwX/FU7GSX4Xd1EfCRfbyAKgO0QBVCVagD9vgjJR8NR19UYN2835Ikf/1
xCtcpvBWkx4HqZ1Me4MV4iiEa/RXMDd6Mt9czOBSSCwqDO69is5yz/bUFdiVvtR/pjvjy1xXDbn4
IG7ERW13ak5RXzEWckLjP+y/bKa0eVkh88tpld4MRJdgwTzG3dZpZLedpbd0+/DzWokgrDB9Xm9J
D+JOvAqSDephthlfIQFXoN0j7usM/+DhQmRDw4g6ee0cxD2ZKAY5WQZ1Xo86LTlhywq716WUQ5FA
VkzD04s77CPiF11HhAz8bJI1WB6rw+Xid9lN2bFSb22LcmDihu0mSOkMwpzY63jXWknijCvllMWK
D9/qO1B2TLwGZOziDT+zTEjmcfNR+0Im4rUiDES/IZTwZSktZKm24xj309Pxmd1t3IjzoNm8PPZX
BjPbCFU/523qoGWgKVp/oDeuSbIjsxPraiyzWa1PyJVnKquR7somgTHUNDSKqbntIXEkI5ATzznZ
ezf1apcByROlsNzZIpbIa377BhNl2NMTxYd6P5uk5qbITtKzvbMbr1ch97kAN3TrNjg9C9MMA8jC
zLhN5fGFxkBzAjfghMKLQObvbFNjRtLOO3eparv9pUdIVVW3bA2/YwzrK3FX0hYZlZ47uZS9yIvB
uzNWLtr7kiis8UOOPlHPbMWU3ezNpu8sCsXT7t/nKr2xYnFsyVcH4JitIo8txsclCvZYzmbp/de+
B+rPt9e/jpttmd3biUN7/BdFf7aw5tsNFpRurEyFl5wo1//uaCsPAcrKf0UWKoTQpuH/uMtXWemB
I+EAkMK7AEo3b3UierCPru+k0JEg92MY2Dwv/5ktuIUidZrRwmCllRGxWLIKXb9EVD7f4Fg1LWoY
KlaFFRriAkAoG2gfK1Ww0gmxIaUmAQwFja4RcoVOCajkmkkyeKzllv9vE1MY1nsC+bNPd4vqdzpS
8LlFrYZsqZWtRH9bOd/1oTLNe8KbXYTbqJSrShcPX8xunvJaUcwVAbh3eu4xI83puuDPl8zv18Jj
E8jRsB4GP9lMeC3kSTpb2zH1iCXR4zf5D1jEn39rnRYzPqhdw8Nu/qqaRVvdGLY0GtV7OH+Sdftv
pgXUnv+5et/P7SVswGUOPS09pDIjvcw7G9yjdx8l98OYLgOerzQ4NVVUsyo7mJ7dRKsjDmRiT8eu
CSrHt1OiA2TQFPIouav4Iot5fiqJkm6uAw4jC04D6gr5DNxmVItRFR3oqJnUYgWu2lzGoL9dDf0p
5pSKREgaz+oYVHs5yTCxkM1Te2e9sofvUnJqNWOMSEL6mJ5d8FHogz6Vf4iUc8mRiV948UwZBY73
NVsO6KtX+4aXtCruZzu/puP7TUMhlXgBmUKL26kWxDxUuW02ja5xOp/AYohq8mQYTyPNlmydFfus
K6K9c6U5QGRjF6tU9qyfhoUfan61hntXwqtjSvW0hfbtit+om8xreyGJahAw+jVSnhN5xxAaef7H
nLVJwusfSUDUhNthbC6HK4beWugh7Y3ZIadMgBw0gxjpYWN/poH9irxK8WS28/4RHqMJ2u31oaQI
0z4maeJYG+GOiPMtG4KwM2CqytXgWoDeyEuOxbszLEhtii3gnLgMZdBBaI5EdbToukxTqvdtQ/1z
HMtQpGHb9oJcQzdNyzFwhtUYNzcpmUneb0OcEgXJ17C37KH0ZTH2EMZaH+Z6cGrlljnxNuzuUdM4
bDahV3+ffGy02vzoYJO1+3u5UzKZ/PQ+mPR8TxI5I+pKlkK2z3cMCnjtCwqBHXRqurQZiEtD858k
UPMYYXBVX0Z3b1MHK5N2Vvj2mLGbC+XxG5k5jQ8PZclGcIfFtqtlpj7PNk/22fELq49MmCFEVW4Q
uKMHFhccBuBOX5otHG2If1kdP/fpHdGb68rS+8Ab9gq8aPeZqECd2X672kT1UKceHnHL+1a7G2Vm
rQZX1oGGkPDwTMuRd3HvY/lYYIOYH5YlRZkBH4C4c9EXZ07i/R2S/19ZBlIvSoV7kSxII3DjB8JX
GdPEzkSk0wMdCNndu1A3QiTCrcvvhDW4bhfkVGNP9Tfq9vaS8BH07wLC2GnBZ5/y9tDK82V78amD
pTMhdAH3nP1OYDdqhCMwVmYd1kwf24B643ZKt6OgAp9Ps7s18+/UYlJWrZo6qVgwwurq7DHEu4xw
5Xwc72W9evJEAFmwEO58QhaHFzz2hYKasUK3YVS2sQrc8nR7O+HHUF32OR7rBK16gM0FUGi7wXc4
ys5Ck6khTj8f7DhOqui0uWpNv8LBefSDTqHwHu7RFW2aPLSAkb6GXmNWxPmXqmKB0ptO0+rjmO7a
MR0fv9d0rkMnpoekKEXL6BIbBJDmQw+wLPj/MNR+R7Kh3Y6tS5ZWi2DjSjGIS6U5/NA65v3Zju0D
Zcaz5+JTOeM32dsfEK8XsWQjP9HQYLbq8EfmbsX6AtXPRoEIWyXqxH9ssCNZZiCpwJdkcjW9sYVr
0HOGTafvNZufxuAm8EzWtPwKbc3qNrhe8aFdijcXdvywtci+4z4uBBSDKgEOTDyfWRqYx47I5MsW
TZvkv7/rf4FOHPdgjXfWCTJvXlIOpRwXlxcG7igUGSQeTglH7C2kd3Bg/OliOrpTKljuyJoGhYYb
sLYHA4JqDAP9eQZ70QwZ/d+A9jpkA9fbjivAAhK0NOIRcAAmi7bnDMVbd+LVNQZ8YihB0DhBuGkE
oDtiqvQR6wzu0WLUw0NfE/YVhAqLRQmU+T7yeC6PCfTKMdOdVcubw2lFrORw7nxR5fFwUNagIIWi
SbkJtFP1e86EFh0fs+P9WI4sAZQCw3N4RAYkmz48VrEU4kNQJyRbi3eG7ED6XeEuYw/X8CKAxGVt
qzUgx8gDbaBEqwkyV7g+nm9Y2MFE4uS8YyFjslgp98cIb4tew60lvvO9UI3xfb3fHhJXsZm9aoKG
q6xKqW8ua51MgBOLFB0P7WE/5mgCi3rQCqfuRfhya1ESJYpLF/XpZNZqvEEO/R5GzT+h/G35AzHS
MVh+ewvhVhDkLDy3Vb1KAHxF4kOickdhhQ86Qeiroy+HNk4qsIOgZoO2sKl5+mT2fv54g510Wh6x
neqSRs9dlzHkdho9zNKM1yfvP7o7zGEI2gxz02zHa+eKyEdaFa7GJ9YG+N8GuMjJuKbYf4xzaBZp
zjXYIatJaIDC419rjhzdhqYywxZ39sD6x65FfGRislWASLHfU4XNak1c14c5LBDGh+zD9B2Ez4b1
+FngNEGc0IDT6ezMSqBvhNLuhga3EMgLWNpWd00XLA6WzfQATjMsjXz0sJCo+wNT02vGMNpd7Hwv
NsfSgEqJN1gvBqMinstleR3GArVJ5zloiphK3qeMAZQo+8JZMvUwG4CxS6D5FWOSWVBSiKyF8kOZ
+ao1WUdcIRgU0NpWJ3XEFn2ZSXFWrkmmckCsgCQXORYwdI3Sb80JrOfR8Nb2ElUFmA6l/Zh+g6xQ
s0irwbo/k+yeI7bMyCMvNurD7FQPVG/CmdrgvrPpQ0nw97ZTkXIzTHaTGr7mSH20iFQvZ7bY9OHh
IuxYaeuBVc8xpwet5SW9uUcHhqA2Lg+9OAIA7ut3TbjLIzPQ/DOXgcxzBnfvSxO2Ms9YG/o7uhED
/wxlcU1I9doZ3Kcnpm944q2ShHeo8xo+PPri/QtnVBHhooaw3fEBBCY5kXNuwrm2PHFiNh78hW69
yHmbZgfs+nrcH+5T17kHqAzq/cso3PZ6bb5PWSnzR4bPS5PXGCgFW0OiARmI34EIzstXZit9W+FG
Gx7xKryHgvdi9u9NyTR5dhf+tiWlDtwE8A/tDw2wlo5XSkfajduoov/kwnDRXPpzCaDDpsEzzujF
Tnz+6rVgUW8P3VngXcfa9LYlVAmeZiK2FYCJaU94RYEfe0KvNO6ZYCGL9qS4oYASDdRPqsNDLXPo
bwz6L7kxQkMvA6d5vM9kzKMlbP2Ip1pAL+Yn5nRS2t3csfvclC54sSeg1TK71Y4mzj1pq8gFvSaT
35Ls++d3CxatdSeHO2nSY+PXVMX3FKOvBv8EC9dukY8G/tRChIK3yTQMyj8e5XTD82IEAZPXSdw7
/qRjXL9WaSsvALTuyAOQ7IAQDKYvHKb4jmt25fN5/g2pQHcoUsh/pG2GoeUmWnDAugeakSaySKJ1
isQg21epWz5/4hU/6B0J/y2gGRXTAUr7cKGJeanHB54+9fe6CO0KYWhkIGmWRcvMSh5OW9pXED/R
PCfoJj2/ygqQuJqi5BzQ5SOnJzEOpxToYuCVnAGOFWy+oLNIrPgGGxVnr5uJFCNEZojP9OL3AhM3
yyfRogAe1tIBx5hKEQ4C5MmFKi2EjEBtuBf0IPkTwba9aVZonldcKcKMkO+9TZBSCRVHsR8OM0Ds
SDH7xFNuxP4Q1ZQIqHx73Yh6uevLNvzlgc8S19zLLJdo/jQuXAqF2aZ6y/OsiNk29Ek8QxIoRbW/
3Yyw+js2lY2vl/De56mjz8pI9+CGXrS014xVLPWHFnLo1F5KkYuhCcOAVT/7IK4MS2nvOrt+rB4w
smMdf2iWmucm39apKso95g0OnjnVyJmiT1xv4ibCG26f7y4FtUD2s9yj58A2Ng/vLZcfrBcujWtE
1moOeTRSK3s2lZTfLgtPoWTmlZqFEYmAAeUGYzw7KjNAsr3VaPsXeia/PnWHmrWPm+RSGcDPnDsH
/W4rnPe2vZSsw5GaC5/rjZ/d+2N2xASNvYqxPaAv/9NgbmcoMUFimlgnTzYUCYJjlbzkuW4b2d3o
BU8/wxhdH2mZ5rtYlgQXTXsqYehDnqKZIBd3E8jZrJ8p9W/9/Q60krZQMapofEakbIw1Hq/FWsPS
zQvtMyV43WzY4oDmIARC8Q51ZSY6ji+vJY2GBQteK2ss9Trnex/5dsmDjbsQJIGYuJJDvT4NG+s1
L7HoAEVr//O2JANhOIAfUk8fSUZgdbuWZhe7P24MOH0XDyQ7k1pmJwWrDpbd/AiuseUqeZk4MJSy
t95cppDiE7+aPY0C2h7ymazHGRJzfM8yczAdGF1AhB+UbnmjoK+CvkSDtdOucsKmYLsyfFqJa865
tcOzzMzUZjKaUaaSZx3FDggDFvrDZcIiG+0IJ1763gA1hoDDo2YVeOt7WQ/ZEW+sOxridMoHbxTK
CWbF73FhC2H39Eh/Qf3AbMeTrf2B2DaYYo0C4zpa5Vqdz4NMc3A49RRzqe6TGfclkg3R2BGShXFs
Bj4o8hlt48/CucdkvvPe2NLb+xoj734uu1spRPhf/qZj28gIjHbZPjc81lb5XaxG4FQi/7T6JHLs
OypuDjuAMBAl5i25JPbkDeqv0jSTcgldrU5R+qqZ7QdXwdQIaZg78CB6U+20tJb/x33h5122x3wf
flgTNeojfY0FE5ihcfDPBeYpoQIq1eJNVuRWpANiJ3YuYBQwmPTyNx85+dZiYSqXmuTFsFiHhnpM
ABTThSxz8K24NEWObxr92R4948YGGBaholAvn2Z4EHzhJzm9QFXEkA8G5M4dPyn/tchE/HmbZG+Z
fZ9OMANdvevj3MQ0yFf+Juvl6jtPTOVy2Eaf/fnUqetXHGINvnJRW/NbdVC5QjSyM/TECmI7Cu4x
FwLZmNs0nFBJdVsnKSMC7r36Ftammcr/vqKBKEMrVpONVDp3bMojhOY1whPKwMfIQo5WJ1QkN5zD
mdF8W4mc47A1tlR7kdPpzx1m0MpBEhsqLp52G+Y2zNc1/XRVblZtjlN4wXLcdwx0Guf92xIDhv43
B93BbsG5dPR3LHwQgA1wLldpjmn4YnAQrzCgG9GyhBCpxQMWCCskLh0AQ1TR2gCE2gbYKC5nzXqZ
dX0lOBsNACFX6Y/NZQwh+Nd281N+hOw1nxQzy/KIz/M401fgcyE1XU80QTeLTPA+wXeE3jADuycU
wyp8fTVZTit7FmT7eot/Wker6L8s11p2sM4w/yJYr2YqSIy9rROSBXAtA42st1zOPdVYJRfNiuM2
rimJWAvfs4BUP53akVZX9gTBfQgxPn7id0fgnTipgNaN2hLhh5YOff6pG1jvdLUvtgJdGsDVVvvt
noNO2JedS3NohbBnk0pUoLF83VAHrT5Yi5vJ0jbmgnwV+i1tBDiCbS8xPyFC1/b6rbnrJz87n0Or
XrCjhcukh/AaVzWIEypkIZsob4IjdThP1EeO9WaUmkljEkj2YzaBxXUCeADvdBLb6n0niX5xyF0u
q3BZFsNhKK0ZZ7lxMnxwDigapg8C10752Pnoj2Z4D5Z8wf2F+/xZhb30dmdFQjlsSVNAzHJLlJ+H
AWU2Wqkw0S0kmO7apQm0BWlxnUs5LjkQFADLQGT5d836UhlxniwlBtYhXEHZufzOCA8enrWPLZyD
qLe9yggoqfn6JJQqznscbfCEkVs93AVoMMy1ETPIKdeSwIUZzaRESGmFQOCx1l26oqk6H8pKtufN
w58cxxbNdvPg/53DHSOrCkw35tgHzXtawBQAtOaTo2LPcDTM2Lc2p1io4qIAhjezNj0J8S3hC4yY
lgLv4HjUR8I/gK3LQkEC6cpPdtfjGIawSINI1Fn6NQFAq2tEoHJ/ABv46/wwhTS/MhCenJaqoTdm
Ur55P/Z2+m9hwFNceQOcP2cTVdaVeFUhKUEzh2u4lT3Ax1O3Hl3KPdlRaf7Ie4I1dMaAHRghNHqs
5LcwZojCkYyWSJY+SxxMIXgOwMpAF+QufpD/IAcI6vgxx79bkMbxE5c4KU7l8jMyBL5zUpcRE1aQ
N/z5HaqRdnaH22ETBUsYs1VHWR3vbonXqlMKuN5V6I3IIxkmxdQKskOJw9/4K0Bh8R+BeNvpACkj
NC1oQq9EABocNrWeBJ2e2Lz65YrBDB48IINfe7hdPXWLeS8lWPazNp98LC79c9N4poZ9wfEpzyrZ
ewllzFfHut7/6iV6FZNSeSkxWhKEIlOd/FztCm3cOSMqM/Qddo17X1ihd/rCrmfUpuKTyximONHK
KhYC0gSagKWDPXxAv/4YPM1+q9bmSaSutzB8DC4pvvUws7M6+4QnKcj7Unz4UQSOkKb1D7mGSH46
/jl4Xd1tZUvq47+NuZMZkgSU+4Ai/cXGlWEv6HdsSaUw7Ju5mxlY93WkxymsmPm2sAtKLnU4Wppm
GxQ6gB/GoKv/BS+5skf8kOQ7isGROJDYOiY/Cj+LuJs7kEwGR0uzKnXvjf5bw3f9FKopcPmyERIm
VLMw1nFKHhjyBu7MPq/YuYnfEcMFWG1DA+oP+iXTxO4Lu/a0GG1IyNnNPi3UZ8LRE7QVLtf6icRY
CKet3rsWL3sZLOmuRHRObxL2c2MazJoVrhN7VNViAvmEOcZM5wnghvqs78VIJg02gYACW3fPOsJN
Ho+bvAaYekD38UFNhta46Ctr/zQmIWdfggwe0XS+64Zf4ug77yoBr4b34ButplqTZL6Wi7dO4GGc
8YIOg82j4rx6xcRcImDgZWNRQU44+67CGzsNj+voCwRmpw3X6AaqiHSKoAnh4imL73tz6ZJzTX6j
1oqWBVAN/mb0oMOc+3XXDYZb7vFYE+lzx2KL79kJvxKTElZoOE47LkUgd4S+P1VLpoJDc4GlJwvi
4xiPJklY0TR2/Dtnmao33BDP0OF8WVqABgUOGFKkweUNfg1dl6Rh7MK/f3HDTG5d6AhqhUIOoIrR
BZYgwRs5RbY4xBZ1n+pDlMjW/SSQWcy+p1DdkT9owcHve8jbLj9gO0+8xm2CNpGYMpIHDl+y5dQw
Q+UHQ0ewv5JIY6CwgELhyZXMBZtABHSGJEswWEaXSZoHtbHggWpO+x0JKGPIX3A5h5Q+laqQvDH2
VOqScNgxJuTmQyrkYqxpCxM5/O1E1ZcAUrAtUscYjTD3VPa6ekHAs9hrPJ/2H8xL5rE1JdmABo5S
Qgb3Ouv9BCMOvDqcyF5l3errjsYMRqOKYSMIVqBuIdvsMSR0zKmRlQPEvLJXDyzSffF8WtFAaYLk
abFkNPgRNktNkFN7dzx1o6LGtOmvvZKs/yc/exl8bJHHD5QBm6FAhZ8O49Ae+Q5aVKGHy0Asfzwd
IUOQjEGgS2Z4DWJD8eLDCjy27v7cqvg9cw6A8HLVijPGAlj2DdAe1bulNyhAfdXlKpzN4mJ1LrVe
Jm3xZaaE25ta+Ay0Kd4C65VM5PBfPi20ei36b06wAPTLLWx+QjsSxcAdEcBlvzZeF4KShBhOKDX4
3OjhPnDuxepFEUwNqQcg5oBDTdb1lZdycGj+ekp9cm5hF3FirofKpaVHst2MxPudTbBhNsmOUXbA
sOAqE0/hVM46YZp6KCMMvH7VKqSz/Dghuo4UYPOiXoeE6RfVf/xdpiq/6oGKUovmCDQkpHjluB1c
7ietfkIBc/RzFheU3tMnNoXyiiT2iSPl+gHMspS72dIr9E6lFZzjC5d7xbOHkZGoc1CWsCH7szSQ
kcOhFyD7kkrlJMtPrRK0CDEC7V6vRB4KtuHMn7tMm/ikAf8RebYxX79EvKE6iyME+Ntz9gdbR96y
GjK84P4exm45DguIonwYfQFzLmscLh319bp9SL+0GoUlumf+QMUj8iYZliIl5YdD5Q9mAilZq/hi
1BriqJFFNDK9XlkuimzzclSV7hke2HDhOXrAXlyiFy+d1zBkD4XycJ9CodUQT4amYBeVXLmkiAg0
tcjPsHx1fb+ExjBf2/bjmzdyWleeXhE03y/wDqzq0WiVqC+sKHFSSFrmw5eXZJljbdOJ9ipe1Tg8
w+zJa7/HTJQxkneeg0FBAn845mRXahE4WZ4fNMlwFJv6B6uw1W2YiRUvFDxnVEydmm5dUQtkr1t+
2HVVJzLimVGgxht1dAyTgh+xhmFffCj7aTxXt4Wr+Emrtu5PZubprloWTzvEfbDwxOOft1D8pRas
mTay8LFMPGLRBSIanFqGE7UVBxFyAfw0IpYmNkFkWCwfR/i/G5FKPmkTAltA7lb574C2c5E67bDf
3g4HHPOtJnaAf6JY5xaPmPikSnoZpkBY0f+/j7sv8z3nprFyvIGSes1blg7Yt6iYycUf6te7XGFI
CQyVwJ7drASSaE7Yh3xM5O6PPYUs6waCFcHgneaZe0WjuZCJUB/osFfi7sscqxJWjL6V92EEGNsw
RBYPBB47Zou+Q3H/usb5U2uc0EEgx+ZojkefGL2MNTBoShGl/R/lcmIRE9Qmoxlo1B44D33Feplv
43tkS6lDMPzvEgi3l2RciWZIynsD3mbtK6bpgzWDSD+8RaX2ZigJqyrMt8kFOy3foiK5ygUTi1eu
r181oHrGi5TKvvoFQvh1NU6+fAxojt6iexJzhFFU4HtTEQwFxY7dofy2N0u8KeYxnp/m3JhenOE2
K/dKxlYsbESv2lTilJDXXXWjQDtW7JZ9KGsa/cgb0iefl40LiDnWBxq7qy2I7SmQrmA7gmifqC9C
tDRsrquYJoGm+Ju5fUO/6aeqGEYwDVYk1jAEtQYzMWBOmGmcxpHcWzYa5Ix95+6Tn+DpSL+8sIj4
46a7G5uZZgOH32a3MlxWdpzUOkd1fnWviJlJJtI8iTXhbdpZmuPsRry7DF0XJBLe28tD/5VDrRaI
iqLKRPkJahIzqqksEX+Uasn2DyH9pwfiFtRehWnzoD/d13OcpSuDdYkTIP9I9k5De3i2/CmXdH9t
DGAsKGJBuC9wPh8Z9VWxEOTeQAFzN8r8PU8/Ny7pGyKoUBWKRaVfpv/HjvcqiBwcPuUXCc19tuyk
cgtRmlm7ayv8/6H8K/tudgl2znkL4EUeOTzK9ohJHLtizS8eD8FTM3Erq5vwt0uLTwyaDFFt699/
QNSYFri+XU0ramiraKidc0h506tD7VChjwmo+z7vCeY0XywNVKuTNpBDzDiSWT12SjNF47FVtQZo
W4u9XcrebGWGkxkD6tSWgBxLsDiz2eaIfFGz40ukGrvSg210DpJxuqhPcUHbShwkw8TUBHGrlg1g
dkuZeAadCs4kA+PmdqbZLpgqNFvHcFbhtZegvcEtC8y0px+WgiY2fF7OnUOJyjmnxEspbNFomziK
u3vF2yvX36PRojOeQUr+FbSyW3tNxsdwvrD4hD6US/YYSdSxi7JXSk3xKWKKncB7icQJm9ilip1A
+HHSk3VTqftmdY5PdMoEpgspVMlLIkkIgxxs7Vc564qdnWBNJeV2x2mom7TQli9BILiDgoiBc/vT
FR3/PXSc98rKkDs/S2HslWlZnjgbo8+Y9Lry+xlJGxaI/UN0knTQZAlEOlYWLPOvmgrUmJ23KlNC
+WoZjuyjHFFeBN+nsKg7f3LCwldXxmiQTOJbcxBl1yJle0ZEcBcQjA1WWk4ero1gWE0l0lk+VSMY
Vlpbd2ZGRdlkmZryyFa/p71UxuBk4Adws08hKOewZCvAgrdEJohgXs7jGST8OppOo9TkHZ3j/93+
h9IS8Jbu4RYW98ylJSXBvnLxdUL7EkphsBhPWGiss3AouSWKGTGQbcVDi1f/a669b3W9Rny/1eCA
aJ+emeo2GNHKqhzOn+leb7abAvc+Xnb0wOpnlmmfhlkLg886q02Jj08j7ZRWkpv2Drn9cnng78oD
dOyrHPPobRxhuNB8ftK5Cqj4c63CyYboBaZ9ex2qunPtrqxdxH9gX3T3srFOOzI5Imow9W7p97Ax
w86NY+D7d62zns72+qJtHsBytdhR3O9iYhzz0D1x0QllNZvPDEMxcJEFdxwWyVw4FzyaK1k1vgRq
OVbs+Zjlcwd5I4NOQokVdtdohQF4ayKOGFdRl+HPvRFe+NxVMVBeZElbSFWNIALFzS0dY9GMnZFT
xPkxAQyX4TLJ+hS6Sw3HH1eZpyvwZyspGaJG3oBLQwO0itUaAGA/iD5JZJ7Y//mrS9j/ZSThA3Ec
QBJe9/IHZ/CMn8vtbLHF9D6EavSd1kmV4Yp2+cMGqXexjOS4QecVv9svKjVZOs7XDWsoI/MqRGb3
VY+ejhsr0l8pKBpnFQZL4oXcTaDWE3WX06ZaW47yg+Ji6xAma/2dh9rcp0DDrQ5zX2O5nGlc2tCQ
RNCJ2QKUe+4a21yaYQrreHcYKwwOTpPlT47IShptBKQDdvT9s4mM06o/X8ozgwPzS1DKe9E/Flm0
bxzDD4Qkf0tjxtqcNXmM25ZzIczqyYQIr93U2W0WxYCGTZqmFbvqKe5HEMRNBdEnFwCQ05sx/SeX
6CzOX+XvNUqRItdOUvdBYkDyPIpySdMSvLa7aBSgZtu9WiMDd6ETreBwZmpwrX2982QgY2gJn8Uk
ALP1R9+m/8aplEFY+VXsRHrfYh+S9bZg4jTT33sS7acUqnAQpSShfB4kwClY3HATCQ6iPLRRzFPe
SwDCaLuewYlvjcxL+Yx0QkxPfR/ShsUe3nDdCekgMu6kV1oqoNEdaoNY7LibX3hpPO2ykJhlpOiR
/9EvKytJMqjh6x4e7F5ln9JdJ5ftr907vG3dDBlp0WkjlSngQKl8tuaa8HIN9J/RO7wcp1QlgKnW
MvnfJgmHgwL2MMEivCSUW0fZraG3utWWFWVYorISd3VX4Fdr/mBpDZD3LdkNw6WKrOoW8fkLIhzk
zZpxMFsHF+euh5VtVEi3XpOG+FbQNs6ugUYYBEcsne87YFDbjf/bhiSJplOjxTZCHdY65tJ+1Mbc
sOXpMfGID/WLpkfhXuZUSXahhhLMrPbRioR/wm8cI26QyHsSpXE9rbP0PRZEW1959jJp1iVMkSW3
D2CIEtoIz5s2LH5dRvG9c9mV85hXbht8KUSteQBeBXTFZ1wRLnKXzrLATP527ps5FWEFQImdPaa/
fHbxZ9DWrBu5nAU6t13Hub6AhUG+Zz/cnsTgUxheMnX6lU3XQ1XrSdEzQcW8GahBsF1fU6xGM6Rm
8m1uYU20lzspQ6uBEW7BVB44ALHV3dmJ5Kkrq+Xz4fYvw2djR2ViUhVQodBAYFDIlalmpN2fKZ6h
xocnyU7zowFCLgmtl7irFDAcXS88fxEdZ0P7rH0zXxrY02ePofydi4YqGtU37oIn393aT/AApuu4
Eep9w3oLe6uD641BwQS90jw764bRwNs2lwHwPyrBnEI+p7o8+p2ll+hL50fKx2BHajguSD+jtLRS
lna0jkN+ZWuH7Dq9ohF/JhsLq5q1TNrvQiDiQMCFb0U6rzgLiPROBQ0Tt5u9wC+86AztaYtfLw+Z
1h+ejE+a7d7n/hP8Y0cYt/vxZvr+xF5WnTwo3H1yx2u9XMy3zRYfspBWvnYaU7xx6wywlCWwOGWf
+rxx4XAgq0ImBjNS3lktBgL9vhx77B3QFDfAh8GYCB7I9fjhj3LhoQS2mgDCigIJrcqeuagaEenv
eyvy2XBBUf4NcNsIl7pMwkgZoQxXaUpZNT8kQOfPN7FObO8K8mgMdq1NRjoQFRAbNcdq0ZuRX2bD
6Lh702bhxiI3lpuKcbKIXNBR2nLiA7ILA1wztLYuJTwCIIzpJOjfUob6tgEBotqpzZWi1giuqXhQ
AXEHTF5Bm6NB/3Kvmjyi07XViDXnVxZewKzRZyXZKQBpOqQEmpkqkYuHz8lvBE9JTB8pMpEDNyM0
DkGkqZ6BHtCY51EZexgkJR+B6gY7Om8H0L0XYQZnNa9tA9hgcQj9YBhgRvNxq1HBNYMU3CfGTBEe
w+kKEw9PGIvifN8ATfYPxqSxyyKOr/VyV0sVR1zyaKhfjjB/F8R3DbWqYLdCisDNX1iFlEwe8EmB
7FLB2jdNvaZ7CryUPjAi4qxEc4E6gblp2ruECr17bn9oZ2vJL8AEIOgQOj4oe3TsNeZcwHp0iWHP
HDr5kAByR9GXl9li2Veif/v50AJBEMPe0i1Uz/+OJUQ46EbE9FINLEgCll5RDtqTamWU7q1Y4/29
iDnr3XEkH356j8PtiOwWj+sOpK8zpWqpsQY6Cx/NtQjvxrY1OekHiF5KCgqH0HsOfQ90gDNNBWt/
sJrL9Inpv4ztSGwrM4D5zkAX6eOEeXFYuULLpWmQvX9JupZ8xjbo5TCq8QwVzCewKxUBV0hP+L/b
hoXSfPoWDAAxBQXQ2oxRzCAHqC6eDqMFALrL3X8Do1qxxkyZSkZXLaG7quwS/OMDlO3FQGToBysv
463tbwe9FQO4W9mPvaNeEEbu2kCVx+Yllc+CffTfaJUNfNBdYatuMCXXjvSvyY64luNSADmRWwWD
uutAqpW7UGKuxJyAQkshdklhonl5UsHQCR7cp0GE+0YLDYlRX7AL74/dt1FxOdlLM1lEtCCGUKYO
4RQ/wRW2YpPhtwxCmWpdXHz5Dq9g0+WQtq82CRotWI7jttPkxMDUvPBEGRkVMr3pgX7LT2jMDhXF
feWyA5jBGwoGRlTyJOG5MgtBGdK6+C6tRGjfgcMlQ+P6n5pnOyVhOq+RKQyi93egYciR7CIKzzBD
/s8Qm+8XXK/Ru3bjI8qAFLinvX3DjnnTNVZBUjJpyRaVvZqNb5INA4OMZ8BPrHvdoyJmufsrx3r5
WrnQtp6tI4oChnBA7ckVKMLFFsEdULHDRHKll7CGDoZCC+4yHxG3zAiRDHx5sO85IVpxmnNAONW8
S675MunNyQeuT4C5jPgyHmXnsGRu44BrXzx1ey2nI6QQ8fwen6BYdkh6fSia8tli1FE5W6Fljm9G
Q2BH3X0KVAueFx1ChPxtFJT4omGG4/RGdqrQYvcXTZkU5Hc68phQE7hsxrGu4GeynS7wfLjT3gb9
vfdxeOtycJnD6b1ytKXOWuU386+mRW0XkYEmHqlGfYOnjmNT+tyzfhIHPpIVEfWQdjViDU/6eshR
Nt+Y6pCepdzCSQFqWne3qKhhqMVGqfpQpUQeaofG8Qs8mxMQJ3rojRCxnL0Fwfe1p9h3nPPEmear
kGjVcFYlymJm+KJC1NdWKIku2bXntpnp3r3WdqOZHrLbILWYKbQhQNlX+QBDH69ZF5mb8ikKXcwm
TSXm5vw2K3j9732f9P7pyplvaGqd7nlUyXH249FZK2EK9r/V1vwIxbgkwjRj4fWnOAvvx/MzcqzB
KM5/t30t4UA0CHizPLCzlcktVhwUkuqldmvhjT1oY5sUSOhTVKFZu6N5A2JfYb1cA+mSYXunMtRl
j3cowg0nlXzf+QWntmv42YdCqhXbfWf4RaN1jeHtsGESj0kUSNN+ku8/LEE0mStIn19/zwrn2ehL
dN7jqZr8+diWOZnHPzJGQ4wFMB8dxAVcq0AaqY/cFjHwzw1RC4DtFHqj7z74spt7W0j0mRUkMavK
2HZgrrGwO83G7wd7LSRpJ6WLJfqX41ICW+4mCDXPaH977tlBrB7VKODI9dpHcSQdCkYjhtrkXnPZ
YxDToMg6PxUW+wSBDNtrGATcCh/f3d1ffxA3+bl7QCQi47c8uCeXJtUcGWB8fsLD3unhjCxd5U6+
N9Kk7gA7KbUGVfZNXASR++DLVQfg8x3/XQuC6o4BerEjNc33jhQqyIeMFO/v3gMQ7RcPwH+nhrje
xBjr/UP+pyYSdWP2xq/bfYP1BGa36LMdKEEwf3JzRQzi4UU+MkMK7Es+SN8xN1Jsrdev7NaS4VZz
zT6EbHPPgw4+ZklpwndVE2AHnEFlsayO3tQNj3ubLQFkHU06NkbMTgL8yEn74e0CIUbSQ394Un4K
JDfKbxWQTlNinOMcmh3egTKKwO2PULsPRFgP5hHuTw9dM5RxWEN5xtWkLupRt/DqJOOMgCTJ34U7
bgLdaov68lqN2IyVYUrM+XaxCe2P58pYjRnSDTDonnvfu3Ilc0736r9InQTZcR/8RjKxyhkB4kQe
yNtAbTZA3RYvLGSNBdtiaUY3QKJU3P1jWljcaQJl9oinsBMOWydM552n06jMWkvgDzQRWlH7Wcbw
RV5XJNYFik03IIN5lWd8tsaT5OFgF4fazH1xRxn54FMFKM6TeJo6S1bVc95AAmoflmcU7Z6hJeHq
LdfKM0SeIQKLimsYXUlfhrrsGp2lDsdENKTsscggMRt1sGiwtm34XQ5W6oJkOnbc9cGWQLmZ+oKd
7YAb3RCOX7bV/Q37uY8EMYCAMf5tIlB5QUFBWQsBZQUtTFjkN6qR6YozTDl1EcmUwXYzyq1x/ReO
CWK+Wk8bi93wfJ0/et5OpmHMWNrwy5MBuamb0g4yfv4ZoD0+6+VU0TK/1i2TZOPBeRFHUubJ+S6n
CWZU6uEDq8vdvPhx3LwvkwcU4xWsfqnx1sQMSJGj7V53oJgBqwaqMEmBhlmwPE6KM4FQ9yMF26fg
VHP1XFaKk5uTORgAXOKqTtoSkPkaQ83Y3jdPf3QucrQM8oPo/OkxEe4zv4aq0ws9U4xoWjPaRp1S
0B+WIce1Vwed2bc6ykGDBB61ZjE3Wfu4YJTPQa3GToEEMeTaZc6TMM67kk8/VLxg07NkyDJAn14m
Y16PVe+6UmYUZgCmgou49+T5TVG7LqbtjFEPj1Bpy8tfq/lz1IMLu8sTa/Z2kNupzitFoHUMtkK8
/kBJwEI7HO8mq3QiHnm8P6WkOvTj2ml4c2+sHQmwPnQMYXPfw94ZXywoKKHVowvMf5ulHbo+FaE6
q9hokP27wUTIgWnRFxHX5+aEL4/6jnsbKVhkxLQbKP9ZKAwo/aBv3SUw0zPOARDQyg/RpaL9e8bZ
BlwIG9tG48ynEf1Jd/7r6iU7JQ2UAk6F5m2FL5WaSi5cUeVkjhChnKnCcRytXoFV7XqPgS4cjON6
lTtcKVYNuOtgKwDPXKdSMrmVtfg2iZafWCQ5O6+qSdJTKgkLsHZH3FUnT0LVFJWjWKkFYhsDpvDU
2yIbgz+K9J2UEKy0p2Z2GpehBmTrkdBQ/2dJAcCRr7P0R3MHzkWGysu1mhFekcPjEfmGkaA0ZELI
b8AbnaDC7zKTWXHPH2tDZs6DgUa/jIfYnRG60w6oUyDB6k0iXUM8DAvL2Rdw5L+miuTQ2qWQkYZr
31LfnsRDLi8tKsQYZ9gkNkSZhuytCLFOzCtym415S0YNrF8ypfzR6qvuVfq5gmSgLiRocONRiuIN
wEoONJckuCwjzT7vtSBFuC6iNejw7McrbMyhawyx1wSv3lEG4K3y02i8hWWyBkcC0pfq0Jhocn3L
gVj/mriCTLKFtZGVY2i8BNsB8yYxqNli01rth24feJpMEy1o9vgVJMp7+9rRXFPg8JwI83rPtev9
xJPq1eBuCPlVeKXEdbHQ8l2MwoaGrl4Sbrmmf0jdxuyRtH3L0ozAPSzXSfILhJYLiUheACmmKFx8
ULOWO4I1Qf2oDTirIzgkbI1hO83OIH32B7K0K87PfbD+gHgmAC3d4agfeG8wlRLwAnd33i39wGsI
PfNK1aw2Esu6N1kTC5J0zm5OF8X855n4ARfmfKnH41IPwwahqEm6BUPWA54couR/MPMpa6WZtgIM
l58SVxCuncbF2kQNJX9tRdDOxtauVE+wT0DJqXt8aqx3IWbvbh4TyoB4rl/YbjdHkkeVJKiXtKfC
oeYpeodRPxNb+/sdIG454npIN47zJH+tGQn3mEMiadznOLYvCL2pKBQluPX3P8RpJse6yvUmFcG4
ETovNRxo0yKXabn7osLN6k1HjvqyvXDNtNNn3L5eIaYalFTrbt0d97YX/c11KRRfjR9zXkvDBgRO
+UKzn+87A6iplx9UsiPIfYafqpkKBHa/CgxonL8JKjuWpu7Kd+Qfwl/Wkb+tGxAKSkDtbIRERiRP
SdJJtMvVf5eFUocdOmssqvUqgdN1QfCRljF3BhwCU0uRBQivrvKXApYZLFqqExSMrlbm2ckxn/JP
ojkJh67gAz9sIjCawGCaA5+JxYKmBvwC7NTRjHHVaImqv/0+ipv68jZme1UyIHcqbtbp2RssA3iv
MsQx8JSue4BetvxBU54ygtLpkUuwD7OPS40vn+mkkir9zjw1NwqrB/+jcF9kHIBitZ4MMVwjWjm/
QnsyhNmLXRiCLVQ+HO/jd2p0yOnKWTCCZNMlyGytiGcCr3+NVu3qp2/Sx1V9nBCpdHKyg4nGX/cY
HI782lfhN8C1nhKU4r4BPH8oHjz5ZPQbv2Z2xeP6qp/z85AVT7CptUYEUYUMTw4TjY27WD3Di3f2
cFwfjYWUVP3ZXE4tPvoUfIsmZjHREbeBdPntj0UbCvoVrL38v6deuGN31wFgsfjL6yMFOZrxLFEW
pRjIe/vFpA7qqUBQbMDGjwFu1YKlcMVbWr39p11e/gYn+A+NdLiFOowLFjxqwpnguxhxxmh1UnpK
U0+05pUQnpdaDaEdX1MxR8b/VC05xBzC6MQ3SfQrYZ3thmfHk/ko9StWPFq8fpMUKagaByYJz9Er
48RCaC6zK6+KQV6OCN7Irz+KG8k07NXd9xbJGyVWH8AasrDyUinMEVxSTRwi8smrHNUJdE9ueSCR
96OJUrw2HwQ2C2Wl4tr6YE7S/ar0ALLBd7iVKYLM5TLixki4iQPqzLgbMW+xX+yHiWH9engI6vyy
q75xU/+qDfNiBfeE4QDEICi18ilgrh6nWT6XTkt3HGSz/GwUUB0ShJPyszdQv/fZRyCBZ7rEqgTw
sXBNUoNBy/26wjOfsvwoK2K0yPk807bjP828tldutOeGqgo5e8YVbMfTC5FhXsURn8iINRBz/NUh
HsGxfhD9yDIID6B0d9iTGHpuNBRuqewl16QiUdKshQORRCEelnmSgbcCrcPAX78bbaojdIc33csd
g1bQTf3Q0Y2t81wvVguZWOV7ihUyomThQSy+Boh2WDbKsuxCIt5WBIimsrDW2CfBA2TizfQS3aNq
rydp5uNQpdckh828DZba/oaysW72s45vgXQDyuSaJDdYkJyMUZ0DovSPXHR2qRmD1mqNJwXghCpl
nh3O/PAn7OMyQrAg77cTZxNxnf8hNdmv5exhnjDIlImmTO3fC/xkbi0AXXG0Zj1hUDOuIz4c1mzm
1DlnY9JheQ7apQ83yBOVX2dUnd8LLCVU/galdvJutzL2WdvyXjr/t3RiKEhoynGuz2Ob3/4068jB
/YTDYlfJq+cVnsdxHc4gd/GXvt3uwazg/U91uc9MdCdGzB+ym/3M0PvQbn+kUc31w8DczRVD7u+S
lVh6lnAW2gkVRYPGZiWRG3q+7Z/qg2tEjX1RXJ7sJmVJW/Wq2PpVMDaEUM1CbnmuFJpq25BUXQvx
dYROaJXEkLp3L5S48o2YkG7T1tdTsa+N0Ga/AcGtO3TV17HZnAzHDz0bGiKvn2GaUZsvDBA9Mk+M
NBorrfd6doAm/AGFJkRB99V16N3xLedXbawJUpEjE3jbaYgHvu9a1Slg1CagmCAc+uC5KjibT15u
XVoTcURr4ZY+tX2XywDuojesvr0fLl/oL7x6g8hkkWAYL7oRfxtnVubeDIJCkWq48/XiMb4p+N/N
Cg+7d2Lp50cTIKrsFHXMV9bHaMxTL4WdazgwRvQokaF1yyIqF2K2+ep18M4ZEZyUMvJ2oMWNjndA
ZqhkvqsflZyR4nCymGEtr+kDnSxVMaB/3ZIWtoPJHqnfjmymRVUigyXftXH9KWO0M0jrdI5HSBw0
/gl3pQEi2PJ1tJGxCcu9vkruof6m2VjcvWOlFpxVa5vGUjxlEkNJr6KtaRPexc6pKT+Y7LakImSe
Eb68GMJyCiTkjGgW1rucjxfrimcpyO7q4J5Qti0lTS1rNtTtSj9Aw6n4zKrpdzQX5IZduGII3byG
6yay3PCas1L79JAIyi+KTmISht4n/umfHl+QElwqSXhqUqskZu0u1ijxmKq46e8vqpZ/2zJX4Iv0
UGdI2jHB0v6TwjVjIrySMQr8zV0SX5fap9gh5Hdv0V4W4DleCqhAEYb4lxuBlEi2tCKlg7i9J0wl
anHz9IQG04E7jB4wgw7hciMzc8imXJzti+IdflbW9dPakseK+ut6o/Mpz6OA+A9ghJwV8vUKtQ/I
oZwa665aEZ8zc5ZAPmdf0TsML+BXfF2mRNuEky4TWekLd/Z3XTdggq1lsy6ukYgHFxOznwiiwqTh
Gn3l2Lp0IMCK/OrrNRkKAiX0gjS3fLLf43TzO4hGhP3J3RQk2Pk6GKUW87gTR4PqsdOOiWPMbU63
I9NjCkRk4frK7Ll6H0vdG4mRkhOdcbqbM/rTIpdtbpnWQJQ4CkYsIf3Kf+C492J5xTZhWbNAfR5v
qFjDIlazigz3vXElzCV194h4mHYiNo6fWdGI2gsu63VotARJ6gdl40R9HeX5M26DbkLEoP3MpPEl
SUXFCz6f6kEwNLF8FqnJhx14ZVw72lRETw3MZBxbJux3wCNvgjjQrgfIZ4c280A3WZrSvOkr6pj6
qbw5vbI8+yGYQHxjt9SJXZ4jXXH5fhvxHvi0344dObisHfJYgSVDujszwku5DunjK1BUd2fTzEOv
QSsRGEPbxEVxSTupEzol/0mEhA2JLF9rcqXQzEE8e+qmQDrRoxeq49Ny0//LzmYvyxmisFZ73D15
lVEwhkiSC86K+ILbVuHj63xTdpR2Bb7UsVhM99RwcNfyEVqenS95ZzFdGqylGvkfT2c7tdqAZXtY
RfEkdshLNbqK4bcTftC7prn12PB4Ot6cWY5NkZqMfsvSgsiiBSNYgp5IETb0uK3WBxxTjYJ2voRC
WK0PpU4WA1kcHLadHbw7K2W9S+ZLu/1h0bAqWZ3zz3XA7e0STnpEbnzPWr5DYpLJrCQF3unOgbjF
n8JyJfCklAdVgHEtqcMM/ANyL22EEG7K4ivwXw7m7pkeL1TDnW36fYiIpy8wXoYBff6gnmeiuD9c
aLYMq4b7KW4DiMSnK2yH8lP7VLwRY+plFoJYeSfXA1AuO25u73rTsuzltesvyes9iXuDbzuyWm1o
f54w+qMP6uJzYkZuv6KUqOLCmyNOgow/fpAbfix0x/kSUSDfvsqYVJVMcH6ZXPkOFo1beWo8s3S3
Bgea28unwrWbGjdjk/GhxgbBAiPu/qYikWls9e5hwwYj1F/pBfhk5moyIgqQ1ZuQh0aH7pIoEDKf
GDj5lV1Nu9uYeDx+gPNYau9krBWWHcp1IP3JQ5ajGjhVR9jG/OyfJeRR7S3sbeBxvpnvRVIT5v4k
kT8vEGP8rSJJTVuzhFIOpnd10BFhy3+8l/yxW0npTidOPnxs9HrQCj/KiM3rTqrrbTUaHjIsg4GB
LomzlxQb3j++aGG84m20vh7XvTeRYxMLdHGogqNAzPptRa1Lslk8SMafF16KzMzkkUzpJE+htoFh
MycAmBh6clq+Pk1pLZ1ZNhvJsw8DZuD0GBIOG+/Vvf58vFqlCOru8oGU1ni7jopoUcyaS+8tnLIi
9hoLrg5q2Z5FeB8QMZbMW5CP6WUe9hVoIO/TFxbx5e4QJ26mCacU1RS+wABWD7aX1A/+nvJV65KF
fwPlp9z7PbJGHN3d3+8mNsWSfEoUuT/I5RcuMEg4KWG4wt1pm6qqZBWZRRIldgZVHHDev86I1h/l
p+24KuPQp6LiEYifEZZ5gD8dtJPwTowhSH9tIajO4aLSM8yaBC1Yer4U/lgiq4T1NCpsWUxz8hBY
fxSRp3DZ8Mi5xdy2BDCMlyq+ynutQ/CBvJE8C6sKACir02x2FLrlS9aSln7KKwK+pv/ObJ/cul2F
2V4U3plJGGHrTdEcxo4AU+MW9yu87sFRCMugCcCWud1n/z1nowRDl/Hq9zPCQfZwjyxjU6dXo0PB
sUWQI9KOem9iNnm0cwIaDQed+pMTd3vgxfxGuVL6uTdmC4xKyH2Kf8ntac0eKdcyaGU2BukdU/a1
hD4U9QoHqaDZ0ImHBF/p6i8Np23d9QyeKjQLpAcZFw+pT8rMCfnW5nHjKmrW+CVBQzrmdgMyu9cb
9hV5lCunLTIAvAqjpv1VQPBtaz41BZRiEvhcWJbD2RqVBm1kS1Ozl4aVt+HirqDMs3Va4Zjb3Yf0
Wub4rq8jW39MXASAmKjbtXqliKlxm74jOzBgmgsxyNaJVhzyk4XfLQWVnOdXcnZ1QXBAqVtl2Brl
B+8zEXr8A8F8gjb8uLub2uHU4IPH4LlYArUfBAfG2FOzW6J3QwQXGXX0FzOiquBZZWAdX0jkqI4X
7O9jpO0VZDPxoAAzNPkzWbtIiJS51nnNl4wP+1vhiJFBUYIvqX9LcB95CzNwcaXdcYK7Wf0qdanj
vVicl3s6zIwzYlgxhmRH/q4m/OnNwBDHDcKULKbqW+Nh0tAM+WnFvsgO3F8YtkcYpacUiSm+gFjj
LifN7oy32NJJRMsX+2Mb6n+iWDrCfCAJ8pdGfRJ4+oRXw6xtRFZICv3F2vuW0aRO0bCAm2Zntlra
3yHzHt6/5KBsDdEHMGcmec6TgYO3Q0e1hbLsuDjPL9MBK9zHvY7MCqmRs5dqypthYXRIfr0uQwZx
7NcZ8QqEo+C+QgAiDlY7GZSUTryWkTOC6Z2nkgc0/mbQfdZ6l53KpG+JVZ2NPkSgf2N+CQW1jbkP
yo0WkJb9zKevj59ZvuZXfEm9vZoyCavdQTTJV3jA2hZPfPyetrNrnsr8vd6dPDtCBtk8WDgu84XH
ZKuENIMfnC7t7nvBsCCynXNGySlKiVmWR+eJDmR2pmClxezkoGIwPnNDz5CAU3ZBOFii2txOGSka
ZGKa3KyzIt3LAbfcjt+IXJzhC010M9ECz3c3i2tDg87er73g365I/aPFTr3a+vPm061DKoT6ZUHX
8Pqm4eckydR1g/4j6sh6VPn9EPi9J+Hsrs7MVxfzqozJQTX6KWl1wgy1G9edOGpoe6cc0aOoouf7
L5mPLFaZLMiDExMM82jSVQPGcoA4e3bT22Y17c+mnHKE1JIfOBk9GpqbMVqSVoGEjoRosOzenBxh
WizbkW1XHOgmqH+SybDuS7iG9/cZ06cYMuG+Jiv7Ai3IsoOHRuoGu+FmJwV4S1+A/+gtv13w0sMR
ez7OUtBQ618Ak7C+lO7ekSPqeyx2/qGnBK8G7VPFFCWjgL760Z1fPrfCdyBn3eRXTKy1aR18mMTa
rN8KlJNtd51PWX12dhNppr5SA/+VdqAgCTQP8MCs5wjQxjXHIlKA+2v+pLzCUbYCCd/2j0o5KD+F
wBJ95ZksVEDyIsNKIYQTd3ik+0XBc51nSzgaw1s7HdWM5kCSvRtpf1+cfhE3CqiNGiorvY7Pe4Er
kQYHk0KfCqgP9wnvn2Q5EXtdOqUVyMdixXkT77VTX3IAnFct+DlVehNe+79elHmLJvW8FWsXbVDM
nZoHlHZ9jlNHCsZ0xw1Rn3TYrdvS/NjmMFeRvNVzEB6PNatVxBgOIM33jgJlMCCzAltrXy4eFLVX
9tWDnrMmEEjScYWOgxQ82hQRVozMxqPVFyUNLdrxfIR6s8ovBZpSuVaCY6qrF5cGm89qsG87ngz6
4qFrpGfnVflqUnuujZzBBDcA1xtAy2iyYNW8aHrhBvYORlsSCzcHIP/PRl3MYnuXOHDEIRUFbj0b
idjeeeaw2tEQh8Dv6GlsCaNbDNC/aSWWMb8ckA3TNLDN2xqB71VPc2WuX/AGsLuiuHqbVI0qYME1
uV/DFnp95CuLyhJMDAZyprHCed8v3OW7/CztuZ9mtO/i1KB0z8lNqYX+MICxsqIioNlqcdAfbL9t
0Obh406UEiXMO/+daCjiHTj+O9inXhijL7/lghvfBCWfCbk0mKJsVY8YbJKUsinFzajiVwauqNck
mK0lE/xHf2eswHrtpEC9dxV1nbii9OOoXfCmbEJzGj0FZlC7xxKd2fvbDNSeRTmzYTgXawH+Tf70
shSnzpfH9n+NGw4FQJecD2ysXBWFwkV7Td6sXQC61HXcqN5ufcARiAhXvb797CKcQOCNYbmnf86T
10PwdlhHkR79HpCe3CG69WsJpzj8y/ASajIcA0NXuenSGlcZoomr+1uabBhy9TEDi7Obh5XTrqBs
Ib9Fk3yv7hymcnhrorYo7g3bWtaZG9z3I0FSk7d7nWeoi2G90SjfyozIvfKQG/Ks17u/vcsT9pT8
srrulYprqyFV+nde7hd4LFXQcTzXEbMMvnzyLCaPYQH7jSrUGZjtveK0ldxHvhUyIf5ddFg99Idl
scN/daWwXksFLA8Tw7kvhcvRVuhxGvaNbAWalOS7VXt9rL2dSog6YAwD49ao0zPhldoNs2G/XO5D
qveCrxQ8Ov+esnGaRt5nAuhysgK3jExgQ9RxuNHd3x3XexPLYpYgmba0vHfwrogOerbOqw47QupX
bwMibjxXK7NnkHaPpLZtu6FlAngVy1FZntRt0d5ofVcGjxFjyLzFp1tHmA8xk85Wy5RLWFIry3sF
IhH+IylXqaITg4cQo4hIbl/i/njDeJM0SFJCg7YpNsSNCjIlxywXc52lpNMAE7wJQ12jbG6V50cs
Bjjdd/hSzOyupmTiIUkzSZ2V0RqdA7mYS1BpI2Agb76Sw0yQDVgfWQZBuGnXh4bKa3fsjhBKZVCg
4kWliuCA6K0dOVsiC+9kHYpFyZDdm2YYAWVOdB28fqQRGCQb33j1VKwrW/ZcIFCoY/nn1d4rtEnO
WU6zonVEIWx1mChsTlv4VjLABi/pUuoZbrv/QdkwQXZw1CUD1Go6RShdqbUQaleUf//6EL9NPvNY
4cnNFj0CrOaxtlPTKco+qplNnqqOvFfKXKgF8an6kFudbHYvtfJmFgI+X91IjC3fETPfItY3QG7B
9xojB0G+4AUu6R4OOuRgsXF4G37eblN+9wTTnnZ1UC4MJ2UWqpWC0KHKCZfMT+rMcozEuclL5piO
03jiYzrEAClcp3VS6eRiWgeefnjBIxCY4wq9g7tkPFJfDVsCHFhvgjPdupL3B3Y+H/1OJxoPqnA6
TL9aMORTR2pO+XKO0nkqOVkbMiKTaBKvfU05vV5dSzZA4tijcgduOXPBT+GCy+cTM41ZzfHEey7d
rfWGqM2wxRZRlh7tcogEapeNZ9AT9KDNtxr8VWojKMMkiVqqjIOIriA2+0Xyzyay8C/wSLQuLsKE
RJAEt0ia9hi9zRMXDFkDVPjRyhhjTUBo3HbTlIhmKjPZjagd7WDSaUa07DrnxoYXr2jq33wntxiX
4On8AJVWqd8l63NmFnT/HBasjwBJ25d/GsH9LBY9xMdhqeK3HFSXUVTuizuPnoxQuM3HXkB63E8K
q/uqFW3SweSSg4lFn7n2vbvBkq/1+cGnMy3Sr8duOk3PHUXrW4N6sgovQ//W0VvqM2RB5DPI/JGu
v9s3cT3U4k1KJY1Zlqad7I+OETwxV1ZEZhpgkoZPrTRqMMGimKhzFHVwCbp0du3tLREm9EBXv963
tcNaNilGDVjjoJcpnySpOOMSAvHNY18sKYWxf7/YqmgstVwBhzBS1rwOnFtqLpVmNju9i9H3COIK
HLBSmZg+l3tEuDT3bepjvFmDGSqrV2VQQmkDr1mk286JQoV8Y0V7SuLamvCNRdkb3Sgnmsgnb+fS
VUMX4pRIrna9j/SztBf/J05Z0MKLFe/9/WbzVfyb1y9rGpoTDV4rkaDCvtBgzgoWa0zogtZ2Mdls
eA6VraUjX/Td7Nv06IS60w/pki+plfHHkbVzCgEU900spMutDXBm0OH5U9dWPUO/lug/1Xk6g6at
Kl5wYZoIsysYWOYnY6KHdIdgpLLAYmrplcskYLswvxJIv16oMj9PyMJUKi2+LxwfAdXNyOBdavuX
hdXIPC8NBRNg6bMH8QFJuHq+JFurtWNUekHNm32OieBNWY4nwl2e42HJlwujNEVDow72oW6EKrEa
R7PRQTWFksK9GhoPYnEMPb50/PcfG81Xz1BQOKIZmSKqDKAsX9/HOrYU4tSAztnz94ied8AcBExw
FBjcrDb7E6swOyJlbIUqEgkDhw4Gz/YugVbbbG7he16k+Zr5IPcV28dq4IueTJHOY84pnM5DKyHU
6NtngFQZnqh8XnUjB0ee4/pfjbPb27eJ0cwbR+2NnC5GYbf29m6af5GeVidKIPBIPYiu7GSxqcVb
1J7FnD3ZVFJ3Gk4wWxeDyoZMXOYustUSPs9rrwibFBQtRM38pV3H4bqmRbS/ESLBWI/k6m6ytrrD
xtYp2mpgM+DoYCjdliWPYGsNi/aiy4VAVEm7B4GmCrKCqbh5x3ehH85H031OacUwYoi5Vjr9tr5l
zMWPyCiZZdCVVOngvgnZ6ldhQfW+15R5KyX8jQXKpzoqEvDj1arXvLCh+Q3GffW5bXuRxUMxuH7v
MEMAYuhoqqQJWt5BNtwsxsRDciKrVd5mE9uu2IoavCC0/oe7kUvuV8K8ojmEhpT9OzCiMhEdDN3f
UuPh8II6VBTf54MK86rXCA9RHYMo7Fu52E0aPXxIDPNCpCsU/cv18FPYyumiusPDcuJtYwUKx7vr
CloJrOBo9PxDaXu8R28GkO4zYhX9I6ZaidYMtKubWa54IHTUvdOB6fYRU7xa8KXk41/HPqa6lMgb
3sHiI5sd/cmn2b/vtnjTQ2s3DQHy5xpdWrV+nVS6HCUa/trIix6gIUuQpF1Ri41U57KOSq35729/
3ZtNvWzKVEAcopCHli8PUSFt4/2bRrglvTka58jHoMQxL6xTsWTlzGpZci9fJOzEr4Xzczw1vOx7
JyyMlLJNX5u+gLlSblcipprjCKvsrIbZV+P5mafRE/CKBfkdEzMFKiTOJlLIMFAvO8PJT7zodtWM
YCPJuiVCSQtRlqOD8pFe5q5bRCz4K8iP207+MSOZmaKFpWIa7qLN1dt2kBTGmdRXmZjY+2nN5wSm
7L/EAx4o6g3fyFGuapujYqQLYJNCbX4KuN/yICMz+DdmByHaAXhHznZfYj+Dlz4RWAZqe4/WxLP2
8qQOF+Z/27apGYQ1T6SvCldwe2iydBE9L0xQN+cDRgEJnUfI49KJXCyprP6gAbmHOaZZIjlCBC0C
bd5nxRcBXXv4yWifoCh5c8I7vmrC+CVE19WcbMfi+qRaZcUeD6LFPVfoUsmN9pTG5R8XFoU+7BJ9
m1XrIMfDpmP2wfPDpz4wqCGpKkYMm/L/njxBfVIUUBGr5l07EPM42D/MZX/b0jUnkGh7hsChHPOd
Slz5C+rc7tf7hkMV1d7it0R2hrgs+013AQc+K8BMgO5vP4dwN/IDykYm0ZP0ygdqhb3IPV441o43
H615JllQm4ga8qNTQTwbPkJexMurBIR6Y1xdSbnblzvT8T57/cNr3gqlMu7eLKofo5FtEgT55Drp
yb4dDtgCwtELf5DENqNoup/3XtB8rUYxIUSexuYn4VXr48Y6gC68n98Dnn41NIDpq3cIPZzOJQuC
TZSaeQV4zN3OnvDb1GGqGDWqVcR2UaLEqnEvmH+9bGA6svuky+ModCxE7YjRsb57ouH3e2MNTw/h
3f7xg4IkEYPY3VCli+IEN0GDB8bfKjEy6G9glS3jt0yN8R4v4veSZk2CtHhgZNQtm7I3f0DzuneQ
0NIEycjJN90fNvbIJ/YGus1ugJS403jvmNyZY+wCRh1Qmibttjx5kQK/w71d+rtQCPOmXsiprBEE
WZ9zCnk/FlEY+oNbVo7uiL91koxM7SFIgAhtqcBAlN5DN1VQQskXZXdiRb9Dp+kF9oxiBzN1EYwq
rc2Vhfuc5d36we+lVL5XrFlwCX26pbeBefe9NjUNroFq2YoDJ1M7PiF3OCw1+NVaRP/c0NFEpZwI
gyRFXE0StVNEZatq3Aju+xJSq9bChBwXq3i35q77LFAPCzIFVxDcgXy/xTzJT3DIxpqrImuOWbAk
ueYO08SCjN+GxqaQn1bN1+BtYExcnN+5aVN5JJj7lg/bvNU6QovjjpSKAgPkWSNuqJQVvZp8ADeb
mTaYdmFf/yAD6qD1eGZK6EOmqtfpJZvqnwFxQCGJ4e39ewqu+YoexHSaKjQiU0Xh2RXAHLesvDh3
aEusbAIKdMuCscx2xEAcvmrsBLvi22m1ng/ff4omHbPrJ2zyEQhdMcC1vQEbzDGwou7GK6TOBfUe
C/tv76dX3h3mzuhgl9tpfTTEIlf5PvgTGtE+LQKnTF+2D6fWOEJrFvExKlsE1FBobCTvBZBxOzcc
S5/ep+dgIDXreI64A6gEn2DC5LqmcSvkBbHO7waEJpuCEy+6L3A9neIKAGwM4F+YPnpmOKQXK0Z0
BT/mMzTpef/ixTLs/CqKrwuo0HJLhu9+PpePYwWTZ8y/tIDhavS9f0xEG7k7jMHVcSTVD984fFib
Bjqx2VEJYN2fOc33837yoz+tjkuwM9J7wEk78NOUdLu+kYLSjZgqxtIPNfD4QCKhp6ksTc8RtmEX
WE0cdLkFcY2u5UPpeTiTc8YlqlVDG9dbAwtRp84tG8DtwEjQbporB5QJL2jEWoCTvCZt4fAQEjYp
SYalBAAmbrZpsoBjTRFM7ilm7tcScMiArd4UHkWRVnnhZgBl/a7JFTMNoIzfFj+OhY00PQAGi8Ju
sZHwXBiG4nbTU1u5mrN6wW7zAUHFCGs+EpnFyHoNdcH/QSoAmlFtIlt4ZmoI5dXE/IvsnTxlCwKq
7aP36T3vg4Xa+R8V2MOc/vcNBb5a7b7xE727NEWPKxYag59htiBCx/dM4/6AO0ohK15qMNOSG72e
+NZvnokjGlkDDYr1H/Hn9OIIv0kCVyZ0A+tB5CzKUAbWa+rnxyD7gWPM5Ohcld6kKzMH9zs8GWQ0
lvp8ZHCAlVym/nmXFZYWLXVcBJ2Eyn695yFBDnQNf6oWWmDQ3mfmUyCqYCcKQ5jxdKhzOehJINh2
QkPxf1DWoZ0JzChc59gCswdJ39XXB7rSF/ebb1NZ4q2dLt2iwYm16BjnBJsl2C4RerqTY8dQu2gb
J8acfCzuBEPSZyyuQOsi7G4Cofg1congThTQgtdoRp73FoM5m6cjcATUF0fR31JondwXNw0kKa5O
XhzlyDWLLIRNSOr77HpGJB4WDIlPDKLXNP09tR9iG4F3/NVLFtNVr8u63tIq2QE5JoTUHbKg9VjK
vXVA80/0hWsGwNt9BiNMbu/ytyQSDH8bC+3CzRPrV6LaCZ1Nj3p8XLXeWOtQZzV3Pmjsid+nzPm2
pjrne43gVpUq2OknJHROffv/XaKyn5bym81IqD+8saLMCa4/aDjQ5m7rDefZ7xsXYyD7YCQGlfZj
sbXeJhKWtI1OhTASYsHYvuwuLU7vjsgHorgVEMQMueQyQ6aiLIs310aV8f8UF1XoZdi//kC+Y9t4
VWQZhtFoD/nDVW8OWYfSy9MJdzCw0MKb3RM1mFsy+awzuU03uyWClSdVDNGdwllKYxJgcPNB753a
2HKTYVOZ9+Hz3T/sd5eugs6maZZLpL3g8wpsrgPHzD24MPl6ZomSntOnMrR5nnAPOkh7fAPYtnzn
nBX9GUnVVMT0rc9vGPEO0GhTMbbiTF2JUKpVW2Er8LSp5qH15B01FCCvdFex/qT0dTc3LrH/z1/s
5Uiyt6zySiFZCNntjWY0OC8/ubAHEgsovZvN1/R9v8AM4Ss9Ru1hFoHUdEODDwgoW84n6vyoZazh
MYGWeP66cXZIvHNs4ZJCmRDje6tO0tk1mCiODmrCkgNYnZItMYDANEkz7cRnthYburL1YioljEc3
k9LY3U+Qe49UqeP8eIk2KqMsyx2ZHLrMmiohgtOdB4UGaaynSjLR3biMDIR688RUQI2zu+lKVYuE
vbzIU3qwmWkPNZyhzTZ2txa14+8B5lI+jLdDeIcni0Veg8KDJH3UCQPnw2lCyTj+OB8T1+xVXZkL
3Gdk+tPu95MjJgwz4CDuxkeLQKKbJgrRsPweZGaDZk+98+N9tOjHjB5/0/uqo/HYjER7w3X8vGmy
29yiAaDITx/k+Fxs8qfCTqtmhgvYobVFDWiaTtk0BFIhFebcqZ8bEPkFnC+zW6Nj3F8/1eNWcpZm
NSiraKwwhjsU5eOBj6d11WNKF2EUaHRn7OSQyzHrQ6Q8UJYpfNWB9IVoMvTsHc2RabfvezFmgo5L
fAezGHBpaMdE/HN7u3O7GgbdgM4A1VjZvztJneqrmtEs86TLF1Uycnfv5aDCxGi+8Xj4P1B6OFxM
w+fE7HwfC5ISl2IH7mMSjq/58mRp+vOPIj6qsfBkFn9gPWWMgmlnGmdWkorOISkRJQgcwTQpTsn7
c2uH/1FtAP9r1yyS/gT3PPwyFf0/BPcphrs7ROMs5F6d6qJzeE/POVbcWGW2lzzKxwaY4lyiwDni
qXKOiPHy8UTnEn4y9v8xWKZw2HReLt7zhlFB9aWa04TnNzzvxiM1T7eX2pu5OveM1SVPjdHK9c8U
f1aXGD8/pX0wz8zsTw1KSQJQ4SSv6jjzdaryc4hItMtAeXUMwNlBdRdEeoMiIrf3+fH8thvpJhXI
roLogd3PlHPrkWzmgGzJ+h38iwPwYJd4Ns6SCBjPpYw85yUd/y1oWAPRr2bDjvTppPBwnWCATg6O
eHZl9p3k+yb8yropdSf9gqFD3XWPPKhFEAjCwWCq0h2zFX4fd3Qf+Zl9EbMlz6lqQ8arWldwWSV0
crNRb7eIak8XN1ImYv+mWWnRMgTnqCJPu2JSCT6ZXNt79SzAUg7oDyhBdoc9E5as85o14bX1Yv4u
0gt4oZGvFyrYJZAkNMATFZVY9wPQaJtVd+GYEn2fEQkuwzi1Qv+QiJk4i5hTLlAwhMVyrZRawTB2
JX9PszL9+SB+pku0f6yxEU+DxaT5wun5I7dVkwKv8XubtTh2ed3phSYk7ixsiHrFc2Xfi9MvZ+HH
XymsgVyU2mzEylGC/7tIZ+cwla7AVEI915I9n05QznnU7ZlXPd8XZwqzlc1IDtdOZ6oZfOLTy3G+
Tc2f1dZh4ZZw7HVhvK4qfTCdl7SOOUrmxegPZQIMGIg71BABJrMmn3q9/0zk4GgXEbfJG2T0Xlli
o+n4akKTUJE2lwML5BCmM2Iw4gjOGiY3Mcaq0Jl+4WMo6CgtWwLuC9KmP/BIdZhnO4hjjQvnl31W
JWG1n6BM+HbhWOmwGO5z/9zamfR83dyYM67qh1MnU8cPcPr8TA9je6QKBKR9QmWq/vuTEF3V1Q2L
gQltgxiqMDdcBAvwxHECQFeua/r696Kb+eeNWgiuKfbZ5HBt1l0rNABd1XH7RyKlc8azPhxKBI17
718ZaEA5Es3W3ZxWcblyoyXEIVzDsIs1Til5mX5acoc1kQM7JkrzsU9pAiAczkxbbHKHqhWKzVko
fUkmE06e8u15Xcc6yKYqYzwywjuMSTaXS8i+nZy5VWsFU6y5u3Vd6daGmOzC6f/bBfbKzw5rTIMP
q980fJr1FKQAt2EWEfWTuDltmEPU4NQCp/JJmD20daeUAOfwwyimDRflpA5Q60cl7ixIptNBKsyg
QHs5pSw7UQPj648n+bQ19xIhubAes/A63TsOolHnrPgMG5QX+9BvDFGccLmd7Wnmcv54vIqv4RtV
3pdRfvSZa7qf49/YML1/ejuC9dQxnNOyF0k4wKGFctvc3QQik2ygeNHKHveo2mFWrF2mbA/hq8f2
vP3m6/08EwvaAtgFqIpMxgCfSLE6fwxYTp9tJHnG8H0PcLYUlx/E+TKmi99614tnBjjXjndd+jho
8S4UxntL1wqtxM2RBXJw4Sr2wLjHrUb0KEcwp+LK+25cXVdKCnre0BWC618cGrSLHdE9V+xXSOrE
xFwKJ91xBYfq0e77TugyHOcdcbeNStZHQPGpW+sueXpUHbGcxUNQYiUY6xJfh4vI4UTuEupTHOJB
yvsU+Bx2jcGXcBWoXCWIENWxXaLbSWEYY3r6acxz+Rh5OD5Te7b9V4nyUMzzYL4CEFM+lXjrn1tj
8zz7fXFwAE0bWUpVu/zqTU9jMkCKaxUYqa5v36OzNcNG+ay8fezGsICDEkkzwAD+pJpiYyCyBZVT
kXc9rLNSLhxZ5YhA2n1s1kPfiLgnBPh+tZ491foX4H5zjyYCzhZtgLVsoQvAQM0kLZjO2V19NcuJ
5GafTanLsLEJ2xyd8fKYGrfv0X13v3ccxc/wwB9Q6s/vbxNZ1USiil17lB6DoXtNeJ7CqKASzfCd
J0HDuRCJIZjNGSVLe4deUTKz6bxGHEhNzeaLAEETcadAE/AzZDEaBj6P4CwU03385qASLKr0fhY2
mvr84jEjXCGuFVMlSv/aroR6r0r8Ys8Up/9VwDfPIupiX9fkPEko8wO7ya0Bn21OgHypb2/q6zPu
4RmjObqdOTqEjC9oEj2ZUosgRQknxq82XPutF7JN5TIbReS9n0B0cUkciBlvwfyFSYNgNn1dxes/
XqiQ5jGa+SRhbxZzaE17DLLO1Oz9xkRoLq3B/RjVZ+3fRf7fuu//+LPDlESPbpWL3WvyM3STdKsE
gYw7h1XGKffWOeAHwvyOPLS6lQ1Hrosr53Ph328dVP4eGO+j+QdPjVjZK8A7I5Gb+3sfanUALaE0
VFFQCZ4PS7nmOioUyCxStMJNC+6OoLSiJa5b12Dt/e8kUdkueMmu/7om5665io612YWLNe/dP1RW
4x/aSkjV3bA4nci0EAgoUVxlp95eW7BaAnhxk0HLLn3hNViyKcjTQezQzHaXXhSIWcSGQuZ0NLjv
CKRouDpfaz49MHTNaSvaF0OueAym2SF4N6GvnerVrGq9VF65WZUgHmGJOA9kWGvSOxp7qRAna6Ms
XOHVr8xkdqEdnxynKNhCNtNuv7TFmRl6fEKyW9XXH5uZt2Xb317QUpsmSFEx6CwKOPxQcmBvha8W
Q41ozdYGtZxAdo9lSOtjF1zYUNFwwGdrUEaBLdhyKofa1jqSyWQo3RTjxtNTJdO4LGpZ5bE5W+gP
sEpGxEcvPuSv/KyoYMLoUoaUmv4+VHYp30xsAjNzV+VTtpqgaKjnY99Lln41QSwBr68lTG879gNf
RLJRyj/0E4zgzA/q/zbcGqOfkKl1lAUKG7UuRvgfWpviiawOGUvPw3AH6lSTzqfJM9zxqUCbyiyL
1Sh+A1GXtAgRLXqaTNfxAsErYkCoJayL8wiBsPB5M+YiWdRls7dS8gEUwVhpKXILg5koTt/1uEfM
PM3y1wI2yDPa0svzDLnDtd2AEWVVTVLq8e1sIfGpQHHXFhj0bXfkH5z6pjpls4ePpA4JG+UKslJd
dvtYoC75hF4Bi8egrJ0hY0WrS3rZWFVmKE1p69/Wwn3ZTN1DPEYyPCQAT+Ek8inR2YxjF4llBr3l
k241hRIZpocIxhdrOzcdIFDdu0syIKDM4n/6VothOmGLpv4w7FRB8aX9ECDVjNYI7nXIqUB2j66T
zwqvM24csp6ONZgw0eGAXAZic325af3qMkEU3+kOXYRKIKkA4lZYHAiAjPZfSdSn8tysgPoc4l7N
7umuaopL8q92e7KbhKpyU1yWBjgSf+SyJwuzWLSbBqAN5F51SfOxVX3U0AoQQiv4SyFjONenWIoo
8mAYGoXMM54qeg2yt4/GD7glyxnfuEziJxetoRYco1Tan/4B1GCzfsWy/7kS4Lq2xeC7UXEcvUke
U+KwYfk5JBY90T45uZHWpovC67JfIQsmLYTwB573GC5sDAcqkqB83R+5dJAvoSmy4P8dFuDXnIYd
fv2rQJO1a+VLKVWEj7xI6ju2h1scQYWhX5bi912Ly3yjqIHrJCBuirXixRSr6YR3am6JxJgTfogj
yukjggzOd3E/nHB3heU6Lc3cvlT6F4NiNqtnEHsTVNVyvCk+vbnkbdc6/avU2pZ0yw21GLFatbQK
YTlPahpMAWGIB92MJKG4rtGp/sYVg9x1bk/QvYHvDF3NlnZEtX3Idr5v1XeZOguDfw+7NaCoZefO
G2XxK4kic+Q92YeH5akhMH7USRVo5XRRViYOhclQtot1/kAMUjF1UfZutvJp/DgSAfyG/qLROhkQ
OoEDVdI5gvtyaykC/fnq5L3Yg4frDo+sWoPYiboOy4jQ4dwSmULlFANWqHFlRYdVlfV45FnzPPw/
VOgChsa3vxeOG0GUNNSCRggAfzpVUTXEPrgRkm9mpE/VL4g8gyjjXByNmM46gSaAmraBQEp/tC9E
Uk4ukhMnCi4DuXaJML+yBS2TELJ4gwSDHTLUitGonHnP5eEk87FVcjoliVG/mkjAWz2w7acer+Zf
mVW+GxYXu4HxebhQhAOX/Bsc2ahQxNxEQTMZKgIfrDW3dVkEoDpI+1tDbSN7kkvtOjJrPNlZtmbY
nPiwtDXNjHP7WmKNqFCC+84sH+Ko431Sx9z0BCTBvFFcjgTxion2o2D0N3h0YerRq01T9l3kjBIx
MTpJBpuE8j2AlO8z0oZZLD/38puQ1UAdOoXMmU03oP22SvG6gKVQTTt8fvB0bthaApho98vonyTN
WXQGQu8ngKznLxcT/elBgKRAGk/FhfXOQ36J8PAJDlw22thQnFjl/NYQFlg1whFeP0VMPda3K1kD
RFMO3zclNTl7cEMesqppePS5Job6uaWCLYtWGgtuXMfc6nCccHZblXtcKM8aeThvU0NuLupDi1Di
2T0BsgLVemn/PXc/P9IZ4qWD687hYB96njcYR0RAb8PXVM0LkU7XN93VAq8mAtBtffclR60D9VIh
EaFBS1QHKsFqUFo0f3sn0e6dX5x2VlXRPy7T5xx6gOVeZXfrV0uLsRJnGggTkLYCUvhjxDhBLnoi
cOIlFqKEFWprJS/B7QJpi+KSzmlRgV6bxNWuR6HRlnJLJOsR2y50Tmdd7XcZSC940UImdxvVbhJf
QMN5vholLtngsyjl41X7N2Jkb9iwuN2lZ/ODui47y2qr4/5cWP6QHIlNRInpkxmOI8vhQ3+6Rx2C
2Z1zI7DXriGyh0jwmHka9tLSCL1hmtjdDZd+iPRldTVOclkeBLHPM85ZfH26xWdaJ7KbgXNcqxQt
cM00vVYYnoFQ5UzUBCDIg4YNSxbTcdwOHQGXavh72louOCMcQuy5gX6qCrXJ0fxVDnw94Qhg2yEx
A0RuJ50Q4m6LY1iPojRIHWSXQaJDVinyMcylXLFhNIu1nsLsF8QzwZkE+IO6jtTXeDWxe01wcrxa
ddVPut4lUg83tf/+zOSs65+JJXFGYpGT2Qs0//fcnrcBDMKFHaJr/KPYZ0RtzvRh+Gzm8ne6O29d
l+huhIscEBIjyFKKJ4Im/5qqFQkJzyH0D5q3qJfzzrt3BLK+5DyHJhiFa9jQmV8/IDs98WuT4QCg
Ik5FGE9sIIlY2n9ruCzqS2J10uMptCknbyihCdoRqnn/jDOdMETdxUWtBMTnHlP9sXTJMm0iRGEd
qbX9Nq4R6XaXQhSGkC9num1/2NlFkuUfiv6dntMwtimzjB6E8kCw58gU66VJoPHR/Se5tEVL0qIe
X4J9Eu0biVs2tTxuZ12re30e6wx2wqYz4FJ18wV+IxW6LuHD6+G5pLFKvC7BYFSkrkv29sXjfnyK
FrUjecilE7dc3jo2Le3Rbq6Z39renDCGk817Xk+A43bbWTJouVjNJQNv/4cPcvYF07aMQeVawIlA
UqFL2yR8zxM9rNZf3qmnOOTlTWhGOddanCfgo8PrMHY28iFo6DA3PhPpNVVw/2diYF5gSB1IXNMF
wwOfmCGvKXYFbSxOLSey4kBqAt+d48Wl8l0LHdRf/LFcxzcx43dXj5bhbkUvvkqN0QGRUClKM+79
p9IXzsxWdA+6pY6DsnBlywUb4S354ZCSAQEWmoNI5zHKKHo6QvZ7sfVYY82ecbE+FDXGBF88AcoH
Aj7pOtXBoTlmFXRBtbfAyztcqv1BTkcl+wa41UFlRwFs6jztHEmn2d/3pD1EQvHZqvmGDziQcjrn
95F8XOSI0/yDc+eZsa/fePSTxMvZgmGTRq99u+3WDqQwxaj6zhEGog2EnZ6GZRuQUTP41CQyOnWg
wZYYTS8IPEH7/Alvl6GKdOvHC0i1mUdh7TKcuuxCr5Y8locJNMWfTDKWw0Mu4j8qA30HC1RNS30+
IQB8lDLcEk1/LSY6tbsq8axY88zmxp75LVQgTi8ZA3gACLtJXf/iuslzPo1EqYAwR1TJXF33AH//
NfT8cvtdmtR+4iCjQe02fRwrys/mep7SGho12UL4XwhmguKemMqhlLRWdMwBrxpGGmcaNowpt2JC
Jf9RM5fhfagK5dTNFBS7goimzxzapExg8akhOeSAJLzlhdGrOlGfxs6vqHrq5AR4fJxWQhp8SZyo
jaGdRuSWazFltl91Y2o+eEySL5S0w+0IevukM/fQcjaQopAR+HuN+jzuzC1kXe6k22U+Z8Pt/cEl
nundKoxDM6PtrGsDvQ0TngGxYOoli0mzB4yG0ML7eAvj5mztfuXqmNL4Idk3kdtrkIMJ2XPrd1Sz
0Vg1JeZ2Hf50wNFhNgIUKESYjCc1wxNq2kuQ1ksts0CMWYHc7sMHgUoAGVf8fHmQu1JUMop31Xtu
ssjyaQthh+KGtkBhTBeOtTUAxvwLrBJ4kp2BydDYh+mJ0+S9hoMQiH78gcABJC0zxpdYAuvCRazK
k04bJnMrv3/XF9EHKbGujPQZ63QiSKdAtl0BKr8223liCPyyekreoTiqv3xKak2m79bxvluPIF8r
jv/Vq4HESgQsxmGXe6p5aFmP2qptH1iDlSNweuJoZ3Co1iHDbTyUufp0313bPmCvlaeaIeQ7qKaM
+M8ylfkKFoNwUIiYhjCen7vOjqxTowcXS4Kb4CohLRE5it13Nw9cugAvJT8yxe406O0blWXFoEmK
pGymqX7P2V3baGWJ+TL6tiZvteIoAyE9lTqV6IDX70c/Jngh/hsOeJs8CPv1or9MuOjDDrdVUuim
NI8L4l8Fteamq0VR/Iyrilx7saZiBC93Xuk+yR+qiP2RA/opBfLUze8ADfHEmSFBdYBR9uKYW2nE
30R8pPvxAe+6Qfv3CI7IZuIsjTEbzPQiLCh4loTzvHABFWzw11NmZK8/IBk0DyDWyj3U6t8tgR1U
RO1fIvVmJJGf8uyq07OK4y4P2j9h3fg2jGvjkZ/NebaevYLywEVPtKlTgdEkzBj77tfNBY7qgf6O
dVxIEtHs8tGbdZOWaxP7oZM4kIczTQOxEufVIIzSCiMXQcmDE68ZcBDGZN1SrVV2mq368eLNe0a5
5TNcmp+Dmglj1859bfkr8I42EBbkZjspHpYVk7PCcpmEamIwUBxz4KBvyaUPzmVkQXKcckrdXT7a
bAkiJHv1lhQTrOLC+wGGB4Ip3bxXwsKqRmwUMIVWQmMBTSiTYy3hjG08faKI0Z+RpA9Gj3Yzae7n
KpY8ApGheVLgKY6p4x/85QI+l5AIYMIiTejm7Vw2h2nk7VGpe+25af4JOYn/Om9ETSbwr3m27Yfl
NWtD6kzxdhP3jwcyl3VCY/REmOcGx8zlJX4Oj2HP4dN2ANv44qxZ7+jgBi6+a6mJ7lQUDGX68R0W
mnC/4CYQn7jwbaSo+mZa4b5MQoGmEbyEt4AmzlBQwGbr0Y8PqZ+qvpyYeg0f6lNgqndgAPvtYnrl
x3QB6hvhRl60/L4At03PJWjxas4i9sV8YNETGyxnmaw7ipCO4V1FCMorCBX+lkNi1cEM6n74MVrF
cGboHCVvfo8e/yNhQvYhQMyMMG9BjGKbkQ4SbaSKodHxP3YaUbyyIG3qG91eU2DyWrBrH6w3nlWV
ws8keW9vGWKyy6qEtDzRIcqD+KdceCYQCUi66PxBO6mpSnrH8l2uxNPSOINOkF95GP9h6ao9jKKV
f/HLanRbJnwKHwyxV/ZmQnYjlEoH0Zrs/qCqa5+m7KMk19Qzds3cVifozFUI0E7O6YhUzHCr3oY5
JpsR+QeKHhbUV3+Li6J5eSqadrn3/FMDADvbcodJ6vBO5Pc5X+WYW4EI8ziSpB9Ul5CfPZjDLzn5
j5pzKH+5z4YMz8H4tenUru/NDkDv4LA/OACsLZave/7a9ys/YeAfj2EyWADcoaxv9Nq/rxWGuvOJ
VunViBqloTm91dhECfHwbe6HV/sgmM4n7HOk6sXe/q9IYdRXIGh+d1DENnNmVGO4Z1+hIWpTQfeu
4SgZr9K+wtZDjvkz6lmQ1+kDItZk7a8UUYAbRYMN0H/QHndOCyaxZ+vHfjDVJ26YiMP11oHmR94i
h/KKSTyXGCwjZvpA6vzCGa0CPeuraazsguAnxAssyJFiMfmR2fousHKjqVtHN8Z+cHMM5HiCB0ul
z1OLgChQ5pwgn2SaipSxiJbvEUqfvDeqcojRR5dzkCeHVvQp9BPGhS4N/s7b84egQFTSsE3+8yor
JbmC4n9FKUxKYN/07w/LteOQl8NA7Kq4YwRL1OtRgjsugk+Sko3Jb6bK5GzD+gXdF59hxKnLMzqq
TWpwJWYEDAawpffU4CqooukvhVfgXO1v1YXYal3k6FfRGlJyrqDoT+aueH73ng4ta1M2PWnJ+mGW
oMAfFS3SAgsRjROAL4VcNRNdevaf+k5/iLbsW+wbl7RV5yfrJG1BA5Bdm2oJXBu8nD2sghIAZbo7
7CEY0uf4U8tpcmI9kv4kX1xGRFvIj1BtiV9VPBhHP6w3fsKZvri53H+Ukt7B7C+RbO4maMCwPuhl
nI/qfS6nN9mrW1ID4Geg5UPMrCkFFfT9IuKRMbGCMDXCQqQ5pMLvkjNeWB7irDtHVwCCtkVlBJ7v
0O4pyhSHL5NuI0jeZgfIEOTE3xt2Nr/2Z08ieZrpyoKE1BnQiOn4H5zy8pSSvEOw+Cg6JeA0tMi7
FAUgM4LcFVjnJzksaHuuylyTOqL63WEpilOeW0apQC8+NUbrXEIOiRyR81+IzcZsZ7ewbFS3pzd8
a5+uLsN8eDKJW8O7vqkBNLIAtULJ4FWUYO8rgRP55C54TQ7xTpMRrtnKcfTkgA8eyy0BK4ILJdBL
VjgOt5EKLZnITdst+jpYCu3A4suFKAkgd0iunZpVN4dQqVw1myYSVXt+VBB/if2ayoGRe/OB59IH
2IOfNx2QiNXsT9ssIVVq/QzLOL6KQ/1rMrw6YVr8cV8GkwdXvluLvyA/y5fBfXfnXSXaNMoathcp
P7ZcUQtufPxJ1vbod3gbFtjZIueYIOcLSMtVA5byZaEOTnnyfD9y8fxki0AMDv1pTgy0+NYGpuc3
Nq4J8oNe3qxZAE1CG2UkRO8Bcs2Ugvtdj9oMmkQ/IASFz0Yao5jpWUx3pgQAUpzTWkhVolSQBN+o
+5g+f6qoQBfV5B8ttx6sznI75ihutPm4PZxlAe8PP8gwFUexxKeMrVN7sezi8ioD1WqMQtn7vSVn
hdPksQguKtFRtqlLDJ0ue3W5YanCTpz0j3zGX7+XTXBKuYJ6TNel4F16mEW1rTsXSBhdN3Un1usz
mLUTr7wrDyG9Xz1mkX4u36+pon51NHGstqJaLC4hUK6sOHru1Ph6fYn7lI4uJkMnOGrFrstPFipW
Z1hAdM+YkuEv9EMVAd0XwgYmFWX9ZY1BgJ+eShW838Pi0O82RAAh6BCDn8rE8T5t3HqfDGuhojDn
9Fkh85BSy/w5oX3o+2Ysy0J76G3P1/kcvI8OsTzcjThaqiaFfPT/lkV59JoY/fae+NI4ouPgOAiA
ACVKcLt+HAAjCbapOf+DICiIzH954s8mGIGn7pEAtbeXd0X7NlfR4BYZQ8+o1BKaWZCTfkP9SfND
mGG+wmBtRTJEPm/l3mUwMteCow3gLsP0YsFGdAv+FSQsMY9U9FbNMDB9Qkjk3sF8ordeor/WGgIp
htIspn5mapmbFTudsR6rPH+P+STUP2jGaB83ljObaDMwqmHZUx5cd+KUzyEaUyrBNvpU31jCdtY3
uMd+di2BB3C6/zGUwd4C/4i1SF5k7VjBMn++nR2bGdx3duzpkj5+5eE5eKO+1Bq3Qgp6qWdMHv8b
3IKus6dPxVEKeC5xuYNZf6pB2zqTE6gXGBlvPO6/O6JdF9o4MaHgoQm5dnzyyCKXdnhE6WypH7RK
K53x5RjiEbm2kF1Ywq4Zsffa88PkIquW5DoUIlWsH07q6uc+NnkameHZhxXEBwxvL5WDilwWntRf
s7JEYGqh1/SDApp7AgdZaQ6ipDvasnoC7OPjeB9rq+3Uz9fmwooNz3//jRp1f9pPUSicyEHMWiPA
7aLPfS4II8yU17lBoNlm0+VEAFTu6iLbXS2tW2x9tMbQWBtGWoQB8wC4cJsK1wDDDroNJOXHfkvB
Hs1N/cSvU27D/WCi4uZuKQdHE5Z9wEqocSB8fIZjRlaiYZNsdOkzavIx3XQs+xpV0xic5fNQDBf9
K/uArTmZUT8Bwy1duTF2cOLYDM/ulETFUqTYqANz7VmVfn95S5E+yBz+xhF5anaiSLv6H+Mc+t/Z
ttBepz+aZ/7mr/t9z9jTfAnhtF97oz+rsh0hMZJqNig6yzLgel8f/4Uk9Xd16jWxTS1YGCtezfMi
DLPz4eue8kzocmmIKrr/NwzEjkvvwCHkURERKJYwPzPpOuQ7+skd6hloki+NytbBDJ878qwumC6Y
12czgTaCJ/z+P6V0C0+3P7HZnxTjxAjC0K6CaTrFKoRpjAtT/MiJugp5oSD+J9txCaqeqMWDS6eq
qW6zkeirMTQ7bZISVN5QkxBtbo/wqd0sw+vcR/KPwTCJdsQ13bgM0dzXfitzkR5udlBvH9ftHbll
lRTc/By0hTxCKM+WCh5WYvP8pi95OAgdQ2Pxl07RUmTeJ+mJ6vCpTL+QitcsE1NhCmOPq6ZrdQBz
f8Shfyj07FPLuz4oTDHco4DnpvohPjWf865VO/YZTnOqfgImHjsun4rRjNuvyZ2fecxpOQWavgAu
VUNcQt4NlX2I95/Svf/0i8CwHDUBzEEM48sHK4vMSQVvQG3OYS1cQu4abmGz1WRbpUaH0hy86cjM
bJ4yQw7OauiuRJ9MsfQOViQy4CJsifnfDAtMaKY7OcflOR97H4ZGVhXBJ0sRbZO7ZytfbQxWDo/2
AmdC6+ujhjQIUCA5GtyLAvZ48yQFxzIXkzE7BZWFFaqSslaFUODwk3WHuCm3/bHnf/6PwnJWkeKk
Pn6pktNIRTZp9/KeY0RsxvD/AxKjg1+5SZ9sTjfpRw2y9TnyxW06ppjcaB56wkq/BNhBHuXyezp7
APHUdW1N4jTp6rYWtpZy1pnOik3n8MEaN2BVhVYM/zM6iSyK8hDB4cvOLzMPW39AMpto4ZYnvx/A
5CbOqlsye51i3fzxfiAR61vRnmkY892yKx/3maJebrGb72CsdnGR3epM8iOoWTivIjaNEyuUS83S
U0qJLgbKRfW/pAIkLfycMxciMQ981MRjbgbFvrLMPNEPXVNIcmUTz48Vjgs8nKzYmQIS/wTvIed1
bVGF3M1yOMyzPL6a4lN0zy/srmqmHykqMkXDMH5G6dEd/W5KW65iEbBPSYH9ScNL6FIpUkjgRiGH
6Ni8MZL9rUJXS0PuHuXUDgijVo3hKX6Owkf86NtNrGUNDybYyJDFUYOsAQ3bU18V833wJrPP4PQa
PKFVEQjT1azGpDo7KevPbnDADJRmUTu58QlVd7HSVX+8CwSY4WIGZTS9gctRGeU1A+O9b/k/duk9
R95UHN2hFUxh0nkahXn1RDX7Y25jDEDGuGaPePxotVVgCE5gn4wJjL5afAoxMZz2S5JYFBQmPfzc
ZWwLrL/2mOVop0YppBO8KQIHSkFcp+DNF4HJYx8CCNUjWhGtJb3m2ELLU7V+nG8PlqzCWscyskIn
2PJrm0Sx5pDyM4GpJYCCa+jiKc0rJzE8xDaLcaOSwAfRCBYmniCpwHh7n8IbJ8R7WloT+F5lBkwN
lSj4S226vUNiTBsnqfiuqoXiqkK7HrFtZxqHe8R0O3TdBzitNWHD3Q5Iie6CPspS15FxZ817VCUp
jmv65UIdvQWpOHd2LsLello5RiK62VS3e2svdNA6lfPegOpmH6upcj2y11FDaaZ0uKUJKct2rDHu
OsMAw/KXczY+wAJO934Iczm40vngcfWWjpg8SFN2PHRCIj698kq/7J3hOLj+2A0XFAvcFnMRTTXZ
vPscZiWG0qLgW/npmZNl6rEfUM2o6eElQ8uFhn/VXvykJX2rjR0fBZAnpaXoeCN8qdb8eFYvnjre
WPBonVPOEi0JwuLktGPdJfBWZJMAVv1OYu7yYMM6XsdHJ8T33YcwzFjXBQTs0NXY1G/NkgAVM2nh
MGLxN3zklKNVImrBaWVMz+lL3LnEBzJIZBsU3bJ0pIwF29kuxygbWwZK4J3PJeUXKMK0AodFYxiA
U6/cNIeoHA+6iP3Glurvv/n1uVMQwoVkiH+++zPc0zlQCes3o6/XmqYMTPA13bQKu/9si7f747ku
rn7KLb+SxSadtrH42FpSjqUwX0YX3b+eBIJppuCExzZfSq9vdCej/x6Nu74Zt9XlVxjuOIKhNDqN
jH369yJ2MA6FUWidLbSuBHjMzOeue8FfrQJyY6Kp8E3rCYL6erbUElxLYqK61KbDqFBHhTmC7dR/
zPMyo1S7JrjjQuvkq7s6ITTHpJhdlzxJf8/6ugl04QCz1ZUXQ25bcCwsF5AdxqR6tYNij8gjY3Ew
ZZx+8M70MtqoLxAcfSOdFf6PR9/kojpKFWUk9k7Cbw3l1GnBNlrpavNWH6MnkGpu5w5Eee0q2/mG
lMHD8fM8aomoPhkw5QyLFErfaad0wlO6d7tSdZhkjGsVFCmcjGTurlphi8rV8EEWuyzWxVMadTon
T/XKZd690aFM4XcQ+qts8DhqPnJS3H/Zjs5RMBmeuUSWzrUY62kEaI1yCOwhUCT+BWt8gjnzwBvm
34yrpFdczGhPAkOBcLYS9wOeHYmGgs2BJRrkr+SXnqjw6ega8CWPTD0MvqMZlKII0A0rmTTpLd5e
bNvNquBF1UahSG5Ri8Gp1UbR/xP20RuHFdmtKvh2bpbaX0A5fafp4D8MrWvSBkNCWKL4O7uCIjuA
REdJ4e0HZ4jEngiP/n3jeVCqeQ5dbWnbN3pT7Yoaic1BG21OdZtqSE+JiTceA9ViGcTGpOMVotSP
Wbk34VrxgSIgJTAZKAGV1leF0bf1iX7R1WkLMk6b5Oqmme7GZGT3Coct5p7LnyC0Y6OaSy5Ydreh
kxb+CwApVVcVR06oVFfyMcrJHTtaesBa62YXX741U5dghYEUVJaAAHpLPY9OG+lQE8P6atnInAwm
ZHYxMNK6CBDu+4/TaUhbhiePRQSgVtvmqr1bb2VIB7+jNNUmrI2F4VdscOMR4Olpwdlm+ZSalw8v
Bn2z87HMWGvLhEtPO5QegE2pqQ/aDjTJaf1Piujto0G0C/qerl7I9msNcQfWfLhr3s+al+exEoAn
B6x5dsypOrbKlfNmuiS6lCgN7GOiWV/AVGetj/msYoG4jx4esvXwAAl9e4CDFIBweXAGd1uodxjf
VnGYqmN8v4bdvoHUDp7iWIEX3BvbgKrDrNKDsASIj2QAPQfYRp4E/aKHJyydjNjzDxeBq2uHd6t8
OMWmCySYHBdCbDQKZIxiKRwXnW2kvVSwk0mBKZfBZ5ZJOR9W5qWU47Jr07miTo1TLdfLwDuDN8JH
kr4NRkwH4Sgrnp3+5uKMJyGUU3X/hL8WHQoZYUu8q0FIXjzxqe0X0OuLRm7pVVRAm1nDnCIKKUPp
SECOD6KF5S/xKU4kUUbZAGwiksTM9PbHX8NsGd+LZjtJYs4jjCy/3ECsAPr6n9YXLOej7nxGK4lk
wZNoLi8n5lzDELjjHsHuwb6FTVCBdSExRnY9wHc3n+lstMVcWv9DVvoS8xREigVrnjH+/n+CnJx7
IumelXEFrs0TiWkdQQMAwMvC8Riv68yQ+jZskRv9Tk17VkJ7uDfMwvthjLwXnoZUL3MwRe+V8iZh
jLPkuMoLm3D3zIkVpehQs2edp0Qo+N7vYdyg7nD3XoJkH7TIyIMCrKqgL6V0m9GHriAVBIeSLGTm
IUeufcAW6h++aF3jrhA0TqHI6MbRkX/5krbnQ3Clw4JfpSEuEEsoW2m+irRGLI4hs4FL/+T2DPu1
b61Xp702cYTKA3RngrJdkMsjjFx1FfnQfOVaI0o/MN8yZf9a55mqr4koPK3s2iLVL2KSyCfj++0L
Twj4ahq9EA2Ht9HJr4Ok2xK6BkBdGxDTCJeICwbwCg7MN5A39baHlnfd3kr0WDAiQCwcjbY4YPZp
bOe/7czrDdKagOCIK82Fr164De+XD8MogwPp6WqP4HRILKYKdin4+cOt3kW6qaStaUeuaKtl2Xw2
n7zKsxAxlBUUYRJqIUdsDmhSg2jlTeYAeFWNv4309CPbZ0zq2inq+lNpWeCDB/Dn1dlsYVwaN67R
VdmtIPLW4hFiCq6Bm1pV/H4gi29Zbo6McxL4+8NqA+9Ax7aIho+hJbuJlrauqxo8D1nqoKLOf39j
yHNmsVmrK6r+tuT8fMtZSpoVbmVuBZFR5iqAtZ7xl/eRsVQQHgnZg4et+Ws50UCkcA40PNN0/Tzg
zUYLqOu4GCL0MaPyQyeIuu3VZ4EY43TYFfDNYJJbAqqUiPBR9hEWJgxEwXpWjBwa2+Wn4BN9iQed
lwgX850NZ/AOox118ngcrEmkBLJ7Wxw14t4ZtKH9j5gxQ3dnRxA16kuRNBDecKXMUgaonxKPKxFS
LU0ino0lh87DUfwrQz4tBsov7cv6gfeUC7mL1179odwkFBj82KbLXPvSnISBKRyoiKjPuNRdAL5o
xHIX7FkGXXkvgPmQ9EvlIGlgjz8gZ6mhqnPHkISO/s+Uuj7kHRW8GJEW1GhdAl78ru4csC8C7ept
0+kxBLbf/to7b1Vc7dlAJhuF/D+jghjIQmztTSjM+qKD6PQEylG4z3wRPZ5oTRR9LGrparS1B1Gm
m5mDqSa2UjnA0bAVpg+BvRdkmWiWL3HUHljsAUqY1tY422U2bbQ73l+Grxi+Ym82QYALF3/RYhrv
+6JmNxXr2wrg6XWmSKlPGvF8bOA8y4BXmuV3jUvNIE1jnxoQaO7mZgN4xQGNON799AiN1G9v3iBW
kQ1O+xdlrlSVNOCSx5xfy6Nj53fkpvTUGvsj+thFnRyIAaYLVrxvh9KbT1N2OOmDDv32sfGtCYnI
w96vOI5RMa1tDcSmCn33t+n/fDNy4HTM5ZhBSddqCIFkEgYNoBNuYTbODHxuj2CNP+UyZdaveUYv
vNcbaZl7PzVAhNWr0IUouDy/de7oKYz5dzyv6pw/7QQMrYkCivvOvRY3RyGZcofkwEgKMOQSOIbi
inqswYzAC8ag1y6Dr8VDGuaqreuaeWV29zzl0U4zKnN+Hh0VAGe/T6f8ZEqOv0cePTOzE0Xv5gca
aVswND4WKLKdg1yXE9uJjkBHzJM67it0+abmOSp/Ef1xsigAdepRrqCnobrlprwsuTuXmbsPRIeu
MfiPAwvqNh2y1FbhTGuvEGu3uvwq22n6ESoSioKc7UdHpk08OAu8X9YnWm0zbQHaceard7Xii/q2
3Xnj9C4Zpk8UZq9Ok3nsmvK2281hoQ/PGeT+GlZSYiYc+gY5cBKF8N3rZVkPlUjMcZ8jzSjlmuGu
USiClw4ewaBDP+bMqfzBmHL7fWjztpuVg1spOgxVVYIwloWEV2rsD1rPh8/d5WaPhWE7mbaxclr0
zuxkuJ6+8kb4XIrPswCfQPb/BfEetGtDFKLP7GO1axtQEvMs7UaxfUuzbodJP8EmxDnW7Bxnjfhk
ieMkItV0MNfiqm61R8ziXLZqBUL7if+RSv6lx0i4J/PRziTGcV3wBSbUsjs+nzbVP/lk+GIv9Fgj
KMHskYYfgYLZpKTRaGTr3BOScqchyEteS4PgtcKb13bp71Pm619k2PQUoV2aawNwSru9Md6NjQxn
N7YCoRDHdyVISyJNu3Tx/Vg2bnCAtfPfGhrHAigYfBEek5yxWqLUUnYlqBpHoAKBV+e85mj/w7+7
MD4bw1WX8zDT+vL32DtOaqK9sWXhWSxqUYJFMBSSk5l/9S67qyuaJiZJu3aas6ravKNYNBbOjcxV
aVfBTrh1pX5vB5dO3qH0neJPFeSejv1n3o10yOASGqLtDsuwJa5LCNFqArw/X4PFMJ9Eu8923H7u
iSUOHV2axEhdsP6tpB+PZqwIIILPqqFEChrA9gPxyCBOt5MMpz5Hw3xQMS3RzsiIsquD1i9/bAtG
7fAYmfkRDAhkOrkI9mDOLp6Dcay+VaaUi3naYF2SgmcUmf+3xciZM6fsEbsCt6n9GO1qIp9rvDcY
2YLXdRh1g29LSEia8pt6DeUqIXVQKguCSeWwFhkWMsx6FeeamJpopLl52NeEvpxaUxe7Bfb7GRWT
w81P581OBuSC/q6GY97pFA1SZ2Oo6VFAw7/oyxooHiu3k8+YQcHuc3CnCXeOlINQDCZDjIJE6OU+
gZh/qes2Wey8Ub+43qj09TC9wdmpm8LGwxDLOEu+seUYq9nZo7j/aX4N+MHHvQbOGLF+Czu66Oku
zE0wTCLxpyEU9mtg5uaIig+tQaFvE/ziMmUKHPqzSawjPDfXKqe5u1QsboOBx7+Snwq/0YBpPyJF
3O22A2iSojppZlGijw1iaua2q34qsD9kmBca7Kp9IfqD6Wi2nJ4vDLrAd8LC7LZgbfK0MJ9eaKdH
l2Y7Rf8EXhy4e4/CLgIwjs2swlSc3SMf3Ej96tV5/QntWRS5POEhtKe2zAr8nQSu+w6sZaxkfcWz
o3XAD+l1YoIWZFz2Fpk0WZfbfiW9ZLllQMlH4ylLm1dqkOT6QiUKOnUYJsGfJ3N1TN7Dv/i3h87x
W2NUBtyi8A2vt86Y22O0W1DvbkPPnAXLzGU34IerbnczdLJecipp9dAR6rxqtSt7O8oK+1AvzH4i
u0HyNMXaSqnhPT5ZdXOiuv6jj9RnVWgkrTDCeTfutg97F27m8NDx/m7ukGm30A1ovE6Z3s89YN09
GpKkW/DT3SO0K1E4PHhOsIcdBJKZS/WOrGAe3658RkMrDAP8of7c2zjVHj8z+18+/NhzeiWVxxER
ASh1bN9W9p9tlW0EEmniv9gBFLdDkUCQ999vuJmUbaXN83mGgkbisGwFop1Dsk3QX3etWZ8Bl7Nd
rWrxZz4aEwkB07QeJKXMjR3RnVRP/Wvk5HHPxmpJ01i5i4iw1uhZbSMOpXWG1TY35gtRzoaWHfY7
6XcQNJpl+BSJ2Fb+iRaBMVEfYUzbTiHaMs6C0VWdDPFjxzxFmWNUG92PDz5Fue/V119sbxeoIRxQ
E8BfsYYlSuD6Y0fRBCADrD9b2MsbILg5haUWqunZaBuqbRh4cWDSNWLwfrzqMeNy1FV9eT6suOf1
TsFMFGkz5+ZRiOW0AXclp9YAlcC8asn++OCVPYwpdI/CQJ1z56bcxxqqXsHBHLBG2E+uLB1MpuLx
eeiNqKAYrWlURmoGAFpFCfs2w0Srp87ueyZlEW/4iRB6CZB96QIfRXzTyRRXxGbFhnv6OFmur1eb
Tj0rkoRWvUhczHhv47QzrqUM6aGAzp0RoPHfuLlIG5NGaboMnANVANNHSaL+1iLtu+YD7ArZW/xw
IZSl2lrEeuyUR3LA0XIYCwaUS81OW8Vsl0WJLSQj2+bIhJTupGNaCsE03/ruheaSKh5nZC2CrSZw
kly2iRVLIwGwErLdEPjs/G7Wc6oGwDwXcFhC3nNNF8jpZMgYkKhjds1caepKAndmtAAN+BnqsTns
9r6srBLFomMfrL5RoXzdXnOoojmgS6HRXXo2Bua34gChWsI7e15BX+Y4/j3LV1wyrwH+wSCGnaoe
kHnyM+2rhi7gaBjfzotok6+SRPgUph5aiAtl8lAhWZR+mOJe2QPe4ydsF9qmBxVeomv5AJjVa2Ks
hQK6THKLMxW6jNjHHzL4rS9UGV7Rfyxp4p6UZ/Hw3cc6Lly4yp1V6awiizreh+/mSxFCGdZclrcx
ADFfvX1ektzPC6pdYOY6T+OCgvzZZ0KsylRfiNlgvWZ2FmNtWfIBP3tj9QwmnOLQUJPE5eYJ1ipe
y572mVY9jXfvVXJ7XuJXrIcfPknFio/L5CV8bCBr/Ow9cZrB3yHHtwwXYWXl4iI/GKideWRIeqRT
b8d30Fo9wfpvzV14piIZ0OmaKQ7bIB5rSyjSiiF+f2xynrjHf0u6km1QA0UiYocp+hUN93ClQTq6
B09rH+aReNQzT/FUNBC4bivv3AxPcyYFSBgQUJ5wo6ZA9Q4bhwY7nt66mejL5uq9PQea6arsG4+d
I2lvyzaRurUKgsfMM81RDnFacQICTvodpkash2e22hNJXxu0ztRmDlcmHEyypBu7QdVM8kr54Avl
lPE8vqrKEof/5Ni6JYZ8MuU2z9KGz902QgX8/+ggIYh54yiFESAgEdi0dODYt6auamq0UHQbasue
z5i8VZAgpNNNNjl8Ww0MweKT/afGcUH2zDIg4Z4bOv+8KCPRw71GxT6BnP0wt9RWdgLc51+hMpTq
7VEuMWNm3BNIU2o625uwbBt2GCBNLNyFJoNy99qYDR4blIcHBnjC2blrmi5BRL0jWsqW0Lhuqixk
G6d45E/HDtvzsfxM3mtR6AS1pt+j/1D9dafX1QRBosi5moYZlXg0fabYetof23ny9Dirq4QWOtuw
dwoK7wY2tmptRx07l+ezz41aGs7juDn8/eWC6SlDBCr7EMKRRVkJbELs9ERJXHkd95gEAt7QYvg3
WogPQ6mpmYMAONta9zeSOUxqhaD+lnqi1bm+YSi3cS4me4JMB+e4KcwkPW3yHFATdq4YQ5e8kxrI
7ABo+mMGQyZeau26SYliE9y/ki4VkD3+mLsfawhLqsCRZASQEyJOxZXnte4YRPeyhhB7jZVLIdGi
ZERt07FuCHNdrh4YaWLdvh9S1GZGD0QpELWaxeuKeFmqPmzVgS2KHuwOH/+zn9jSP3A5dkWi6rch
KDRM9Z7wz4QSpVQTCNdF1Ca9mGD3nPiukdP76DkPjwDsnkJEXFM1OyIVdfjBRGePEVo1TkMSSEUN
lSjJ6mfsuphtcebmBqNDBKjljM/Xke7ItOUhPkhXlZRLPlVDtoCtiIA57d0FZJxB6SfYqLsATSur
vfyMGKvTocuyZEXbDm9xlYF9I1W1HlEXi5W8eqnHQCqzzoedxzxGFCTmGlThK0jgqj5rdGhzF77+
pWc2I3dCExRUQbTeojj98B/C8DMRdgfUfFZC/lKkq6w5kdids+fGY3qTWRzFdYIzKgIYaVSs5XbE
ArrOpa5qyxpZCae53eDLf+7Ud8Xu4CgBJ6BJJE3lbMhBJAoTZjT6mbC4CqhMKUZt3rJq+q6vwq80
nHbkTsD6505FEnqJvhKLkBzF+uM1M5HY82POIjPEZ8wJqUvzw7BK1hXliez67KHbbfFeOOjfPev2
AU8IhnSdEiSUZlMOvYlUloRvMCK5KK2AEUswopNjCZh76+Kiphy5Fc2tr7b9+yhwa8P/XGUkq9z8
3wL8gOkosnBvnSWSKrqp5wUk3BaOZoK4npSTa+Wwt3CCiO3+2OnRDa1qlBZQBtNfvIbC/kooEty8
deiAgblNGp7pVtZnS2gEFOigSPBdONYSWqARjrdlyOmbkdohuQXUCM+yXe1s/g69zkjx7nIqfDcX
0Ps6oJKzEHrCOSwbs967fmGG0Vk3GH8jpgvHWtDMAtcgHcimFVGal17QPAyGZKV4N1/W/6bo4v36
TaDH3OnKxvDK+lBYbDlSMJsoQXFLrLQ3VU2JgRhqMEG1VB3xgcky0dXFqKzGY3avTkik04lMiUo7
yBQ+85vjUlOA94zGZVnHHi9BoBM11+ZQSv2GggPlV09b2CXIgaslZKRc4RI6NjU6XZOUU1r6H0B3
VB4Fau9zOU/BeJRRs8bbTQmsb86L4rpQh+mHUbQAc8JGkb50kAbf7MlLZAOsCn7zioHKwfzGBZPi
/J+KmO3EPtRPx1aND0GhdZzcF0xP70s2IlAmEx6j2tkj+eGbTqwB5/bDrIYdznq0Pijz/wL8DP1Q
Ex6Ne2dirC6YuhSCj54rAW8zGwiLUmCoEgOY4xvTP6ffcj4VcKXCjVdcGe5YPnp3MqW/QrJYdbil
qGZaV5PXC95dDT9Advu/J0xV1b7BWSsrIeRTQxSqmMkJuvQyPSYuvJR19Y4xMHwkq3AGLEfUzO/3
57wH7GPb2EL8vLWG6V2IjMy0ZQEkJSY8gUrkeisafx9nqVKHApXn+WCuXNwMksmgN9YnDv+X6LcX
9DLRDB2FfW3+0PXvojyIr1jZ0Nd0KkCLMs+tK2Oe3UcKU5mj0ynrUueRl74DYknqh/pBshH3av48
c8voUEDIEosI6B9ZdjkyQf6SW+w56VSMbrMtNw2mo1vkg3g9OkVYJ5t45uIquFkpWYP6OXaka1D4
GyY9x0S+Gv2lWwPHbBAFSyQVP0OhS2k4znNOkwM4x4oNrcJOf2/q3MffiRaSYBwApYPQqvRvGW9L
fm4jeXTwzZTLOUb1O78BeeMcTpMBc12Swzk1aMDvQKhXis3L4N1KZEjaOgRI+Q7xyvjJ3NI6QxjR
zPPNA1nfdxsl2VA342WOs8VcYy8LE/YQeRz98fBt7Y4ZkqYYxarjFncz/d1FiJ0ChKU/c7NfoEx2
OiXSoCAP1FtYXN59vG3q0goJUi2xZ2J8uT8Minm153W6NLIkuaLHXnDdTYgzGmpA8E/ntXGWCdz3
9hp8dEuqJo6JgJDFO9SFxG1J2SPIxQFqOkSEvUzXA4UMeyBNmOiXdqxPGyrmuwioeye9k1LrCO6Z
/fSyB4q5uQYBS0hRuUXas3NilarXjDXGRKWawAR7yFWgATHP7/FEawQ3ac7t5SyePJDtu33vShEN
mBcKwqNcMPVS6wjmadcI/ROc+ofP3aM6C9wwIjHcW/eObQGnABBtXWHLrtF1ZCnYxY6QnN77/yQe
hvyf+k/1iCA5fZaZTXfKyMxFl3gw3tqNNkHzo+05Trt1wlqqUzaBZOjCjbZCw9q7eyibBUsTLIuj
xc0Fa3qo+J18B9Lu94RiYmn1MiiBaQ8Y6EvCXm1q/aa55M8tDGy8ZN4+hwXSR7ph44XplYViNSJG
9VfPJEmm+uWn4vtvm7Cauqs3ucqqQdLibXR+pJH5f6/r6fr/ChL0ocSBw05DMnPLMoKDpPcQr3Ir
p8z9ErW3XMjwGB/n43J/W6q4Y9hCCYTFKhESIpErL+FuxWP0ffGk3VSlspgmYyNzxwtS0i7mbWh0
s79mZokOSy/hCyPsHeAbUQzYXd68Q95tVJDAg7q9XqyT+2GgX90DnmtNv0xDpakK0ROfTin5EP0l
s2vOflLuJe96y/SmYM4HKoAeb+1iE3TpwGYT7KYjnMbpLUtB9fa+RivMrrMFr8JxtpM2CdKRag+9
NseqF33Ux4Lm7gTnST0uhknhdAQsdAmuXZDw0wSywatlZQ2FYr/vs1K08k3+BEVEclxGmtauc5dn
IJcC+iJ0w2JKsMhemN0ucCx1JgkGk4ppS7GSOLb2JZo9PKkXFzhkZxepYPjMLONEsfgzl9Srs6T4
RboVspGcFCRC5vyM764msiFqMKEQcc6PDRag+ykajPURarXk/0ybqk0JkbUi1ppS8iDB1HAF/f3n
lueH7vCxoDp5bIFK+UzN2dqZIsG8luyJoL+E6vhWcMG/jLjT25H+MKrhz7ExsVy/d13cKMwog9VY
cH0Q5p5bLMAzPUuwPachg2rvIFldVERQnZT1c8H43FWfMEScXXVLBoFBSMY8UZfqqfqsOYChVbU8
T+c2oHVRpg5YlY6ZtCxkN1nFJ8KayHyK3yEnhT9ML7uW5ywz37NoLg01Ixo23CQxf9N6TOG92ZSf
3vbnrzBjfXh+2/nxW8nS3/kCrfUmtLgHya4pLDeKl9uA+EUI9XjMkeUGF87kVap+CGDWwcOJUAgv
8N1ox80neMMkFJHRidcy+dcVuVgrPs2zsmTWuT7MN5ud3F572FDtta2+yHWJ3AWb2Nom5eCXSD9K
ip25gN6mMsuwq7Zp+jnppjGfZhuYyzkZYLbhwPj2TYoyJZsJZnF6yG+iEFCHRfJSglZSp0EIlyqe
1Eu98m4w1L+Brx78E1F2qvmOsEuFs9SsLr3nwdSi1A6Kfqjmwod5cuaZTmVvvx9xeAMJI530hXg5
dwvO5a0aVqrf8ygH6eYAN09zOmDpmMZ5GFoVD10jTgu4kdRuXGd3nuLrDyn90r2QPy/16BYHWt8W
/wlA9ZzS2/oIn9eQoacMbVtjWJM2IM5l4892+Y+NCW56/N/xCW32eMym7hzhGF5TAgvo9BzdZ1qd
uwFZVdhUg2iHqp9zed4RQyXVgNITPOH3JWyqOk90nAeTB6vcUwwDMoQ+Oh+GuIgCJSc73gxJuHTD
dDXmNY2iNMsoPHE8ODQ4PXtr+wR5OKZpHqdGvI+cCi0S0obbmeWEO1C66zEoQsSJkDnX8KZOUjYp
dguwhmIMvBgJRqAuav/EvykbVECuCvNBfrup62ywIIGGbj6Iv9e1qxGGDgvxUpJAKSXlcPheVm3L
QUUcNxZs1qafTT8jfDA55Pv1NrE4hS4Bj6rEnlHrJ0zgMNNob82jUAzVyogRTRRLmuUcREunIIqe
1J2hb7xdO71vhGG061zgbU41AWTHZVntNpLF8O7FS1ddWtTUO7/GeuT3LElmCUApC+YVfUmBkUkz
bNSQwWS6CZLz31/1sZLUWABQ7lyv6woUe9T93CjQCQQs7uVb9yWz1lJrkv0YXnN6znyqB9uzb2C7
pSka8S1XbsxX9zPMqZZLQ3ozBkog9PaGllt1Ig2zeQ4xM989rOeITO3t6wJqM6i6GFVJe/JykjzO
uyf+L82O15Q0Y113RL29Rn/Ofm7oppvtmilcCiJlbOG4xM075ZMYtziXF6mjr5S5iYMbPPo2gDjq
lh8tyDPYiO238O5UX6fjDGhfyiDDMxdtbEjLfP/HE4z8Ru8MxJAlqb03YhC4PPb2O6Yd6keArikI
BIsq2DfFFXGM6Pq/8XCEpXrmUIzBp8/uEzua70e1Ro5x80ydw3Q7h/Nxn079tzl+vujc2KOXYb0Y
trij5rErtCUDGWL72hESlqSBI2rk9kcFdfs18E/0aY71iNN3qVuXyvaJytG+VqKSn/DlMBXBzHC0
x1WhFyHlFwRZOOH6ckYtm3LEq6zbyhYTBhjWVAueHL6D7nCyYsiXsiYPDvPFkkE66yYPaGhM6dm7
rwFwuUn9evsrMzxgGcvUXMaOKmadKXyWG14s0FjMKEqYllMF3e0wz+bCDxPOv921HiiOudn8+yYD
GApafwOOUu0DkBRSKW3MMvniZLmnqJhW5AbZmlkv4+0VXyin/KyMPcdKlSQ+pQnCYOhQ/8UDvblt
IyhbNZzneZPTTsD4SicVR3+TxFjNjFSIWmkYgVsqc9U5Dv6wfycdMrKoBgWtPccX37KOrX0H0SXj
z2EcyuwWcYokCbo2SKkVyK9B0JrIYSZtWb6fbx1tUeUG+KnWT5APSyFaqCvh52lq3IZCd9TaEw6K
m9PFz+2ckbB7o9NRHXUU5vRZTWJyAPSFDmraD3bmUg9RMsg93PlFmvVIBcYE8qK1FCIPeHU4m1zJ
xcaoA2cW2jCIuTmeeujWN3cbCrU6zGqzAwUm51Pxkqi0Gf3dEhfPQZeIU1m7/8vzpEHxuyAXEfYF
VR6DATUfjcrwcKO6fqUvbpxZ3lUyBojKsDV9OEqvrEUZ79ogB1CyvaeQmAy5jN2VgOfXTUljOLqH
rJ+iZvkl6c2aFgpitC4ybIPqguvdJPs67UJ5WhCu+XAxjAhpvAqW7trPj8DiBiiVMGQe9qOhnh9M
ilCAx9nEshSav98h+kJ2wQfoI5ytuYDhJull8OxdnM8vi7XI7qxL+lQ8TdYexC1gaPsOwGKI+FRG
yYYKTJYjZxaIEM3GRgeBeeQrNIJOqnrDun7ux++tCN8mQqefjzX06q8ADFYFuaZCKB04Vm7UQ89b
1reAhBC5zvSuM7ABXJBsZBoahBaEGLKBE1WTf9nuxz8jBALQmPhRDVrX28iXTOLThoHRlbKvkA2Q
X7NXVT4xMQ3iHDfTmnTVbCngpdepoWWmGxInTDh3Az7RLUTnlZjucGZHFlemnhOhR5CvkPd9Gv5G
klO5ZEAP+a/fE2nQ7EBLT7LZkrXnqqpVnC9iofWfZTUXTdqVwqmj3lN3I9KUO+8DHnAzwHCxwzgE
cHvnGC+oYM87TvZTRzaxGBIdJ/8Lilv8IETM8VV9PrajaflhW4nmSQhptdQOtq1J7RwdOqpyflZl
WnJZXThjuD1wnBgIbo+Vkm+Fbj/GDHoPsUcIlqkjBFUYWt0+/lZqlUSYTzWh0xISXWPayHsRixbB
fLprDCN3at6ynisrgZZTUipF1cKN+0luv7y/6Xa+BoUEKigFqU0RzlBPfWqJwf1kTsiQmwRyT/oc
h/jEEN/qJjy3Gy9f7+BXPSUBQHJ1cKGu3kVO1Xz98mlfDqeccO+8al7cRm1B733ifSJHPx1kDTXi
84rvGRI+Jirx5gQouBoCgHcpxrDjxHDdOdR6OPRRFzENN/mpzGPVzBBs58BWiJYJFvD9aAHL8exa
gm0mmAg7LawpsL+uFIJL5uYKN35Jp+C9bwhYGkuZEJejqKCt/7hx+OgwgJh88Rg2D1kw3JfMJqQG
Tf1QLjreL3nKqIo81JIyn5XhupaoUCNmCExlJNMHoLrEmJX7KGPaSOo6A70Rff7853zYvT8IRjCb
d30lzCzsVNjvHhPnYq4zReovcznJSbrN88iTW820Ge4N4qdBlcEsMvkZlUrAZ68++2XY6ovH9d12
E9vk+1VH9lVdSgPqDtxT/E1kcgj0LSmiRiT1lDMnYaRhZnOfrM/tD42OfBe+kl6MIbEr+cn+pPkD
yN2yIRTyIbvxJs8K1HzJUoes0cr1WPkkYc5tESCDxpYIykd1z5zbNwedBVew3wZvxXdzDYEEeU9r
0cnvIAOnbUFeiwiFHV3jdj0jOG4nN/uv350CX1i3lWYbrZgdQjFiLOw/MU6Q4fOZ4CBljE22+fvE
VSI8rsvH4oJCuR2p5cmsPU9ygbMh/f1eDW3n4DjnSo9ia5jCe2z8+DIJW1HjxuZ6hzGQ4rmvU4YZ
bTB23FZiea93/D0N+jo3AJgy5str213nx9SNalwKvCtCVumTbkMztcXq94n1bTeswtOlFZ3Eie38
60DcKx8yzGRCC76Ea7mjOV6Pn0k4VCDUWEhC4ApCWt3yD4zu0QLq7Kkxo8peo5/9/9JOyOkiBbhf
G4PeurbWpqz6DRp0TVQg+DPHJl426LoOEni3ZYAto7BhQFyJxfObj/tBiRqCbm7Z8lCK7txZu4yB
IDp16sNdztpOT7sdb5FXecRxl1uqV4kTS1nm4VEAlFbt6+489ZqWYvlLk1VNqmfg0bRiC2rhINc2
6fF+uHkzLrmRK8qtHooFoDAtlxUvAULCBVPOhetbZ2nr3P1pZSGj6BjUpA0aBqryfM+lYR74RYNr
G9trQnHShQUU1h9pqas7KKfV9i4Q0Jo6eMkpEQdYnaglLacYbctYrFEV5RMtwW9qUhU1GgCBDWJc
yAiH8C02tKbQOmBSYSn1x7A0ufhcmV44CJdMkCwb4ZFUy55UcwR7B6x7DnQbHIZWTTJssrHL3j3b
ojCYKn0a33MMnNJNqbqaXjQ5wnp3wg4waT0LU+1LOCkY2kfkUcOugkUcjajRkOhzx8qexj0AZ01b
U+NdJRtHzjm1m7XGAquEUvuzKWn+4Plokhm2hAkPC4wTSXjbWEkcMAoeEC8zK8fARC2rgAAlSwax
FPm0rJsQ+9vLRL5Q52zdr9lMNZ3QECM6HoidU6R8Be0m3BUlFZ2+m2Ied2tgYG07AyI5/pbtjevY
ts4SQhSoZrvfHPQtHnbOxoCZEstSfeAwYmrdK9OYkFYq4hU4uQvNbFkhVykxxP5RnWhH7oewnA0l
4dqT/QcvT+EMakL8YOmE2+GguSLiRlOOgp70U3EjGQw+Q0hBb+XeVcIcAjP27nvgjQ4do3yBXB4f
LJusRGRNFSyUIGCg5kepPbxUdnKi+hqKTvi77rXzqA9hNlqVTSbAXeQWUO9ALVKmZFIGN9CxGUp/
rTmvs/CUtl141O0etHNCviEm8i0EwM7GCGdTVODwGKOqsp6oVf7YvM7YHzCCY9qq75Eubosn3ApR
qn+sQTUNAiT1+4H8ZnFd+xfrmvXWVB3sDIayQrUcInCVuFBGnzr1qBnpYtxjUJTOzdkmIizuaCJr
MdJLQj4HMBSaAVTtqheKsgdmh1AmSG0enxPeyDA1QmHFUh1T+a6umhdmYhmmCXvw0WdTf7s2uU8y
8ExNbOJ5dtglAEOzL4CUTCaph6wrAouTAWejfxY/51++qm4JKF2Pm5C2PWI/R7JnqVqrPeMgw7x+
rtPIDyj+sEwNZ9cMBQc7LmXGccZq8oTLphynEMU7qO6+ouz7bguMQ+e6pUiTQ1Ucp8FJeVcl3KD5
iXxJaACAnIfsAT5uclI/sY9PZ2WyQUL3fKjxNXqHrjiOEU7BDvuepX1+AZn3TxGE51fCugcFbNRY
V6Il4U6rsCv3VKjZfUvjMs+5GdtuR3FXZ866yvJjXKPU07wNeCgFpd9MBVfhz12jYZWVRuO1bJie
uzFidiaQPM1XVWCtDVkHKRq+ytKbne4dXKu1qcti68/nxQMQPgnOHT5ZhsBcyscKE1bC/48oAWzT
Lk3nMn2K0URxFeORiiyJrZ6Hr3dta7AM6B7eg07hJBjUDQKrhsr4BX/kh6k46xhuZFz4l6ZkP86Z
n/JDrqmAKWEcNc8ylWQEUA+YRMn2DTYbLSrRMOT0ISBvzrSMz+gg320PgipgQE5ApGjlro/a4l7/
g8SkQ05zYR/SJb5zq57G+J996fSudQGxMmwExAsBx+9gu+YR+RkDJQYCIMCSKHA5KqHWT7/2OdR5
Hub4l+dVxUrOdWin+L8duXhz8CAcsYbl00rQmftAf6CoSSAb4Rd2/5mZdJeAl1g+uhn9YwrijGCb
Cf6ul4igSh7Nni7TTsfqfWXBOZ8zIM8htBHrJiDl08BidSgMhe6x8AsRSRACkmnmTwRw0gvykoxB
H233aM74PdMUdnO3szLIU4h9taRcy+6SvKwBHvO7D+QUPPvUzl4BLrjS/1jEkMxiYZEQqGDU1kWt
LWHje+LdUe73wHnjWv29pggcSkTL3ZuQkhQkXDb+95Gw9gbg192TTVpylB5F6v4T1+1iTAlS7d+N
4wFpgApZYeO5pOk0SF+6dNSpVEJJP11unnlAWN8dSmoigPP20TBlq8/Czb3pG1vnKjPxWRjY7Ueh
1ONDMo1c9VS7MRMBfPPa8zXQoz4fs38BhQRUNjxuCqmkH1GQZKHXnPTadZVgEldbmjbIkDWco7n6
0FnIvknRy/ieondJSBhkMDy6l/bpWUffUJzmT/2mf8cIpCZOZdV9o6LP8FutWxHWKbF0nQ9lXFEr
zH166hd3VhFIvAAOXcWMBqskk+AajDtCJARC9QQMm2RLYypoCq95AXM5vuorQTUk0No8zHq2S831
Ahrb6ohLzMu8sLnjkO5H6tfV1kV6sR0s3oAyLKPwKs4RMovLKhHxIvxyoMPGSjZRkmtAaHnS06yb
sAEVqoNrxeHM9odKYfwEIUjDGdj8PsX5lxdyMwyjSXXPlLfNmw951T7j+b7DBfDE6gSXZGBBCYEI
RfZ5t1psxMCQCxA47craWsaHGha3YeHSDFz6YuFUwohXXYtyhnGiF9T1FL5d/yPPFV8dRVzt3GfI
t603/0gHesE6Vsm913hhLb8uys9Dvma28AZXTz8andzPCRKyx9Fo5rX4QaY0ZfaeqoEs/jP4fb2M
XcvRXdlCCk5mfwWR2umqRL/eLCH2/DzCZMsXf+giZN6ETx4uYmPGr7JZm8CW1SPZ2+cTDu4xngDW
T6GT5qLrVqZEfhiY/8EmlyAgX+sB4+Ht+TPQEGIrKtkaCzyregeK6zQQAh7/FzsoJ/+kwPn/c+yc
eZsC3gGcIIkH+Ws/sp0mjcujEwZ9UtK6BXi8xDxUsncdDYULB2ak9kWpclFUJO4I7WQzxmUHHWdA
yobn84G//LPOXEarmTLf3Qu6an5IadPG+nfIYXvrfbCHL0U5ZdlPKQ03ZzLZNIaF8UAof+h8sHno
tsrI1gy/3e0cp7OFKtmUjc1RmFO4URxI/jG2jT+OTNMU4KuYyIsMukSS2eP9NWMFzPVdtlKCSqHy
9MivFVUsvnJQnJjBuI9tJJ3rrTkPib5oMpaGHe8D0SOWp94YGxEWydilmodz3haC7bpV0qEOI3YV
3eqLhvsT0/q/0JlyqW3uU0/MWcbK24tqqzxU1M/+d/vog3lKfIlF42DEKfZbLXoAdSI9yPToXnLj
nfcKQIYiUOKa5ma8UPw7YClGE1YXfPxnGrBx99ehA8exKA2tWPPyWPO+5k+N3YpvqIMRA08Y0FXP
WEhJZ+90nF1J6Ur35qCJNPEQKuh86eEEv18j1SaBNKgENuObeRT7i3n6VR4tAZEjuVGDy049NKjg
BxnvEmoykbtpc8Ef/9Zprfmg5ga+HM908HKORIvePEYE3zRkLnTaMcia59YSaOnsAhL7JeWl2g+a
C0XpioGHpHR1jtBIQ8IRlT5PBC635i3FlxStFj5evwAWSDN3jFrbbUnko4ZpzCRuIt5ukIngp568
NgXQ1nw8/JC0aU4CQKG7eBqP6UC5AQMf2rVHC0G/4TPastZEhvOn5m5Ew6xtxn4wvMYPsbfeMd/z
lqaZtzTWh5W4EODDaF4EJfOHnImd3Z7oxppzTU92qAdNJpFo8H/HMRz//Q7+2RjX35pfMiNjiGC/
E54P0/7DbrLNoDLWKv/5xHuCas3uspPxDrEc3aVdgOcdDygNvLGoM/gl/sfW5NKwV80taqykn73Y
yRY12ubtZAQzIGQpnPUYEW+N8jsVXnEH9P2XHnVjbczjxQ5OJ45EuPxnT6/slC+fE2k2VqrKzPD5
4W61lLu4aPKTzQ7hdoRaaCWvPFVKzdCUE/+VMWWuWx9mavQeGHC9i2lSkcioH++Ka2A3mW+s6z91
KHekXgeLGcVUxcVuamjun4MI1UfTmeY0FzjG8XdxCo9463tZtt/NX/PTHdunVkAPEiZCgk311Nzs
WNsR9RLVN90rKP5vBeJ2qoAQg75oD5QOszQWSY2KJn++1U1LKIRWzDexBzeX9F76L3VwfnWeRFON
5ZwKxEVlY3LCSLfJWLAAP7IE+sFzTkevlDTnNwqg+VndCvM7iowBK0REZZY+EEF7oAuQ45JIQdV3
g8++mqHhyX1SsMnnpxRsZsnDWzvvmazymJiVTfrxbc65W8BTpA19+40YO/XEbfN5NzGbiy1L971E
AfRF48TOTC3oaLozjvFMygVhuO4NU7lfXsl7RmXypsBRdfobpH9ovBXt9WScKNNShS2hloToyLId
OWLhu6U/nNy3K5C9KrZ/x58xi6/QuoAds5H+OCWIjgbw9lyQo1pxu5+ye/NsMQ2v1bgWzOc1lqTb
VfnGAznF4359Kp1pzaWbn3HY9DQzo6SabLK665uYwCozeeEcOYVI/zhFjSyi/T/aHg0Y4T1DlzbJ
iyP7ZS924Emt/YHfSUCRCGhfFX8j/CF5oQWTEJK3TtgX3HQZqdtcpYt2jOG690aVGIgs00xHHScj
620KiJgKyx1UL2uDM5rQD2P3Kgoib95k7FcRpZ8lGlq9KKJlOs1CnXDmxoGXLSNnJ0+Vd5VYCzRH
m2BuqHbZFFkIgdfQFnbfcCYqfLooGu6TZlSQ3xGt9hGdcU7w33XGUZllPzCn/y2E6uAQScUPrnZ3
RCWb45dINZpIccZBPhwmcS3wZp7a3Z8+9FtfWKfG4ZsqHBt1WRVlGGPNiR+a2MLTPttEjAr8vp46
sgOBm8qcHqoObQzTw/kAQyVMhHeBXDLhBud4lc2cb/FQf2TxHU0q4NakPZJpwdcN/c16LmWjjAsz
E8zgbRQ6HyeJYTXnTYaXdYjhe6WRy0CTVscoTcCfVzUvNlva2RupsK0Xn3Pz9dKCci2NWrnKMI/Q
Rkyw2EFgnopSz7zfcZxAaR5GGyjoms7jtY3j8Q6cpI32PgPttUPDBqEos0kmORC7V4vp85ldkdyo
okxXgMQOjRq23EnnHyWsDl0c8owgdneietIYYvK6YmM1ENz94QrYhxVgHU1S2KejpwGpMcT5hn9n
hNFUJWMTpMZw8SLpOORpy80bW/DjEeRJlm7a2KKdsCTMLu1Df7SMggWSMyKPpiHl3BD8yTxC2AuM
y4N+ZLXZghUNJBj2lgACmPediLqls/Wqrw0KcAs7GStgfdyWEohAadfWV3hnMglsoz0ody4e9FqB
pcl/bDdLbcmrPPhSG8CBtwQAYbsgHTSZw1ctKZStEmQw9QExLhtEULQJ5J2YnQpXii0BXislhN1W
K1YGxLre8BVDlVvkCyUSLDLAKtoy4e5wmtCtcy8jTaWpoXDbUb57pVQAcZ+a9m5s63pYpPIFc6WP
/Op6Rjz485HKZkoJh9XbB4W4n9nQOzbNRQLJCLUakOBz8cH+Wa559oM8Wa5o8IPg203AzRkzwmBj
C57VH3X+Y/Vfd9IhCz0cWm9IeX7CVuxS7sdco/Xnrbp7ho3LnZ57zFb4K+hCnRgI+5P0TvAMkmne
GSd6H3D11J6q/hj4GXekQ7iRtosOBTa1NEJuzcoTEJRfW7n5skOTO5o88cSlzPf3xwW3NBKO1QQS
xwPMVLQf6aAg9cwqmmEiwWjNCv9uFMw5nhSPDYi9HCOenpxBCZIx6SpwUELnuS2eJp+Nzn9soT3Y
SlEjGLxLsWnlawSl3OVQJtK9DAseSb03jkpz9Tlgf30toNu2RqgKoKwV66IsrsdnHHyVGdR8iGSX
Yl9pqojuZGnQL2rJa86gsuFKy3uTCVG1Ut6BpggsdwrJmut7McWGTar61dcXXda9nut7e6v1Ikrp
Pk6X7b3D2ewxT/NXZgrk5Y8ppfzunuWHvekjd6ROxkIJonY9ZPYgMWpkX/v9RhJeihEcFmwAnjtb
FJP21JYopS+YeFKW/M7MDbJ5+A1iOKY48TQg8TUmAD2QWGQPNlt1chc9G2ZQaoq3OC/wkELXMF9a
8tG6lRjvJpmRKzaTS00NMzinkPHDTvQ/8YmhYLTfn23HlIQdgyyIhLFLA83Kzwn8TiegMOQOTg88
krcROzBn6MLJocqzb9QidF8TWy5uwHd7NhzVw3M26N0jlMNJ5MrJgXDt2utBwFABUaCOdPAHKE9/
CEHWzQDFkoTBAA8TMa+FLK/+tOFaWmlNFbHw+Ah3yusi3snfAlkZB81i4qUMNgP3jgkz7z/Ua6om
pPcadIliXc0Uk4T1wp6e+iHjNBHzp33n9FIcbb7kbLuhx68lFtZzJia9VS6t7dol2jWJ5/bwlIAo
uQatbJOHaHeGbD5/7BQIIZVrOXl5M5KqXM1EaDtFFiVZNT6ZJpt8r/iVm8M7KpG8YqC1rBuQuALI
tzxljNNS8J60Mo6JvQyJ6oAR+TVnvd2Mo8Yns2oQi/X6GM7Eo/aN/Rv6REGhpI/P5Wi1+ksowecW
VKAnC4n3MpdoR9UaQiYDA7tiWsTyTmtGMSiZQCEifwDZlYakepTMg2r0SMZ4owE2OSajrbquqpos
VKSFmKxOouLwkPgmsRVGS8MVJyDJkXIwbckr24k2qpc02bnTnQ9uYcXIDUOTwTFrRmlC+1B3viQs
bTlDngY5FnGf0IK+CrDHmE5Ocf5cWhCQUhDtKTqOiC6TmiegrFVepR2ja0ej3Vk11HNIKMX+z6q8
d+zEgeclycpfcZKDSEJrNau3OWr0M3c8g4pkg+SrJrV7HHcZijcVlo/gZimsY/FM1MTJsjKJsj5p
VvlRYudEIoRysCF0x/4MKTZ5Pftj2MY82POKWqv5Ge/01eLPC+A5ZQui96BjXF85lBuI6nZ5Krl0
KBq7By84FeURIMp5x6W+UfAMP14jGhplVGR5gltGvIiCtjN62Ok6PwqFzmSGWUuaTB7nr3DpVCI+
TKATmXpova/akIAvXdg3FlP+5r5XToOdMKdRDT+l2TFZCcYiMIlfnVKdOB6z2x+hpy23sr7VK2hI
mLUVIKSEv8s3rrEHvtKgc+mT0YJEp8DSf61+9LAscBO+pQiG0EWbZJHa7fIPImlp4gEzDi2iEMF0
0Xak6DB1/UcoDI6UmTgRIUI9bQm5jeCvlo71dewDxX7w1N3m5baCQgd8H+YLFtm5zZ1fLjG+xr17
nrvoOGg3sU6vKhRUHGZXYDs4IWWYxWZPygviAbqfFTLO8a27mWGCC6HRRDl1MVJ3QTmxGmGA/P+5
EPO359mq6BrfzFBQ0OiYNyiydVIWUL1uekWlzUE+SueToSSiTQsHyAUERWXGpeqkT2UfVzoePmjO
zXsgU4DDpc6MIxVzQmxZW90fWreLUAmJl/Ct8AIud9aZSZescpLkqJcBgot5EQwFU6sbNE5XQpYN
UPOyrc6gFpd3Qu7VOudlJ6P9Eew7DRP40vm9bVwn9Qt4X01paihqPBJIhUL8X09lKyBiZ4rYwR1G
VIKkEOBeo+WS4GO5ub9j7SJO7XRn/PrCiGV5WU8HhxdH6kZNlYCYhLV4mWSWEXBVj4DFOlqV+ni4
F0s0/Ik1f5aF13YlUFM1d5ROj4q/+a9eC0EstuQIArLh/yTbjIuiPbFVxUn19WWLwaOK4PEvrRAq
zo1ksyB8cSV1ddJ4vvg05HsJZrWbdWRvRAWVtM6QByM6KLsSZyO9b8A6VSbROhkhN+ma+XwKYHVI
tMe31gxoYS4sz7V6E7h2YgPqtMSBEO4l2KpVAV6trauccY7MT+ex1Ud2wb8cebtkSx4y3dBOCxhP
QVv3SCYkEk0nLOsx0thESFPNVJX+NaJH9j+xhPMAyn0WQADb9giG/75jVjAC8I0Iz0KahPVHsb6o
9wyEcnhCpWtI3Dh5i2DpzEF0jt2cWAA6JE0FLtK3BCGnjLpwhWmMJjWb72AacVLPnxgMg9zFLd3T
QgBNfE7mcaICEk9oKx8Efly4HHfQFq+gH0gRJjaM/76KKCf4X5yl7vUSTJ/+UprUExKE4GEK7xfZ
fdFQGT+kdvDAV8GnIFDSoW9zSIcJnGD9WmjYVzRSBtSI3yRZjcM47ntLkqtPlr9Ir1rlexXXNR6o
p0kSWOvua81GlDbibhDWqFJitrZYzHDl76ApLcze5NIVD5OpS+OAd6lWgDw58ittC8Qp2O2NpsHC
AnZTDfS1mm+03PX0aP/TnJPGWUR/5wni0BXG9rbSZLHIPx4a7HP5XiWiqfQRYBAbbUKWceIZgFfF
Yr/trEjFQqwhZwxmLQ9W1195O14eDNeRt2TRFpQ86ZQYwAnnub7nYxGgsMXeR2dNKsH0sYin1Ro3
yU9WJQuvYkLOSk9VXtT+20E4wKADY0T3YNxApB3BJ3HJyyCETCsl2a+2rmIMKUAAfvJCACjVYK0k
iCpwJEVq/1mAeySuMgO9QTl2Q1w23VbruSITrWDsh4dmCDseimw2Z+s6cbX7eRGKyes7qr0tDE8o
ztsGdPSzxKcZNKUB97gRCXyHohYVfb+JsgRMVF/UfZbJUpTqCGqwQDjAxfyD86/bnY7BwDb2Onwj
gC8k5Gg8GnY9nTCturHDLxVto0DHp7R0Fdm9K6qYpStONMCuF8EoYAEp+7TZBqWOeMEmU7egz6NJ
t+AvwfOvtsxNmBpW5UyY15H1OMM5IgNqnLXG4fk324H4OdsV9Voujd5u/uA8fadCw/a8YhzIx0Xm
j67VFD6zjhidGTkyrybIFSHOufIoUaXgVkzPhL6c1IYGXEmzkviPrycG2uf9Ahr3WKMh/aiXi9jz
DAOVxMpAdMeLOWwCCKslWzx+7mof/POh5I+0zNIKuEysDiCtiwxwwe9EGNXinpUzx7K4eqQFGJbr
ZeyKQZ+c/FHwnVj2yqp4TZhq7OCsqfOK1N4UffC5BcpC0FIFKzFy9nMizlBhJohFEyrjMSWC/eVF
BAntxYfUHgRvNodkRSycpcqJ1MocFs8ASZT9THzp6zI+fPNCbVqkQuuG3TcFHnUOMie6ku/OdQvR
kxcEe2hiYcz1lBU112opvnkg28FAwPVxV3M06hEgXOh/9FWemMixAe0ravP/eD+CDqUezEhGESBm
ZMgZzlGNHPW1sztFvv2nU0Opm4ejpUK/vvUKj8f5OxAiAmb42RHlqn9hGvzwSIi0uZZN/ePqsRFD
AcEiCB9f/GdYJps6QlgIwSQG6khafVlg5b7OUWbM3g8ZW5pw/3JR/IPUg0pVaD4RiZcEkARqQ/7M
MAOnXipBI7IWruJJlGBL4Oogn3az2qrpI3zNm2UNhwK/uI8suVz/tDmqY7n44st41R/zhjV3+w59
/MJMrRPWPcc17i7zLwddcm+VGYLSn17L+WUnbuAHuyEsfktyIzRdjdRaMb0fFEaa84Tz24fqbUJq
PzSjKOB9LHw5sJ0LutLHcQTL1m+tKSB+yLVmFi2OvMRHJC903gDBakAZy91I9PLcjtxz3FUsuLIX
3rWuAnayZF0/wO6JDxvPgTkGMItJHS+X9NDRDB8DKmvO1zl9Hgu97mnmMJGCWHc1FFEVT0wX0oOF
B8hsfI3vfYv87FcOwFhOElc9ONmkoZkmDsvwBjKx6Xx81Kd8TerY4kdA2jO4iXxBKXUnMnhQS4XR
7UlBATIW5HKwu5DEgTbQghmp3hYsdqeDpCGB78yNX7NOcd+RZ9Q4g51+lG2498NDrMFbkHc3ncys
mcGt/opK344+QFMjQCv+xwxsljFeB1YdcI0l1lXVKVkUlT/9FsBaWwRvlpd21BcbHmrv4x6bEGav
ldSXq2zOM3o7Tepum7QDEIHDa9qlkEfigMcku+hWc+91gsrVcMt6VpJ11seHJRS/gRU0u0PdfJxq
L5TgmKw1OtZOD6L2hqcBlR8WAT5qm9ulqQAel6spf062rTzxaYylC4JJ7Deh9+I1X2f3kEMpapxm
oZM0s6c1VMjtXoGIvK/5G5WrQoZxtCnlD7dRg45a8gWHh4fef9SOItMqIDFW4brlYhABVWathgeu
zd7riAGd5gwshfmj7d0IgLsPr16fWWR5U7izXANE6QzbgcMYaGnOhR1hGplvJSJiQQp9DfsOyNWE
khiiDyLWR86Z4JB5nd7ffslMqjJYPlZpAvFhnLPAW1a4OUnceDPVeLdR2GpzQ9BLmvlEE1m/yc8l
IziLkO6DAy5c2ontZZD9Qa4vZkYs5QBPMnQ4DE8hfb1UNDOeFZo8plUWrpjLYe2QoHppDWRudzaR
yHAqCjztPfmPv66vbLMbdqySauMuYPK9ShRfobj+P0wVGPNQF1cvMqqlWtRYnIPQjZsePqoxdF2z
kITmJmYtWL0gCQxwVAH4J8BVgfECQ135q26a8Jrdui2AXlRT0RxQDGSqFCcZDy/RRU6V7jodhP8u
s8kb6V+2VvSP21o7hTymQx4EmxOPcD+OiqX+mvgwgaMMcVh7sWmAoStHrXmZP484E1cWnX3SLOeF
p6Hji+nEKzOmizzSXz0l9ADSw7HG80NENBiStcK3yvaF3LEeiGaJPqTNrN+R9viggxR6LTD9ExTN
tTgoqBpRAvjMTY7jsA8BFg63gbs/YKBlM6uxidnxeKlc+dtw+mKiedz4TR7AF30HoO8mZkujRe71
cNJ7MWzDlC7jlGzz5ocENaPzF1xsW8GjJxJdbKQ5XMsaYbI0oTLzT9JtgFOpQuhDay7kEc8vR7jo
SudyIuQtAUbrRWzX4/NM0gUfBgsivYnShNyx56X81fritVB0BQ0ZyPSNMrW4jD5+gYhQ4G23RUcz
9h/Wunb2trGdJjgZg5kPegS3HZkHyFDe+sSqF2q/tsopXGs+kyNcH0X+osZ9K4HE00Y2Xll0CHwB
5j44x4VIWhxCRTE6oFE9UnPBSr57cANPMGFwlv6ljcBX1lqSu6JHc1To62hD4zVQmkDKSiL9MO4A
pjkUZ/86h8oc4WJLIoU5xP6deBImaZAP33nMEtz5Z08YJqQDKbbqScd9vVJNZCrFKc3v8w33c5WP
eaHOY+RAG4vaiyXfRROEebDlFXSHRZsMlx+7CNtvcZBIbyJ4HFn/SO163fvZHGBSP2HfrxA13j+j
11qjp9cP/QY1AfMNEorVYLEGvczhf3HH75nx/qmPdc0PQe9n8Mg9IFvJzjlNHYQ95vvHscAR90CK
1FYlGPqyqCDBgSmvmTZYk5G9gr1jmX8u5OW0tCkUwfM7rKnDNIyTOh4Z/uiHrHyijgZiGs9a1kfk
c1Tg6gTIwW6IkYy8vOFezYxHk64Oa9qdMd+y1+We8XcDbw61VoMo/XDuHigbv8xGzdAWb/UPQzGG
iRmnY+bEBqwuOt60g6g2ggIGXpYB2L/w3R0hlkfuNuSaw0vGWMjjctPM7doWy6vEFge9leCW6VWh
6OhWVoFOd1gwKiwkX7BB1ShhSoQwb3vcHDxRlrbhYjRZ8Ne5vd/YtU13STRTA8gu8W8eb1LqIQZ2
f29Xh/JogW0wwHyzHZCgge+qDpAPxA4XSuiZ19+9MQ1JiivelSBQ8eVmXremPGn1k9QmU39v7Bls
Wt5dcRNPzkUnh/TkqMjexEScf+e31bGP7n7C23lX4WS/f5ekrdH4PvX31ZIxLnlXArUm1BWz/Y4a
ip5Or3mxShWvNkzKUIS19BnCIGrfwo2vj75joe0bkRMwmvW6i/Hihs4TreldO9M8ggEqrXxwpsRe
/iSMjUMdGTSxmwiIPYPDOiXnHdeRCUFzlrxGHves+bJ+kGKU6zTQL+kFQFLXH+jbjAaXklRwZjmz
+ug/I+eYYVF57KP0g8HEReEACQKoanDDkCYDykTS+rMV527Uy+YEHNcAif+fZY2w0gDYPsD/Z7nB
tWEQiW2wIRXBo4f1/v3xyK1+G00bt2PvARRfiOIkreOGIH5a5U5teRxJZRSpNRV51i7KQmr3cwim
1zPBjnM/hdSEjXGUt/ugNpdIcXg49ZD8eI/BJuiI62GgNme/e5c8qEq6JYsDLjJQLhe/3wQ3g7E0
alHth5PwjDhelAxHD5AZqayyb8duRKfwb9kZmkusAtjZugflt6EiI8t6f/ksHAU7gQmbY62Kk99r
1qcOKTFTAJle7cvtyy2wnQvpgTPYMIIDEJSoWMaW+hHaDXyi8W2olUC6YraRk+d96+E5iSQABcQs
qbEs5+s42ccCizn10eBDci5Le8iHyBttoHq1tYHIV4HBSxjAEKGi0+CLWPQxpJiDwGR0cJ80Woor
pnIx7v+e966csud7d+hW6hWkkYSwg3jmYZk+waFoB9XtB6XY5mKnjIB/Qg9TmRvAsdlfJgfSpUZx
T7ZJ9w/zfpCUp6GVkZ494y9V4FmSiNtCpD2V/3rKkzEti9CV2VkUiwsYYXMdIARWUTjc9MQJwZ/F
z9+IkGKZl1Rv2KI5NLUQtUb2y3mC/zKOXWUvaAJ50B2OBM5XjNlNjzCxJ+rmUSc28NVSZTMxmfyy
joWmGhy/R6g6jPV8OvdYu4pvzCdq8u6xBlsC3jD4W6a9ur8Zn6hOMsOAWde/ezRYVBfW0MdPPy31
N6DvXXObGrwJQdSUSk+wXEHGxxCqr15xY5R2S75yblTbFVKHnRdELuV+vPFg1Htrn3RCQhGprEQW
Cibfzo9Mq/zfgHUFLSmZhQ8ooWUfauDbvtH10U9tI2kF+6ZbBdYExqaaV7RSS0pnXs7Myn9l7qlM
bwVUfSYbfga1GwDVzgWUactem0hFGuezafqR7plad6N3gvI2ycKgAI+MSauf0Rm5tS69sTfvr+Nu
DcLNmJdLu4Hc4mHUxxURLvL9AeZVtaWNF+dbYV1P3nmf3WR0vAki8r0gS+e4x1foWIXggfZmevE9
Zsqqj1EbrKJntNrBDeQ1T5ALfyauCiwMUXExE4g1joqzW3fy1l0y2cElH5WZknM4bxMczibpIDtw
N9pJuA6yrLVqoa0A12C14j+dRURmbyBQnP9xM3+CVPq7NR10d+udtGTEWQEYxrSkB71PzbSkwgsB
2nXOkvW3N1ZZbKXWuTW7N4FgHpcPQV2hZd4Tf++B5BJ+w07GMoCioMxPwJ+NqSXupdOXSOIX6llO
DBVq+k+/BekgF2sg36B3itt52BxImq34dIUwU4Z9pWTaUIBiGUNqTY05iRhav/D04KBRmt4FFbb8
W051OZTc2GwI5rUKfdQ4mq3KF9uQaNnuhLvHUZBAMUkv/goYv0ZQN0TpuFF4mUBlGeWdGXetaMso
wQVA2PHiPmQLhCEu2EAsR9okTSkIIgQcdm5hn0P5KZj6dLWfQKtlTG6ffWf0anhzphI/K4I1T818
3U1j8Y7fsrm7TnVwyhNR0gzSzk926jbW5YZ2bHDyRedlAwbiHihxohQ1rYWJgPQYJi7TyQ9DBUl+
GgHGZfqRSYKPsbkoHySa9WIOp3TX/DEgW5AXJPn294n2a63Wsi2LCHzk3pFi3CB7kpKEVEgaSl6h
Ya+cLee7S81hv6PHbBdNLbu3L4dPNu2V8aBYjfFLhUGXUZUQMr9kye37I05gC8RJs0hpeTv8FfVK
ELwbWCfV55j1wBsIZgXGGKL/94NYEpkw4Za4imY0tTQiGlIveooX094kx7UvsE//WEMK7px9PkY2
FkbbzyYpemtSnRaJ2aery5qkJbZU+wFMHPFA0GDe3lwW3Fbt/ZI3E8bu/jBRExjokRyMHdqzqThI
0D2hacLwnGailqtPKwy5tl4EhadmBtliQmUcKxOulHySTcfoHZ/YnWrQPBZBiLPINvbhrXHZZYVZ
A5yBF10kEV+LvEgMQwGO0+Jf5HHGlCctBqUhVTK4dBdy52zEd8zr1FUzSAigjG1czRf504NSeOIJ
rJMabrSkGh2yQuvPxKWP0ZU7XrUIQ89oy3esAZLbAFKQPsPTYgQTz1fmpImj19aIz+z0C1EsV5zH
WrF1GBD0CxE90IIZvav7ujAOwSIZ8MPec1k27ApPf79HQoK2RNYKwAoOTpunVauJAobioZ8keqUv
8B8bxvpbop4yZCauskcwSshmLau7XU5QM7Yu0edevTuiZyKjjIPGAd3qPNeARXGTXbHl8Jod8hru
mXGIIRiM9rIIV+XmKoJWjNyrUQzeONK94SnTL6nQNoTVeJvbJj4nKZ1SvORR3LDzFykz8gikazDd
44xuTWTbxU7tsVg/NTR74QBNUjGVdiQDQkaXzlFF5W5OOE4zfQkte6JGM0iHudK6y1om/fQwkPrZ
w+bv3C+9MSKn/2iIwjYAmjDQc8KaQJv13aeycAdGvrr8UkNePwaIFE0E+HYmhuKw0mJAGKfWnQjI
16juUEFUNJsyoWHNBhfW1ZgNFhQfNby783vNp3FX24OQtBzeu1YejkUNwSQBhOa53mKBD7Grjp6V
tQnwfRodHN3Wq29VcUqdg8LkGwGdlmGV5PZzIxOH1nawGNYSlUg77TpPKJXNVPlWyHXQ0aa/EtwX
4RNTjs4eFt5ImeBeEjsN9Vr6Tpa8aK5+vAKvxFUZMQruaJWgMTghN5UdRUtA+q5MCu2RdQWAZVbl
6G2/1gdaYCt8FnDQxFwdHQV35MhZvye+snLNwsAbvZaei5c+D7LHcwpDdu95KqCUPhWvbv7qfEc2
x9X+ioZ2a1MQaoX6B91lbhGlj7YeDi6VDnNh3jUATVrj1lTWjpJCTOSfwFeMu/vHQyo7d9FroNHt
nnRvbZmPIELJhfSauBYj10Adj2yP3cV3p0Qc+UN0V5qiwjw4Rb4Tc8+ZyjInXY6j8db6lRghxb5y
TF+3VjUswR2AVv5tFVJhJ67YpqxZSARFpg/xfz+f/KrqizhPo/mQgAQnDEYGrYoQ2H6Tpg6YbGy4
9fdwkDisxiiDlMBhs+IIkFYe2kIaAhSNVwzcE0rSgHtcVa2gs2sIW/CWFbqfWRsoiE5p0hta44P7
BVNDaq+dxC6iKCVLFbVIcGCHltp0kmelxhlex188pAlA1cnrOOlcwW1pZNokCrWRjvix2qTrE//P
J5qz+NZmNEvbCiQc2LARJ4lt+uJwKnVwb0ZgKVpt2pB01CFbaiSJabXdZXJ7fXbrynEEy2c4r2K2
/wddHx/4dW68UWEoZN8wsBVdiSCMWnlwaYvPhbAB02tD/OOSO48hputahvGa7pRZfmz4btCr7K4P
QO8vRQhV/gxmgv8zwHRRojDeR3TFIIU6XcIv9lVZoRSSiG0bQW+qnXCl4WG+lHf6Nw9+7Oxo1IPk
3eeHJO11ey0GVJ6BsQBwD46+DkyXWmess2Uor4YQv6WmgM6AzZhE18OphzZ5ndsAscp5bX6gFpcB
ndvl/kkT3iWmceH97PGfgqY9+ElSB6KeaFuokA8hJs7H3qJQEEF3CpnRDEfzLOGfg5aN/RSXTNot
hmNu5emtqy4trESGXHP8k1GXkQixSPOmbTm1hEphG/q7RWu9oKuu+BQd6CNg5tr3xUxBjW+6G+xr
8iDE3CqHf1UUPW8xKLSIza/wF1QI+TgsRvmdkmv/fr4DwWDY1Zb9jXVa87owSmfQTOKx4IeMz/0P
MXS9Z5jgqTCWavY+U5IWULzlxnSgRR2LQxtk/0XvRqo267lI/6XM0wRnx5J7MNV1zo8MzonUyQtZ
VPuuu+3nPFDn0PfvcayqXzU0u9cmSTIwvLflsdbxErdB0By8lMiiFvBwX+640S9ZSO0DBzxJm8sr
95eN4DU04dQCT3k3L5tvYCKU84bMY1eTEhKIKqbYSTp+IcztSCa2r3zK36JtbeQ4/wre7LwCYd7w
8hl2lRdygMDSCgKR4HbJ6O4EWqPANeFJDV8ACkaU39cR8W2thM4yj94QNwjFl5VxmPSHdPBiLgvL
DNvsQBfKyNGkc4/eQriMFYnWmXYzqW1mRGf701XQQptMUr2Xg5D0OeuD5MvFMIVq3nsP0OTil2qe
pQ2GcVG95Fqp2k12NAS5LQt3bZlNULaKIR/mC467A2xbN8DlN8maHWE4uPllrToGXyanMrb7TnKX
AT0JwC3dj6WudY7zrWz+XfH0m+Ho/eeX0fQWpR01euMBmhSq0pjnPUuxRjPwZM6oOWbkskeb/v9y
X9Qv9eK4KtchUxH2k/GUmOpSReYKq/Tztq4Kd/NrHe2qrYZXhPe8wcHTWgMPxvC5ERnQ1qcCRXJH
femMguNZ1VnUiNAAd240kKEyYKtW7Ray+dA2jH/SWVIMOB6OwySE9/2//0dzmiZRoe5c4jC8VXEo
tTPeNaJ1JL92zoNWcGEEVrfHRBsPiawfEgzFGRjQG73cxGjeSuD76qvEbMUg11UcA8mRzGP4Oupx
GuRF3oC8t4Wf++MSjrDyLLOQa9P8wiEZroFno+xAmJEvtmSRQTuAz95tJ/msIyIJjhtB7Y0qpjdx
aSPCruyHKc9xc4NLvwF32pfucV6zPuL1EoFPAJLB32tep5ps/N8iepVNpazXOJznwDCtly6j+buo
WlHIJIFTVFOlscPVQtmd22KZJBU6hYLnODcOinCrLq+oMDclYzqmzsJFDzn0YESBPR/8X/ZtKHy+
lfArokaHqkFxsVxsBJcwoBDRcJRVVoM5zkDi3c3sq4DuSZv89Kfkxql8D89aXhjOUmoB/2Qwo9Br
h9E0Mr5DkT0jzoY524xECKl7N7c4NTihIaUwV2tjSMYh+8ZJIsYc4WXn5e56qfF7aV5gx+R5yOBT
9KCIPKWa+gKuDz2uYO0s+l0T6Ju+hWSiR4K76NK0K27LyhaCBhT+GjjAuCnkvDqCp5g+koMOybLW
2BF53QM2N3w4XkXH2YVoEyEe00o+MraxPdVRo+3vCysJaxNKjnIKv3Nqe9VzNxHv+6ns4dLFTVSB
fNdVc94vK2vtbu+qvSFxCEhYmzBUNRhC9jZhgJqhJffE25MBFSsQhmAT0w+htCviPuNQjvhkCeSA
1HVttojFAnfrfgAFEw/4Dz2mxJS5jER7G5F7gpHBS6JRYSl314UcMYeQ05gFCCasgSG10rgK72WQ
Xg7Ylx1KttWeAimXrwLglb9Z0O//G7C5yJWB7kJv9aC5RuRGQHpfJpbAhBFdI2Wu3foQcHu4Vp7C
hXEFPmtPavDlFBGCLcIYjDtmPFTTCnTK3IWEGK2Mn1vyEN4J1zYkJp5x4zKaygA/4ULaEurubyjk
t+qtevfmrgMFOJ7J1VGzJXRkgBmeVBIKej4cx72GRCH45h139C0DoNFWCWME0HWu1i2nW8921z5m
9E9hmVZRIC2sySXugDaUB5VwiSPswJbL7kvetbG8sOda1vQrHTKVL0qQRnuS/3pOnplfObDqeLfj
NbhdEAS3wOjq/JnsPeRnN5fXtiEnSZ0LNnhKCburhcwxreEJtjw3CkNyxQ82PiytBrVV3/vW9f3f
cDKKUg6SmYLznlwGo0gnPJFCXoPC1u5m7DSlDoaMQi+pcVdF41XciolFC4N0iizLV9g1WAu4MURq
BD0/EzyMKtrK0j9r7EW/QL0NZom21wCtXyQ+IHDhoVZ+RAQkHon5KaSGsZPrY4SwJksddMyFKd2U
63YTvWCpCdiEeNMIwgvlj0lfvs8pz646mTVRn8tT//b/lJLarLddwgw2yxhhDdI75HZdn4yq0fbD
xATbrLeuYMqaYch2qRsJtPgSSx37tmvuB6LtmTGFcxgeHtdl9hc2anbwaCnPEYMTql7tKA4DWJes
dSQ88KOCzEJYrXw1+5ND5enwpUZVzCqgYfD67geHjeu1+IMKzuwF/uBzP4lViTWL8ZV4G5Bp9uCV
FIEybITIlyhpVZkoh/7u14m5FbVW4jQBnwRzbTCLezdowFEaAwRKba3TvB4KP/DLkUlMWqXfbXSh
XgF2PAYFVBDimAFM6BSyisrYweRRFCofPpGmqtwodSmrtQf2Hyyb5rXQiZ0oLAHZHx6Xevv9hc2P
qakzr3mbZXKjO8+Qqe486T7dyN8kSxjpGHYRsathp3ynySgKN69YyFTvrEfS0TqscovPOCW1icOo
7h5IYkKv5kmS3LHQKIIUkZNC3ViE3rsn0dx7Q/rpjwedKu4Ld07euTwtEO6Vyhb6I7Ftk9Qye3Ze
+lyajBbJAMCZOnDaq3Zfqr2tpGLiWPGv1MVTh0lpo8GaPdkdFC0jZsXhqzJUuGNSvYZQ3Y84gFb3
rlsLBrX96hcxgENkyMQSZVuWUd2qgGvJFPa3Kg/GJxuusG6ztN3VHc0myzRW9B4AcR9x56LqAOnX
2FCann2IUHKi6IP3BeCLgmsHWP8igfv/oQpldLwxhB/qycA9Mn7XN9MDriC6JaSn8PO9um5mLLVN
efwL6Y3BITMIOyDYsLXnsAWmekw2uqHonYEYaQp+3YBewN+3hImO+fPMcs9vluHYzqoJNCqnIeoE
LH2ovriMIE8Fe87/nseAtKP/ILY+24AfurKCsSqvYtD3qUsgb8zZtnbe2aoV5WoOrOPy0ZkTXP6i
ltuv6KGhY9cVy45KqdRRphlwgdKP6b6wdQt+dk8P5Ogn4spRwqCQKMreI+brv2px3nwUsM9EjAMs
xggudFa8eU8WcNTmLCnxKES43KJgwvp22ajV4XmeoJLPMltqIFfxvQwCwM2J8EnsSmTJcUxvRqWL
4+ubVk285WZPe2Ctsx0/3fx0eOSgmgaCzK8HIIeEYww/2MEg96DjNSp/4u0fV1yNLv9+d1V0R7wD
962/7GRQQc48bc5lFrttHtrnGGJfSrAwqIBVBE52NbSdTwhWiqbF+25BOJLLMqcTrt2MHNWMh13c
PQX7j9XXli/OmvFO/lXaiXMW+CGroWs63h9Sjn+fJUR/2B+YZ8n/0CjeFH72FBQhco7a9hBtsdQO
5V8xNy7y4t0qiWMPNROLrEZOTRgCCezPUKKhaPcKTC23EspJwIVfdSwKRmGpWNBcrZ3TtAErJ/Q6
jx84OvQop2E9D1UnHj1ckoRktm+Ryt1HgvJwQrztC7LAvg5fW0w2FzSkw1M8lc6N35dMqxWMhwZn
BK3jRrnRbX8Po1/wYM3GN7bpc2/OtVmolYW+bq7Cl/P650c8Zdfdkj93gHluv8lXtCT0YZWKf76K
P/VLpRlP/2LO7VT2ShlE4Tck+dvmRaHSLbdTvsXRJmMOI5uJ/ZdFUpwPGSsaqBSQCYXRIsqsFPuy
OuEuvEWcGwpXcGe/wOrfV2XfUpHCS+y8WtLbVuYub+J2cCVl1WakLzWHUJj4/M6DV0kZiyYVe4tk
uPx8DJ/rymOqmERx+H5+rjnqokMXfQMKlqNNXJjoHZCbY90PvZ69ujToJ5ix0nyvfjOophNJswsi
Kp66sQpMjoxT7ABRoMiQ3H8R5C0iPhNs3d1jGWatEhDIevG+yHwRDPR5hRTCjEdHrGWdnwvf+W85
rXk3Uzsi98LXVywTBdg1/ev5Fgog8qTW/wzatUy3341528b5hKBkBb33V/2xsUmwx+3zxo8Vkj6E
EIz4nTm7AGxbfLj101mBZCrBRFyMIIA+8Bo1koCLA5zs5hcT66xHpl3K9AlqsvDJTwnGiEqfMx8M
8zQ2++hfo6Wi85x4YJCMhWMijDIAclB9uWtUce0qdI1euCDA1IfZ6a+N5qjn4pGnXgWxwBkd7H92
VxIph39paYKyEHSeS7oyjG/HQgap+0PL9XnXMzQMr2hU3w3V3RdTeDKbCD/NMTPEgYTbbf7yycq9
v7odpyu2Kb6h4yV7duu201qwvkW6GwpABxSZnMnF5LAdni5nL6Jxok7lZltHT99qg8+fZORuEMsj
FAKFhxLeSjFPRdVve39loFTWrISXYo1SaU6NhPG8q+stGQl/TZWX7WW3d5RS4aP4nPb8LbK5fsit
Z+rkH/adASc458iKhkTS19OHzi6ukp1WiikO4KFRTmHPHi9kOenS+uNtH19NlOqPn/NZWMReI4vG
WVlgAz91AnltgzzqlxyQJsNm7ySLnjvI3v5/qJEiDl3KUuNqROZ63mGLnVAwtmwyta1JwPGOXaAx
9hpVHlZdz6r8SNJJfjoLvbxwyVlx3LK0kczaD6wbj/V8jMM5OBiNipavYh/rIm9uiQ7kJYpqvml/
Mr5p341aAsE/3VoSZa3sZluTSbaq9dbyoMft+mSSsVkjgmMgKN0A/jOujucG9VT8rFy5XTK1ujy9
xEyxJ5LPmap2UF5kNomsVt1DkT5HJ7KFegspy46zVszqktataYAuji4SG0vxvjErKTYZ3o+cC+s7
C/YkdobhnFhkfXzK3I8LsmG7u9EzMb+hpO35k7mAc9NbKGFH2DaGOZQ/QF4vPEMqZmVM7nMKj/F/
EiwtuY5j3RRUiI75KSfIWMPQ2NUK8kurtR0mOWaOMf4vjPN8Smbdor5jvdMFbK41uZUAz0kUtmNi
lezCJwJCWrt12QcTyO7u3NHIRnZe/fyjBDVZvErqwz6ao4imGf2A4CEDsUC+Yl3VPMWAyftB5GGT
Lre6CUTEqE0QOm/ygXLoc+THJc3awIbqfcc0pLgp/ZO9fxbDz4ojW2xzsLSUDYLcVfWvuVkMBt4A
NohbXWlUiu5cQhnUsKYq9Az+JfoJA1JyD+nkXk1eGmDrSZnYYQe3z6GEsN8HSd+SVJElfv4j2cOO
Cki79LB5MtSxXJ1fEIXa486FO+Z5gHR7two51KUAmkakn78tx2f9PHKdsPCVry32braAVFvzbLCo
0SSLSen8ahkn+V7tVBp5U+Cm+cRiQ7DKBoN0fh43adaYoXOv5PLeZo9zDdhhn9a687wdHq5TvIXm
SPGF0ixTaVhpIkyoU7uToBAFzSK/syx/tGnBPqx8NzDiUBQI5QfqCA5lEuAGonld6Mt25SFKAcwa
SWMNZ9ioEv4fGheArPlHXKxqFTYZXx8WeXI7P8Hjxvr/KDbJvTa2le9A4G+5USsDZca3PxMNKOsQ
URh26gP+SjLFL8k490oGwRIcEFgroqKveRXc940ejrWOjIPuIH1JDtL2Z0myGEgK28YEz3YFkZHo
zlUe1SMkQpgerjJtD5AURu4La0FEIs2VuOx346mX8oA052vrCGAK9afUuU3Fr9avQIPMF8WkZfCw
xgsOf89VJMruQKf7tmHpOzjd/ViQoWIUf4JdvoPHFf6w5ik64sQg2DIk1H+zVHVQ5PlSMeuhZwtP
8D4AoBYWjZkJEmj3o0jrZAVJt1/tLg5GuY5hIs+SD6aSz8WBt37kCOgKCMBAqxv0Su6ILOWm/tZH
oq1EBRs5p3WubZrFJC3WOx4OuB5PtDCSmGyqK4UwvxoR0hwNUx9X7NnlCZaff4JqZBG5Sf+LATd3
6qoQVbNeeV8+K+BmxXlpqc/Od1wgqiBRnCbE5g9XJjgjx1qFH0ImY7mplK7Emuxwwm7ll8nOYa0C
66AYtdMNtIFKopMsubnRYRckAKAfIb6p79Yq7ub5ys80Fs69JAYvNtoKeHgKcrXJiT5Lz6LvNpnP
hZDcH+mYs28hc524yp6GrvM7g2MlszXwfvchlGxBxKAcLWW76oyyCaPLKiOSiDOJoHXr/MHYYRSo
inXrAQLi3Ab0J4fLLCJ+63BB/FmocygmT6swfPDMZyHlHkQ9j5POwBaB3Wu3b+8B6jme165hKAky
tX3OTtggNYWJHhndL3jwkRRj61GOIsHiEQtpzl0CHGMCKB7VMrB2BO+Ko18ylpmVeTY+2fkiExDX
wafOOfSg8KNyjxMdnUmvFNcmmDPXVbJQRsm6vZYhMvL1zATr7x7vr2IUqHc/iLPPOugxS2sMdpUd
z+cxKpGKEeP5qrCdx4J1HGjA8mG9CHpvmMAPmgKtm662LhBpDuDo4kJrrOZUYbfGsRzSF6gyBfV3
7HUoKnXi+q/V5uezufQlFnAYcelZAtJpniuTO2IdxBnf+ty28I27XYEtwS5PbLgFVzvwzZpd8qNy
UX0LQaZ79pv5akPtfOZKgZ/2YxhFIP9M+ONqqgS432L6QsOWtNuW4t5cCiytT3Lh0hDe8xsgvI7+
7Qhzx/SYalmXvG5MDmqGmh8J6OZKPTHb3R83CeBHdT2yYRw2kcyQ9Y9qDGSWQqRyUN7/BAFd1V0m
6spKjgSOawapGRA8v5bc2f4HlaLd0zVOdgH+7HLMoVmuymg8myBvhJ4HogIO7RI6NgSoH9cmotaG
jLSoRYPEqYXlgDc4wF7WrlWGJPJSxkusK1crndUTFA69+juX8CVgw+v2WcXaijxFhz52xJhfUshm
TzrhHCloEhHexRFzukMIB6uG4Jk9bhnhh5LOBjyhaLzlRdqrCVSdtMTFBNh6gPe6NbZKZMEhmlCW
7EWxlkM0rv5+GKsnJrF2050UL7AOf8EjBOaKrq62FiUAo0+Gl1sOOJGdmg6Dofqk7rgaRfsNgVKD
OfVissRQS+zZWuQw+y6tsKqd7jU3/1TA/rwr9Eh71ApMhr/1yPyy6GtSdpySgyz5+UcBErgM4lPA
LkWfVLkmR7k7ijWQqLYZ+7Tf2h3m2vCTUlw1+tt4pSR4d7DKA8wIElWojGn/80BU8MjBAitHhUD2
ZHsKGTubCg1jMRyZyL6zQVa4ALLGSikcHutf4cu4XDofWiI3nNvyNbiuHgrvdmvmGn79RUArR80X
SCZniYxO2zNwCQr1YADtFZCZJ+nHu+6YaISMnMGyhrsaW47dhePEe6cN8YhW7RLDpY2NELt49clg
QskCc0+0HGUC+AatYWftKnO2wGRQmIbD18cxyDg8572V6F0iSXvFdC79VeMfavgMajmV5vdplzIK
+CZO5Va9bDaZKBaKJ1oC2fLWNcES7Kf2nCqoFt4zeubv6hEKaaEFU4PZmb477pnH8qWzNei2m6oa
jP1TS/9vrl8QAA8AucRS7E6QOALNr4akwc0odzdjCTujOW1P+Wd8XpA22ONJSc9tyGq7zYaKOMS/
9UajL0/lDwMfG/EkoMHccA69QYA5YH6CmH57l/EwNR5u+OgGIMs9we3U+1LBo2xKkk/SmmWDZJNj
EOTW8fSoMvSyTZphlGlu78PUM6c7/E9VIgSaDrbiDX5EdNDybOY6QfNoKCsKh47LRyzSGJNEffVH
bAwd8vH+Pil/q/HW9hsbmVazXIIDwtcO5RfuWDRUbKTrbODlQy7g1O6ZjdGeBotN3HTfkDgFpWeN
6+UjJLqPmlRP3lcVxO3a5huq5kUuO2vPuVWucJ3SXVY5pem/88rWD+z58kF6X/lkT4NP2WEEmjXK
Rh9knb6mv6ZYSgWqVBv0PkIP596zlLSKIdCn+5TyZPjCLoV/zPRVnNXTPC7zKbIBDv9FZnZw+SNE
b/q5Ws3go47KVb+PAtrdY/Uw786HA5diDsgJ/JwK9qlNq2rD7Dzx7xS3dhxqZSKNNf7DqwzvHh6C
D1uhD9o6B1kFrk/VQ/4pCcot9A3834HAWl0iyMPDoVXIXcrm2hXIwNnhr+qZpdFA9s4gw921+m0i
raOL3p2Rd5+apPzhiPpFrzuiqeTZo7AUlHxWEIB9f+7PmzVeEnPFyokaaIJdim40V8QQ2WpZvO9h
k4+kDyZzmspbX6XNKTsp/hDOh3D7n4i9sDMWuPFX9UjAc5sOI1E7OOeNNT1oKML3C3Eu5Y68qCPN
ybk0ZLHGiwkDyf/9NHXfbhvL4iwolquFKQzy2bMd9jjQ0fU3+3f4JMEEa6htFz0mkgxOby6BWGr1
X5Zzxxc3ee4uUJfp4j6P6tWx37ikaDlfgtlL+tQaducmfD3JXuFCF0qB86rN1aVQ0VaUPfxRgwUr
otMgjRq4kN3TV8hNkA6mx/ewVQPwrzQQv23XlpuS2cokNFXlReLNxHyw5VkYlv2o2HGhbGUWGvEk
9RIfCwWmATdKGL/c7EHGLGjopudXEvXeDP+0WqjJt9gPuPxie7o1RN4MzjSYr9TYPLxuHXu0QiNg
XgveuhisvvgvqRSMnt1AqDp5pIhpb9XFQ2JJotoNt618VSTtfJCZV4RlIsElD3q/gv6uVaRXPR4+
7oM0PtP03hRQJHgJYTl7QDk7bsNxYzTxvHFzzIUavAfp7i/zRjQxPfy8YuvMBuYuJSlGkdGQAvDB
yblbQqOg0AxaFSziIEoe3aTj16sQbdtAmw8VIRAIu3Ll9B6sHtW/oC5PSflmQUW4Fz9PVzpCOzlq
PzSlpZLr8qF/g3cItPTpTacXbV83lWb/ZzlG3cOubW/EaLsSAp7fxlZ61yzuhRg7c2de/DD5ZT5X
QGPRnNKiyE6wo1Kh4emDsDRjlmP610nvFYGZFpsq6XolmYCs6YwvMuGORlAngTR53w4DHOFI6Sw+
szPlyVlPj4PgAfomHMWCQFfMkvzvOzB4CiZuoUd+d43+GRGFNcbJmwnQYj35aBGNn4j/tRhcl2dS
FFRJOjKhubTpIfj6rgY8BUPObzyqpLPEvQOE4iYfMr0bNXne1XUYlqnUu/0KAnEcoxRoze642IcM
IGBq6oidvAWDrGaltOZlpzUVU1lOYahaYFsTz9/mhjOrtz0BDhgIYupDuHrpg6imM0giLr0Pnq52
NlNlg11SHGCMjm/t+kaHRBdqpbGH8kY2AZCcIBvNhgaVLXfVt7QAKUyo8zU2Q7/+mdbxlB/Zq5Iy
onjfWmPwJGP1twK9Q8i3TmRuhYr4P4U9/AD5TMoc0CbBBflS0bYK6x7pOJJcmDOJTDmeUJfxXOCy
g3S/pCcvVSD4QZ28jqFfLZuT3i7BL9R1O6z1MwYqbFYo3Lwnd1tE/mSxhEp2pIA0HaM4supxM07Q
i7faqVp7L8SpKNkkeBolTDhSYMqIDkvIG/Q0v5s+ZQhdv793pZl8YV3TDO7iHjb/9iNkdRUfsJtD
b5oRRghK/NYQ6bKiTT0PhUtRSZychO/PTnAILiloafV5Z0ig8YQn2qDiauEfhTyxdbXInkW3Iacx
K4rFYieO6ItGk7anMP3LajmZRAzfo54jcJwQbN/W+GNs1Bee0SHxmTqljwf34M7ePtgLRbiraJS3
fK4BBrgM+CTqx+q99KKrshmr0lNqY8Xr7WSVvMe1PI0Il+aYkvI2A0xYOGM8ef1RwmaUwJOXwpNA
URv8J6P8dIiDfzv9dPT0PPMZY8PmE2vgx3DN7wm1MWC6fxFF4MdVV0GvaF1HFn8Tb/huTW9XaSlS
u+oq0vWaEPqBsXUxKl29xcKOfkkjj89s2OjPTfQrlcezhHEnLFY/as/5JgnQudMFPLgMgShX3YhU
V8/rod0thDw4f5cUo7sJWYK+eLY7+2N8XKIYj7H+zenlEtgXj41qYepEzO7V/lgc0QtAXD8CF11L
wRolFXTGqOaD1HoBmv+r5x9dV1Uky23tRua9qC8pHDZ+c0dWbScV3Sl/HUq3VVSGicIfzAJA7hvY
K4q7IfTxQBlvAqEDc0MKP9rG1spjkZtQf4fuF3sUYBSOwh7fuzzQ4cgWaldug2ikr2ZwpRDCkw8p
u72EJIYA7lS6YNuBKIv133bdymNsAVwcW1g1P8RzrdO/KfCDdK9opmKv2rU3NPtg5PtAw6RoN1Gy
MIvbhrPRXOvxqoOaYhfUVqSB5h38m+OfqLrf8eZoLxOhOxuOK8YSkppO/GLnxhGav1dzZWLRGep3
tnjs/QMu01Gp8fzijVVXUuF6adbata/nAp03sRRgVzGN48mhMYhJW6RJXPPHjB2bP4TMt8cxBeDW
bGypOcsQvlIFdfqjlHQnaDv5n/vWhaVKyHf3V98P6PtSf9c7SfFZsVhlESE/7k8OO/tny6t2TKSa
MG1k+ZLFYKRtFnBW1zKztPMFCU/3hgtNVfhcZuXvTDABn8nn21JM91l2ft1M0abowPTT7e80V2xQ
8yrXiEDJBYO5o6F365MPZZWk3mL8FkFwPiABg+7p1tPY05UeVDRxM+f5YlV24Vv1PgqPYw7C/mXo
edV76+zj97CahjllpYilptqzsYmFNF9CrNt8ThKXKlrgkYQBCwlaWUmnVeaxL4olrmmKAUuNurYA
VesxLN+24pzXW51qatQy7qkH04bEostjVJxq6cGDim/vU191f+FqK+sHcNyNE/LEZ+vkbkp+dk8h
poJSaLiyG0WV4BGZORo3RfiVUTAPc/mLAXav8jks4HB9zCyKSUB1MCs0Pj3pPgVMXjaMVHYIP0uZ
Q/snx7Ds3O8HXmL52BHx1Y/YmaR+shXvafyfPrQl85Bjos9qCZEs/B+iN5THAGx7cA15jkh6d5LA
lI1zTrE/zcEe9WhtfaB2LHFoJkg99OO8b7ZoK+OtnZJAu7oPQatP97Z4GWtwtLyoM4v8ViEIebpK
gGyZFPVUbDM8G9dg7fesSQOeI7dCyWS8G1FdKLXscFhzC6aRD/MyHiCKhGO9DfODjYSLxicN4dx8
fJ9KuyF/fIZZzlRRF+yC8oaHAC0g9T9V3xsvDLDAF4xbaiOO62CE++D/KCwn/rh5EYyEBdYNoPfa
VwjtAejeYW520k6z5rw6nPTt7RwbKjlEIdxNx8v65vxnWRAsihdP83Mm+yfcWpGrfl5k4VfJs5x1
3WeS+cjMMNjG4DL4xNlJBGFMUw4v9UpH1LNY/Lv8NNFCVcn4MHFkTwR4i9QcTzPK2iBPvL+9I83/
yzCC0mlVPGjUYXgUcACHd6AUyiZnbB+YvwxAXsbD6QI5hquOlzeRQ2TrjlfcCfEFEu4iEI3qvtAx
RGUi+GcvxzewRQqyUNIUdFwXMahohji0QJQ2aToP8j5UN9w/UIZJn9WVZP7LNZpZOXhFVTTYKARo
L6pWul8PIGA7RtWnuIU87XsDbQjDsezzp+VvrPQBkDde+PE/vfG1jxpLCneYq1hRNiC7E6GpnC4Q
ULS414f3SkFMKIYWPPKq6ZIOqDM8CQAH1nrd2E6J/lCZ8H0CiIXRkIOH7BeWtqAPWda5fQqhoU6p
p/n7qGxnKYwYUdhgdfEtQ4qSznUsWGTxwNbfcfjOOgFBbKc5oEBjp6S17ymyAO5RIrqCRge8Vn3e
F+o05pcifQoFeC9RvhW1HJ6Bf2XBrrPWWgrIRXrrfBFB/yAcZzcnpe5fwUhX3MPcqXgrhtn/7PYo
Q0ZU8FHuUpOYmkc7jIFMmAHmQcAN+R+rz/JgQD3dcIzd31ovXV0HqK5Uo7sOnlghXSJSycTGCL73
ES9khuuBBB6wJhselrMoMH1QMPDPyh8o7wwmS1JScnMdJnSN/HXBbaR5rQOpUnD1v4jzYBGaFpF1
P8kg3J67gVIpIoR9YF7ao4GNH1TyTILdOi0SYAJmJ1vc6oHq2mque9Hbz3X654Q3ihPOYXAvJbyb
0jY3rNONoJ3PC2/j/FX5CWzhEPWH7ZMexVOzeMM7CtqV13FH6+K1h73yWsnfmXmboGlCqS+zHWfs
HWs2AgIeajGMjMkyR5IIQRIh8AyXySovTiXm78AUt3/5PFLYQqAnEJj0wuDxG8nLgERIV1EyvZLR
yCyUi7ij8ot64JimMhcdpDK3AuQjf5OxoAmjjms4heYuMm2r1D6kzAMeqvt+pFeSEcCNyzYIFwPy
FIORpGTnRv3+LVenCMSx910T1i+mN/LvGyLYR/mTYVRzUHLeJJgRW5AMiMzgV4r5bNtVAfJqst29
1xJH9fo/bov7URY92orz8VYhWFfm0hbhHUkKMK29rjJQvL/StkSPbfxLb3AskD2k60Z/Ha7KAMp+
g/s9V8rH3hmcMbiXA7I419N4GcXSWlYfHkTi6RaRbuN8Y7S8VT38ALp/NxWeJ9KQMDNmgetrtQOM
Rkf6jzjt8Oy37YKEVdpSAtnNlLifePRU5cCrLyNmVzxGHktLG7UrvlTm1bwdfXrLeWPlGYC7FzB2
mMMZtu9nvtqEKUoHFTqLzWpUHtVeCx8hJhim1yZ2+5UT0jq1icZo8rsoIFNk9wgBL9cO3e4amiP6
bvALBCnd0KExCMasEJEZ1O3oa30gAZ2oXefQ7Jsy+npnwNJ+ub5esOEQQYT/+6XXLEIL+pC+n0+2
quB/HBwycN1Q3yQnjUR1Sn0LewWzYZmLwAm6t8W9EmQ3ZX9rYOzmBl5racsl3C3rqdAhNkklKpWU
1oUfPi5RqwRMV62edhH7qX0vWLgYU//2SLZZiGZntT+VwIDo1RF4OQZepj+GnUCOzP6ijpwKYTy+
rl6W1xI9vp/Ru5spKjwgvMxpWBRfOYWZPr9F/xqwsRcWZ6GkNrRuXV+OFNkdoMPsOBlqqpInZrs+
Bxs4nimxTqF6L0wCgF+EKB/ZNi2RiO4rQdkA6Pw6WWLyU/Q6ZGQjlFZJTn/JZb+aNh7DcwrHbaXz
8q76l+4HY4Hnhaq+WaYsEFO3mCPNtarTSupkDToDcjr3KCstG4h8zKsomeBsJFif78P66TddFI2G
C1bLQuxVycmWu2JMqfaDf4QaLtZIcflDs0R3b2rouRey0FzO6w601L7G4xW+vs8rEtncbiCPepb/
RkNZCnbg4oc1GAVVBbbbNPVAWEW/cgvg/tmBdGWEkNYTS4230hNTupQ/fWzfjIqYnh/NdJ2MfpUQ
i+KORqF8Q7LEzwZVhdV3GwoIW69HzISOP8IFJJ5wrBHaUuucSC+v7MTkDq77L/QdqBrZ6SvXViq6
3I2M/CYI0Cit7qothrFZpFGGX/tMQiIbfp2Pd4sKTdHd4mHh2xuTVSl28jotIdI6rHsrLbmzeKix
VW587Z/zIKcCuEkj+bLNyl1KlyM3q0KYnUGs76l4f5XYaYxpw4qQmiH4nmlvum+n+B3B1ClK3GFD
Pa9OFN0sGk8+89cBzH0mK011IL8XiCMZ/01Q6wU0/yXCCmkep9tMHUaMCHcd/8TflmkeDRbU5tSo
mwE11TLeNRoEp49LPUnQ+udeYYHXnxWiJU+ZzQZMHQBegnbu77Wn7dnDODXluvnhSdW/CS7SraBa
s3rc5Q8NszQwxd+5FHG+UDAlOJv0ICpELINu+noBOJBHCrlWdySyP2GV5vFyYTK9J+iyAWATWFtY
CbntaFYSkWwuTF1eIKdD9FsIa9NfEGCrIGaWHcpjUnCOL0RAqDXXkm8JWpwlt5/yiL6ue99dhaj5
KvTK1hFEbRagLVWHkaMhP4Up9xM402jaS3oCVx0O/Pp/X+bw5viL5PSL2hSnrX4Ua8PVaslNvvQ0
xK8+b4CL0Shd22/cm6zLi/pTcG7BapMrshuI13M6Xwm0UrGVo81WHcqsmR+DE+Ssesb6mbq5AxF6
/63lHv1EO60NhXwZ4uD3lVkxgSC9xuHLmowIg/qIVzeumJFbdhb4soBhVi1MOvs/0fH3g1FNwR7X
3N4uwpGmBSaDgKi5nowZBjqkWxU98YzMpcuoSr+T4H1p9CeAiF1qRz0RxlxQamSO/BgGiGfnPOXt
dsKIm5NsDGAvwIDtg76dJS8UF3jJbcI/sX04mpIw75YGlCYDdk8CtEcMRmYj4VxWKMVJ8C6+qpdl
9xci/tzCyoP2ri/mO06kCGRAAXxHzl9vYDWsDKRfBJBYAUATHuPIP0fbUDppNGap6AhkoD3IYiLH
rfMxa015AXNq+T/i7UDThkc6PmMOe8hNBl981bS3x7C91hr1Tm3tqVA4n1bhVrCbAcVWg3uSV6Vr
FDbZUDfRHjHxvCV90PXXsT0PIYtnmM0mhAjkwLVw8HpezzgLPX+HFE9DDLhGSXibEIBl/AUtgFcH
8Mc1/FqEVgN6aI8haz5UYmEtJWjVjzu2FJM/hFNi+nwjxD4c5zMpmXf0Ce4Y35LBAkQMMjsscFWu
5mjLYC7B/FDSFYaSbnc0wA7CCI6W3B4PRWhSZetJ4xh65pE85vigDmRyGJqyaJxDKKNI5878K1Fh
bfKlqEXCxHyak7HR7Th/AXx/gmZTcIRrlxqGD2W6uv2hHWi3ks/Yw9D65KcXzZjZh6iJf/KAhTU+
dORKJ0JFpPraWhHmSVcCRryDPaKM31Y/R7TnvDC2QwEbhGez6rMfsDH2sMcwBCRk0aBdbkAKt9a2
yY7ctDFkZzMB3TdwX8PRwgcNgnYT3fgjlFVxA0NJoJdBJhPCpq1fknV0iECRWv5O1ZO7aDAbh/dM
iqm+hYCP0qVyt2hSh6wgaPOPMsB8/4+JevdMn5ROxXFaWsWSQVhvepvdg5jHxzRb2Vns2Mx86RZJ
LibVWtSENtvbWQrif5BigrWNBfnwolWuiobdj7RZumzIDsfX2E/AKMGRMyz8O1Wxy2TSHmMfBF3N
fFGH9kL6o5nLLvTH33SIBYO4ya61emBlYxL4qL3A36T2Hh6NOnVgtnzFkzPFSeiiJCqQqQPzwK2/
jkk1tma82daixrSEMsAH82CEkwt58IYTKqrlK+kFT4XEc1olQzi1ipx0Zbi3P49KXS/WtjkkyxAa
51MLE2it1R7QDzVqnQAocvByU//pML1Wa2xflUTSXceGm632UaYpJQSNHJVnIISdzf9ZXUFt7kNC
YwLgWOfssN5F1Czx8P4HczlzpAVJb4ml1BuW+cvve4naeNFviG9O7OnI6smGjFnGEQfCqGQ/eHvq
uM3uTdhgKEoPrJ5oSz7DeVtpfzST1c19m3zft4dYWiD5vG1bMIgyVh151rNyxOfE8+xz0QDGpvNi
Wxsv84Gm2a1KnESPdB25cJ7Pbm9M6fXClCe7LlaWbHBHV8c35rQAZ9p1/zh2k90DLBiXpmkILIhH
gXmCPubYNrHhGUFVmjCj/ErXo9G5isyanuJD3fh5XaaqTrg/a+a2clRrUe5pvkmDS1Epair28wWW
NbpYM8kD2RGmSux6I0G2pwZVRgqfBU4ogStAmPqcGcOOWvS8harDjY7vKNmqFmkIrpdeJuBaCkKf
i1T7nxwBWzvi59fZxfo9vH1TAE6wetw2cnKVDkSmt8z7KoTCQrYFmV0j2xxSBrpqiN/3Tx6oGvtA
JWAmJEs1lj8xvxw/VWFZSIO40c9dNKXKU28m4k67EG09XZX1GVRD+AH0hIRaKMZlA1nlHAZjQmyb
hOl0eJjPoZF9CRhNZ7TODvHsYRXu0JrM1lkocv40F67JBiXDEknEw8kWCvbsyfzxtjc/jVfX+Vfm
oV71I+TORTXaVuLXhzr+/kOZObZsc39F5sluhPJK+7wJr1yygqDeQxvLA699oi2H2eSP1/MCtYKB
ug+UUL+uK04R44Aecn+9MYqVhDBWcfCKGSTpP33KytP6BWMMWkFtstsGSYjTxk8lcI4o/W7T4NZ0
Qv+V3paEXo4Py5uA2AGUCQKJUG3uC0lX9fMkxOsqfAQopD0EstyXh/n8vWLgb5KAUBd0AJuaoQLN
itPiMYUfLrb5xR/YxFKdpVi1RsNwHd/g27TBaGqHxXkLC1DhEUK8mO2Dw45elLKp2YOKKEonGnmW
JbQsNX/hwSGGa77bdaGwDVi3CVrds/v7MZq41nU8HJbvhhMVhhE27edQbLBMHzljaJCfg4DILJfF
vzkzeNDChKbN4lF4GXGEdFqwS7ZlP5oYjcC+0NhlJ8Xe8AP6mcTjFQjKLjH0f8nsBkD3L3RfK3Ji
0y/wBcLBBVi+tPWUU9OyETcXMwjbTNBnPz8ODGjfEW9SefH+IfVeDkNGYXnyvl4yAIN3pS3eV5/U
MDvdszGaimDjcUDDuv7eXKdNIO8qSkPMq3HlFVZNQi6JO9aDqq3ri+csAVbkA4oIDT8py8blq/04
+twsxIXlDPVbnPvHRvpo0GT0NxPTJD17iwgIG5pLSg9/WyZnoQJ8sbdAE2bbgF8nPEFVvZ2MNXgM
J2cgg/252UtgW2BCuHkLOo3o1IJBJTpXZW1/Q1T6xQgL8EppXIh7uUpQ05FO/GG7uqXb145v5Edd
HtEkRIIPrzr5NSOZnyKtQ35rfndAObG3dg0kCjzXabZrCmPTD+wqnSBG4/wPg4Xti+K5vjLbtTln
5C2RdCB3fYKY9B0hTOKfbtA7DK7GR7kWjwICRHMC5JeeYZ5/cn/P2+4uY4H9TEAb015DRECSy4HB
kx5po8KgiurQEciFKhJDW9gV/U5Pn2Gwuqe3/hs/v2cBfwOP1K63k8QtSClsARxCwpArV7K1uWQL
Hat0coj3M93BlYpDTEeKwXH/zHPsN0DlTNE2y1uOZLfxXqW6CiVTlC8E+QHlE4KmoOqp+1zcMg5B
SPlvzRAyNaKz4uzw/O5C1a7LaHvrBKQkDJdZXRTf1DUb+jnTYtbE+2Molpf3K4+RohJAm+ZjJ5Qi
pFlxTmzb4z7xwDd9GZWC7cDNw0meBz8Mh/lStxJZWtYCBFw4qHLhUXKjpUQa41hyIzsFFuzYxSzH
VUQp3rGk8se3F6ylCWg7Fe3Zy33Nc7Vf5f6+rdjtbUZdqicukTuaUA8k3YWwTw4V6i5InB6D6aoq
9j2LfmzmTGS9sWoI0j1OUsdq8fbH8/5PZ6IEFGbzljYkaIy94Rshc3CXyx0A4rY4sXWCkEzuuq2/
SCzj8NKR9N3g77/+0zYk6Y/NDnH8dVQtvgTu4aPp5oXZuxGzkQTEoneExHQuaWzc8g768M8RLqdl
65RIfqLwebhtBv/VVSmFmX9uPTPu/w50ug6I8G6z36/FC5GGt07gxgN3vYAC/mbd+xrOz65eifiy
NXIfAqBEEeaITPRKOy53JiRN6TnF8iEH2otGWsrENt3mxICln9Qa+rQEGuBo4NEgRgPHB6nxfZrl
2Uskaw1z5j8CM+GJtx4/4veovPbFkXX4LtsiKU3ZuLDxXA+JwA451Bvo33l8YCFWddQzqkEHPt2t
D0eQL1aMjtK8/C/dAi+tyQgWdBlTgkcFU3Cx8mMnlacoRlNPmY90Z1ZmiV3IqN/ivBl6TNDQwIfF
2OwmtxNT15XuY9gWhR3zBB+1VFLO60Z4Dvq5r7dRMpHxPy1JXPrEzcXVb7wuMh5/M0tWltUea1gl
Sypfp0ItPpBW1euQKV7XBG8Ruu1jr9ToGYdzT52XZH0sVCVI2HBqJPRhgXnTOCoeFkhhWqLsi30K
mOaxBbFvt+tUbgbRL41rY9g9hh5zIAks8/a3Cn6YxjW30ZI/SV8Wr/1uHNt9XXJziJG/LPJWU+g/
xkURlCPWQ9p8uQLhy5JNcCG1fjL3QA7zfybhlw7HWkumxtLmOzUuyGmwIUKLhZG0M6BIqgwe8d0U
ZRL4LoaoiyjHfozRoFvk+R9N3/X6Xi5KbcvWNkOQ75ERXjCtMZq2zJ9SpvMQJFBG/iuKTV6CuSwr
Wsk+WiP4F1EunDyxeKEiDhU9KAOgijqUTTPYbQEosJVvzOb4VE7Jc8d5IK41kmfZNx51xzqudswL
sRXKrWfY9nHkBbAWPKHkVK4H7Yq3vzF+zGo/kgKFg9Sj+wV4qDkuH2fu7tsUphIIXCsahgHYcusQ
OvbmDuZC72mFTXtYl+jQdzWBGWfSUE/gHsd9z/0nPv2ghiL6BX2P0AcBIK/GmBbctZEcm6/h2C59
IGFfk1X9p9D9n4e1b6Z/qEO4K6HTn5P+PlWuJs7cG/h3iPFHJVtproQstcFb+RjYnGW6NG49W493
deJtkJXpVlE4qZ6x2XUGxQ+TmycdmpiGgWdxLhvvvn5j8A7ZF1BED+jtPNphyGliJYhZg+uNdZWX
tF4zb0gWnCcgE9yB7+peqynwWko1nCniFUq6knA09cKmifqTMxQ63nmeGKLP/jTtLtonrIKtB8pt
ssEOWWycnQxEZFwuJrVpSnaXQl7cY0NSWnzKCIYrw+hTq1+qJ7VZsewnihrIxjQSau8CFS8UOyQ9
QzmteDO2Xro4uVacpq1WZ7Ryqts0PDPT8kCtF1q4IYhYzyKcLyOzGztng8dZaUmb9JuiEbKCwmk7
nLQAfWhVpdvdkZirWHkatyukz15XdU3tkZNFQb3LwZvu3qjEfWSpxCeZ4CNUZzSzyz+LB5dETio4
mE6JEbBxmlJ8sle4rPxh8X4XENAFvUcsPH2EEYZ3vKBGzxXH7JEA1dXmOPeQgHXg5Okk3rsNVOzm
SYrDzWECzw/dHnkTmequDGVH4dPbNitAMOgDx00rkjZ8trxDR1UKVk6FSEauY+cK/hCrBEui/WHz
aIgg5F+jM6pv8L28FPQwk6GsuuLKVPkLfxpw4njaWdHfvhtHVDJqywZOyAL/ZWZYW2uWjkT0ZHQ8
uJVsxCXrPlGK4v1LWpiIq1x6Qrm65gQTk49kW4ZxWy0qrUqnFpTNZlnAN6ISBSUhlzEeeaJaMm/9
J6Sk+PPvAB+k0aFSXEmzeP7x8ZN4SF4oXTGs5SXv8Y9jYczDHTMROY5vWsVNcrOJb7pGTpLY1q1d
mEWaf7r4tITHFjBIwdRdyILBY1OXalYJU4WNvnpRVXXCmcErq+YhWNg20JrwxizHc29APGGioUjA
wKwu93yKrGA/K9DhwzwmbQJOldn9GzhTTuDh2WHvzlPfAU8EI8VOox7qVKPZ89C2xVStE43HkIjW
0AbFj4tg9JkYfCn9uOq1BOtHghuhMonw9kzMlQusqJ2MgceCLEc6Pethu8TWq6nqW2OmpmQlByC7
LPhOZMUi53wOM5tkKJuSGbkndDbLyDiUP0y4SOlNwwkOoTPaKhGmbzHa+NB2eBdHNj9W/XnMOfcY
+Q6+MM7LSzZQ5rVlR0ZowHuloWs29MXKb0H6lsZtjWbUjBLUUrDlLHkgIMAsvPFbeMBtm9DDnB/S
e2NMbaaVPoN6StvV+aG5/ZDV52zwMBVbw0ExilZ2VkeL5z35IcgBjCX1mq9Rfxc6LuWFCIlh8nGb
lZoZbwcRsP5j+VXbe1SvjfwUof38Mf2MejTNEizReo7zxhhjmjQZKOVM1RRAy+RftY8HxqP7Ethd
h0QzkUTHrmZbIZCdQnxW3nzBYsTUF42Z6aeG0DMRtuO/lmmGRw1nt08HBiKhfgBRKXLlNONVpTqt
uUSElNY8gWMVyJ/ejWt4MR9HwvSVyhJ5OL5ugGoUDXtjfb6MEtknbsVgCx/gMtnQgODOQE7KJ/rA
0LEm4TOufrOVcxxyihdnkh4O8B8bybfgBr45Ncvylb3dtqH9jXHGibaqtxgsf3150M9v7kZvB/9i
Xwn1XIfPOZYs0XIZFAf15bUNrdzFbmNnrrYkQHkOV7HAMM4iz8CkJ3spnQjGzbT3mwUIMZIJ163d
9vhCwf8FCJT0BHQOgPD8FHsGOnkAhxAMXs8OitgQOYRXmv3+EYXAGnM425xm0hqOzdDvcFax2ewQ
Nksw+7e9AtvS/D8Y+UvyVeormn/u1EjN/AzhBHMS0XWqeYmWLWWgCPZ/cMGER3h2oqTavoqD8Dzq
w+vjanrrfcfGHa2SuHQ32+G8s+VQGyvjR8WQ3O9JLRDSt+CTGZ+/MS7WZrEFL6ucoFnuEzft6HTh
yQLSClwtEocFUJeT3+y7ZXLSe3SLXz1xMh5hnk5ST93DByiQYI2FH2VV4eROpqmanJgWi+BIrkwq
V2AsDXykmDkm4MUc6qr5Vg31xodrme2/SC0WcrBk9AZNywFyl5cMyL+sx6Mnzc7qbzCuZJAJo22A
yG3LU6dq4rKsj94MorzsIZRqIkMm9hB7UR81YojMUxGpb/5Eaju7ZpmEApqzW1+v+Wt0NMKRftha
3gNpMRK/SOPTZcRk9djkTCnMK5a0sQtsRaVc26VtPsIHad+A0pJNwsbHtwu6m1+/WGu0Z/fgTArr
bLYZYDC9Uhw6xHhA99mS+dREZljBT/RdIcYnszenr7IFysY/7tZVmpmg4j2wrCO5JCgAFsJ3/2xS
yT+jfmHsavo9n98vK62WWvIcKLAP3PjElOb16dnw1ZjPpIzX9Ruq4Z/kiWMCH15yoV/TahmyFOYC
JoOSipXBS8dn6jQc7vBCkQmcHHPDZgH+0Y2ysFXAxQ7plt1XJUocTDK5QW/xkmYv+lhlHavhppee
AdmfdvYfakFaNXfKkr4EuVlGw3r2CLy6ocTpzCeep28fZbGusdtMy11EQmD1unHger8hH57a2vuz
hsGAhL45+lVHV53XrYKkJXWenScnH6X9+zgTD/Iz/gLwgq1LNw3pZs9EElnEg3BDgaXx6g+pY84A
X1LPWMARMkk/MDWe13+YYir5GZfMwIj+Ep6yUZQH6g/YRvTZrTUx5FpFhjfj16vMT4QDsPf661LR
p6P8TxG3KvyGP7HVJwmpYH5RnE3OksQ7S4G5NzATp0tYhD5BRjcKC3y6jd/6txtCJEDBFHngDDS1
MSh1AktosteKSpWeKbsYlVS+xfTkeqzm3KyHagHfHLNVtI71NMoDr26nOFmGRNB3vFh5P8oKe1cu
ohxiIubwOYIO0Bt+3HAraiUFfcK4DLzzYbTNZzmsVwiZuutrzDkIyhypvfvZF7x2shQHvRA9cgZH
vs9oeWhiVBBguB2vndGCyjicOx5XWbag460asKRax5aSNoxKwEl01lAlvlvFD0reSD2RIhnujOyP
VP4vRDC9f6WzC3s9lUItqRgYW6N/1r9Qjku7dFYq4ALq0a/6sYPQIHJHGDX0xnuhSN+gb7zl1kq2
TD129HX0GcHIrHpXpp6zx2faL4pzcD63ygXOu5J+NGllvQArQD4S9/3DQGDXtP5Ksjv+iPsmOc7n
ywIanIKRDFzy38hlWmnaFE9cXnkfRWH1UUr8SHTLEkQwzQQkGuvutDV2XWIDWpY/OfJ0zAz/EY70
3u7vOfI8Woy1YKpMUfgl64dzvbkXTOGlWoATBwaHNfADkCOzyIpnyALZk/ZFZ3ByNys2pQwwnHIm
I9EcmY6Zs8XElSWgJkN33aobDZEnNmAwNfPVD54/B7b6vI0oS6WFJEY9IaCy7r6Sq3V0yyC77kiy
l03w3Eyv5zLZ6GXTZu5iQpRxTqO1SMAAQJb/OyD50CotklI/39EqiTMj3rpbGTBMeUO7AjgXnBkN
g1d5s7E5gefmkdP1zIW4FDpPnYNF3yIV6NCJVJoOtkXWDVihUGXUpgpazlkhci2x2bWhog5bY5dl
koKl1foszy2RzBwIqoZvAnEoKpmxXa4NyVBKvPmpJHjmW7pVgfLP4jkswbPgJ8T+TJhasv5sVWjv
+p9y1Mq4fP3t6EEqEs/GhRBFAS6dcqU2uoawvHTkogkvhsCi/wGzxoL7V3rP/SUw2LC2DW7h1pWS
cAKvsPUbCgf0KpZ4QBrHo1cYFTaRzbqPW9YjiFotpDM20rxJbpBMzP5XQWHiQQiAc5ePJ1U/KwHH
DnXhMLAAqzBD9FVV4GpBp0bI9HZdHA/IsV+FOKVupwdWRYiPU0OMslRweIil5Hr2NmvncP5rjl6d
ct2rfLmysppq5sDVN1Yl9LZvzAosyHeZ/7CE4x0gmEF7Gzqf5l9kibTzWM2CcSaTXkwRepZijMD2
azadtvfrAlUkB1hVSGC8ZHI1nqMmSSwed4VJ/h7Y8uaw5kSRnBCTGG2rQbvi3BVo2qGSxN9nctgQ
HtqlsUVyDkjiQTPFeKB834Rx18WCkv7Yvu+xIAGaW+roUdsW+2CWyEvgUV4sRAr8q7sA9qmBTYXP
3haDHWv1U7F1QsveTV+aUITW6dgNLeM06LtWVpiCWOt3w3Epi8jJL8ScDfcNhzKjymbRJW4v0SOV
udt9FFDeCAAI9jJLcf9l20atdMlfz09Mfj+z+sqlpku2snwe/sK0v9t7iKGzHgIp4/tBn5Cxny8f
4hHfvToY/a+oURhBzOokJ8z8N4bLmJtrdNY6fZtvoHc7zq7Q+iOfadMvPm01L0JU6ZMw8NY7pQXU
TGgEFEeAisDQtCRXfEMfjkDiC1wOpw9sOJfo+O6lFMk79mwe/DolsenkUHARPlDNLMKO4WXxYnrb
wqGa27dLSftD00n9MsLRPBjuQd1Qgn9WJTvG5ymEGSSGtyFurHzRyO5xNL6Ds1hhc2tRbrd9oA0J
ZmVDK2xu5VrdM5vU7B6k9XNWCOVJhLqd4NSbObgHNebMG8zvio5zP4UeoPDTlzR3DzAeQuShapJU
r4EQ+M2t83AgufWuuWPGQ/c93v015GVviTe03D954vhsUgoVsL3oj04rIPDx+UCTZSiuZEcL7mwo
fmc9dppyw/b4TPS49aUif7mKnX45UzB71MlEx7rqsUT1S79d8gb4uMIBGEcC1rD2VX6JEdndZ3uR
efdKdsU+c50vggr1GmaneoiJmE0QWiwbpWt/Lb+P1Q6RBpZRwHhotUW3CEmNCOWDOWz/sWia4vxJ
9gyA3yNv1ObYoNRYMzCDFo+qUWZnaoW/CZ7lzrPgU9k7CprHs1yl3iywheEJNnJ/mZR50kmyW6Lo
TcPAi1sxfOq0cCainf4LrP2mJs+1qcFfdvJN8NIoL7n4EQgOEH0MEyknJSKbQPXFIzBK4SIgeyl2
J2bFIS+yXAl7hhRxCaEvVIEqew660qwiLAT7k0zOPd50E7o13yEJ288rY1LrdkU3Z9BGSJ/rvfx/
Hi9VIPgCbBn19xjvxbpuv2VKSJU4nK0hVRfw3tE9YaX7IGlp8iddwfhkm8bh3ZGyeU7oH1Nrk4mn
GVAsccC8e4jssn7H9BeLHTAcnTmU66oVTCJtN/DexTqC+wCteT0CIhc56VZPJXvDah/woWT4ETYL
8Te1RD5LEZhYkwHm53RgTFgRHwRSJorXAD7xJqeerPNjOyfIJLwj7hFrcBjc3T1jiCtVhETtbbVw
aFvezgFLV6t8aNUVCJgQfV8Xk2QPgfoZT8gpZSmyzuiarmNPrtSsr/ZhMZBXaNJYNz34VytmXktK
xHHa/D76WC8N5Twjl5MVg5LFTgj+4AUSDSVw1FViaFsMQhUtqND95iaH+n5+D3BLNvqUHJf92UlQ
EB68h/92y4/RiubQwO6buVd1/egAmXYCDwlUDBULJf5bTgBmEtFh5VxT2jTRXlzo7U7qZbYeRVGo
8UQLVqrnaJoyAMpRIOe4za81tK0AOb1qQAm5sFOfweIIUeKodXReTtcjBLsW7eZlRA0L0R96xdM7
XLrzaheabUWwO7TqEvv0DKit70d2228XWOjpRBD3mYO8OI0xqFuFkEQQhAMcaY9YKLBUegAqHY+H
8qcd+tZfoedolsvm9ttk3HPWiSHLulaD0NZiGUhOK4DsrKJvyJi9jAcZ0F9Kwf+8wTHT/f1qs9nF
e2YfsHm4zuDSGS/ivTMSCd+G4kx+CvpD/R83ZQJm8PSmNHbwUAoG+cuQUiYxwQ3qhF0MQMgB/Jdu
God8vJNA3VrS5TVsCRRgOMgXBz+Boa8/scfTG0eUyNJ8MZT7P+gM9SV7YkqPIAt0aV6Ztdefk2Ng
4LD/9SmDJucemWHpbw7GUxq3z32xu0QSt3yojiw7d+flxmt+VFlRH+gbVmOVhQ49DOwW1NSUKSAD
mztFX6c3RlgOyIUDczzTkXVSsNjL5k1nFadWhBbyuKnqkN1dfgFLXc/NU994ybffO2fDUIgBaLeT
NrzJTgAPVwlN0oY65wtXw0DNGAgpPl2IJh8WWN10EkNiDnJD0Y5lMZvvurbElyP4SJjAyGuYds/a
9XCTgd6w6qkmeOj6K1288Fc5R1falBDR3rYEeP5+yuTOGxZvdYDo9TiSYl8IgfqsS4GQ28Gn8nDp
qIVc4N4HMeo3D9o9GsYxyYtNBtXqYsT6jOXpUG9CE3KFC/0+rwY/RYlZ6fCe9Gjch36enYq/3Iot
AaqBsjXlIPJb9kOhiahXLF2ySSOznQb5z6NjvEtiMiQ9M+3YxCL7XtB+T20PWI0M6RrZxDVsVjMc
SGYOmkX+IaUvcgWrsD5i8kXGxHMfMAsqTQ6gknd3F/bhF7sXaMXGJQ/Su9+DsZJIEEISDXZH7375
DtwMtYKjtWT72rscE+C4gt9Zm0HqM26QTIWWh+1pk0xCaSP0PIEV8LcMLwe+bDdoQZfDfPRuFxC1
GqGsIYtRmMDIZ24URXCkHlHPI3W0V5sqFdcf4gtIZYeYCDrDNxc/QUQl8OQoOArv0Ehm6/nFYcMv
KFB1KcoanGEJUrsxwurn4lmjENRxEXMa5vzh19xJNVSfeh12LiGQCEfzNOqzGwFWWq3YpM4iDn66
q1SM5DXyGRdPnw/REUCrbn8z1YE0ojhEOLNzSskLl0bHJF6AJWT3TX2GEoOLhoYMQQCRlDKf8vWQ
qY73UXyAsjRzb5QzLZTSm39RF4TT77GqSF2PqIVbXZ365phaeMVfVdvZqRPbHo7tx2AaDRsabAw8
Wn2kc0Sv54y3cdQyZGBFkYFB5Xcak79WyVcYAOEQeVhR89C/a0XZBcte0hbbRAwQhqRVtzHI/t2E
dUKPNLpR16XhLu2fpgT6lvNJ0Oqai2nh6qP8f0SEjxupspiYolFRUic3tbn78xbGrzVnuAMcUmnT
eFsuxuk7ZJlnZm9aO6dQBv+cEHt9vRAk1xy/5eGdxcDdGdX6wXVN5p8lSv98SsieEi+223bjPc8S
RNm9LCabW9WhHJ2tIdwR5bh5Uh+zatyW1qsDUtGCh1QhCXdhY2XwupdpD0UN8ja17KkedTQAnDoX
EE0CgwARHjIYy3GD4GKSZuvDF011O0WYC4DNuZVov8gfwABrmAiARtVpVp8XvbuKfG4/8PTx5TkJ
Xce/lGySQWLGKEwnJd4Tuzi3dQ6WcZbJT+QQLWY3RAghoJwiBio4abbNv9M0IKaXabGIe9+65eL0
LTBJ7ZdWusyv3VPSXwesf8crvGnLXVk36Qq80qIsIaqdC+yNDyg6t1W23ALXCjNTGkACKWf59Kdp
GRsACU/L5WMKXLspMg3IjJtUeFMU6NonJ4PepxdBE5C0OIU23TZdrw7KCiro/TaVNcK2dxgp8/73
J+T7v7R9CfjfZbduZDddJXevkbhomaE+sf39uxXfr+fbxosNUYRBgc4rJD/EQWH81LQ7Qhj59QYO
bgsZ1SMkaguxZYmr2RP16/R1P1hEx3MguPByl8UNxYrBf0Q6TZFFo0h6SZFsXGhP5yZHcp3VBQ0Q
/5hGzF5Pg08Nqv3f10XGWwtvJyaYy1/hMDXgY0ITCMtx/44ficAnPskQ9M9msQjerJ8L2rFwUMES
gcom2TEovePJ9rBXpM+0xqmcq18OmwSsPt+QQlImYExABV0lV1U1KUUNd+e7V1L1i1P3FFMwqZwe
rD6JFLNnikeDR7/QY4LSZAJi/vJzl0WFxvGEV3A3Sxe+yCskzpjnaAl1bi8uowfMZ3/1M0el2Q3z
EHGC2nu92aUlup3MzTx+rFkmx/JZVYeN2r35K0JtfUZRodFs+8VD/Ac02Do+dSADJ+MJTaRXIoWa
uWFLM8sbX6ykzi7UjxT420POZFxxbSW0DalJnIRCpYkVRAM43daS5QR7BR8tKjaWyKajjZ3pcZyn
mTwWhLs+/vuLA/Yz+Br7TTvYNnkIOqpqxVf/r0Pso7gmrqQ6qqLgUXYrDNrbA1+3DnJZeU0iHptQ
64nV09lWnmPKhbJhFOnTHRuurrQdOA05WafzQesQx+ekwZN10j/ACZQOv5ctfbflU/R4Eg9rAhDk
K49zdfQ8AxMsMaWecgNsPHSHx5jilR2uYlXazyxsNaIaByKSnBTiwbLEpZPIUo7tAyBbc+Nk+eoI
My8SDwdDILGwGSvNPF6gF7eCYEwf7ntoGbOVFsvXWrOxS2rLMaScAdRcT8kzH/HrVCH053s+CTus
IxfqEr811cBKhY1tqbdSb8g6yHzaeMIye8shm0ihtRmWVY7qh6YUMTFaK/Elgv/6KPgQpXXgbqyV
VEePB1W2V1KOYozVb1Gi16c9SaGW3uJLqH4WU4aRhHlG4Dz4jsPuvBSsbg+nFwpbcW2n9dvayR+p
EnFqHETP+2szNVeFYicyv2JqrAAecvafdZD/xMLdI+6VvlRQdtqpwLpn8tR9zCXtd0yBFSDZU5BG
v6PhvavAauLg7W++fOYNVFlEZMjtXYMeCTmhXnhxZqYigs4eIpDGcu52UG9Pf1+1iHDteMRWHy/W
52c0byJ0IfyQU/XH+XrTlzN0d9/DqAS4BeSyZADQ47zdDhX3wKH9plfuLhZSjOYMJeJuM/xr7qg0
MDxCTm6164W+ecraaoM6skTdziqlIl+dpmQ9y8tsIAp5qHPlEhQoaEbpsmECDwP9xgJe+fFBaxNv
CQcSr9+4PNfMaitXojPcjsn2XE/P+Bf7ev0TsDV7ZLd4S127MY7xJw+Rgxi0eQn1PTzWKE40xvvP
vZsoHrea200c9qSaEGVAAoHbIxWMKPtqm/wlspd/B4o2Oif+j1dwF3d4izqJJhQAmzfxh/0lYu5h
Q8uQsWxoPxSfrq3PjrYv8NOLql09Sxuz/uX4dl660QZRDI66r9sZq2Q6Gk7XYaW44Qde+hMNYk2K
qCQTIg20o/yWKQ83Xl/6kZ7BpGAVB2U2BUsiSAhxdOwsKzsciF+utXCfP51N3o/ffTUDypwtrzUd
sJHBuKKJiWSdgmzxGWvdDBpA42geezqjgK1FQHFM2Ah/jRreqMQI3nMqnkkG91GSUVGoMDWL8e3x
HoKp76SIfmAxUNAd7gHSkGaQGi8MkhaWZOeCbAojPPtJXcKKOWUpysdQlh7dUnyb2Jod/FztX1g7
ewDZVDKkt120ji1EQ/eXSybG6v8YM/trdE0aK984RMn59gHNt97OnWaW+KXr/ZS/iQdTdY80ArMr
0sk0GbmGB1dnbuyXISdK5LGP6f2nrKbj+mKZk3QVab3HgF3fXhwqwvjDQ7Am8sr/zI7j1NQUX5j5
1A1vVoBJZO4HFjCbnsj00OgwGpKeygBOQytcin6/MI7B9Fcm5z2uOpZ4AKquzRr3dJtp4Kfyk0IJ
hlq2utYpqXoRIT9Eq7Xh/a1sNUbiCiBTu2nm+K7XM9kbpJuv4+QlwDsBO4si8K3dx0tNHrrw73YO
zxfgFEwi+gCW3h0eZaq9vvDSt3v7Jk3u0lgnEkfq828JKFDexzkuc8h8OEgy9Gbc9etHIbMEt4+t
KCjzYXWmXSMI/NvMSg3GVPrn/B6w+CLVgiHNMQKcZF792Il4cYElvpFAKa7WhzyHtm8/QYk4rfAO
Gb+Kj7vgNtbI3tZ8X0WiQZUVL+XeooBrW25RswQZT1QdVcxWHDgPGT2keroIZsO6i60qFMIaKOpe
FmYx1yoCD27cQ/H1xr8yUzZeGD4tkfcEVgn2otmSP0NqYuo+seE7p5kShazik14vk4CFJlJGEmHj
eHakS6PoUCAoTZCiaHGQkaaM1mAJ5c1hZmPicJNWUCNPh4SS6ZJb/35y9swMrdUkbTHUbqNUQEHV
1rCijnqH8Iw0m4gvrJ8MSqBZP4964ofcdsAzQra88OdG2r8Uteh7aNfmAuC9yJJTa9IIpheRcPw8
+qE+ZBGFN5OXvY+nT9VdQnYcmUgUPEyoCu4zrprVircin3oGNSTma99VVBieRva4uyp8QAFesdEL
lwV/kjf6mDa/dYHrxjaeSJsYNk/7JvosvXLlKPpHobIXviPEF/SlGqwkMdIlKn3wBwwtXlZpj5am
kpe7oXkyokqdIXCqUQdqgb/5dPAgEfozSJ+MfX4WC4ltI2geR6CtZ6nnpHq9qSeQTH6xwisd77/M
Y9mKOe7OJXXNzNMlctx5+diO0r4VsU92ROyrffM7PrZguitNOunci8NGIQcH1FxB7xLLYwM/pU88
ezxyK5i40BE93JkaNR6gmf+QTEq+nhzJeen5fm8ieluAPUaWDUopUKoj7Cb+GmItYq00VV9x9dEP
uKRXWK8n4iX3bbGaxB7pqLiURsIPoA+LcR1zqNPMs1AJoL3TLcEvYHWuaKfYbRylWbxUbPK28dKx
hnG49BOxF729Lo7HcEOyD2EMu4sq8m3lNxAx+tTF4BcbeTcGmeWwgHXWAI7bkTrhdKejmo3vSezd
afWXawKRr0HbHRuGkCg8mR+KAis3waCyqs2oS2KcjTbpnI6QTQgWMXHxyknSGRCz+BlPrvF/x/yN
AeHOpksUb7QYhcmIFSZXftSRv/anWZfiyai4xNcS6reIp/Um7YRI5PFLpY+bfZ2x5LNnh7XVAmia
MypJbo8uvkZBgJ8Xc+PbHQ1xgVauu0ToC1EIG8CgoRn1X8sHHNUfalv5ScdklDswyBF1vk75hW3V
rUHBv4Wg70IdvsbVR/I/rPlxPKBkbS71KlpIAnv6aPrRM/Nmz7+isYmBR3Lw0EjxJU8Pr3mdH+Y0
QvGU/l17/m1yDCwmXBnG6Egu/qOpZSq6vFhFeLgCcxMveDczEuG860Ya+OEZ9ChbDK2nBYQD0t9Z
sVxbi6xluGMPznea3L/HzCcOotXLSANj44k1GAiVXNZpXpoKye01xcP6NoaQ5z0VMzhwIwZy+56o
kbPLKc3hBocuVxn1gcMf6XWprKFuc8FmcS2uOWS06By0r88zm4Q7IgOikXDFRTboK6RprDHGL28i
JzPc9iqBFWQprwuz8bR78ks1cXkPB8hM64Xk9t1FiVFJeuIYHfmP5ihgJG5D2CtCNJEjrvC0fbif
tNLw3B8uiLjoeUN28c1cxpIxG702cAo9ASWgXvuAOcftT/s3MOrkx9hlc2pQ5xX34SLuWapXldk8
PiusZrES2CO1r1fZCp8x+xq3BfmHh9XiQAgapFor72lc7Al3L9K+3Q6M9RqtJ7dztlDhuIsp6BM5
UFVgY2owl93GBBjq2/UbJnWNWoz4nLddo7xGzUKxrKdelkcgdWd7Qbyu+G2QTXB7n+Lj4jbnCIU/
qVwSQA/vVsGN31jPGbCPfj0pTkxkNPz3C2NukiCLhqbKnq445mmaWw8dbo2ToR4GPiDytd3IZWmz
lwmmIPbYy5zCVo3beH2Mrjcmoj+lVCWAfrF9QB+5dtI46eS8apZKeJT8tJcqBVey1Jc7xm0YImRb
3bVv+5oCE6011PsKCNA48YJea7p9hMqZ4qep3CYesA6QOp9ZJDiAKrB1ZbxwH6tAsUsg/yLSkTEX
b9L+cdcqgIPDo7QVjmLjtVOPHMzZeKAMPYgcRzJooxVpKSnsnU8R48yL893sprIE4ARn2uEV2uG3
TSHLBWHQQB/QtjjHv+4rkRrXjsYp974k5JIkpqATxZqKTvOGeTUDnDkWbOIXCuVT0vxSro0B5Kjg
di8kI/FW3cC9v6TBYBOXDWE3BljsGK7pyuN2ersLGPpy2eLBqHz7Fmt/2NRxtnZoEp41rQNW+J6W
PSiXch7INbqn563tj1vL69hXEhJOYXmcoJYWp7h9msT80ofsqnesgaMzJ2rjkss4Cldbbd009+zt
iDOleG/zVOoMVf2VdvlXXnfOalJBhbwtx+MGoFb3tab3h5V4QewbP51r/+Nq0KxR3s1rmaupzuIW
rMPQ5+ErdzantoLk0f/9EXBk8bKdRYfwG+gIFxl4g6HM0Y7ybDgk/AH0NUf4r2BGArTXZ47yZhmD
FXJpXTwYSRdO/J1Ejhh8e7oUShTec+yQuqAmzIkAXQHXnCRu5Ep89dbNch2cqmW1gC0DjgkNhcb8
h7te5zU35beQtIY0pa1Nnk0Zyu60ipq9ykoKuHAzK/Vcm+lE+DjIWqEA8Hu8QuXllq/XwblIaWDe
ERyVzbVTJhRUbT+RZtLCqwJOJeLXxcyjBjY/kRu8J9xtP0+JWuqNmDDQlf5i3pgzEGzkH6E+WpVB
MHksMNufd2xa19PTQphUGoTaRBWXW0aCNUjgWKOWTkXqMtFl7EJLMkwsLDcAgORtr6ebdJwN8+OU
to9BKjnrputpHXL/m2s1xdvguMIby7gaQrTb8eFidy9ZCP++Gb7y9mupZTYs0S/O89A+jlYNVWEr
wBxPqFYAyEdzGfB8Ag0INVE6Cv76WHbPfKnpm3n0IKE8nZ/ZlnfmtQ7NDUpK1thiWl7VCuvJfURu
yfHIIo41yCM+Y2FQ16FWCe/yZbJhTybL4j6uuWqcXfPWStIcJh1bXrb2Dfj3p3SK/UoPrjUrSDvI
80FnJACViKR9oQ7Nq0ofCKu0f7ygZFO51XGufy6jQlEGVWJ+4nBKQJjg69kLtPlaZtg3xQD8yOWS
C6L/q92Z4ziF3JgxaauW3dwcxaY2ttiEgHUnkmNfSWhj5/cEbRrafgdHpfO/koTjNHRxn8P8LRx2
jK83Uza+Lvqdb5ZB5Ka9uDiDubxWYgXbJvGTBsSYBc48YWK3Lo15Ua1gfRP3kimsQ5A8yDdIsMNq
K7gqg59eoFOpv7e3iibzkINyO5S9PaPzzrkRR26DIJ61U2fxtiVeKIC1fMQE2u/cMrfMHSolhOg2
7gidfCeY3hjWlPo/S2CPW3t50Tu+Z57/ToyQ8nfl3gPaMoS/UEJD5eZYDSfrROJdQI0aBHOa4xhD
k1E4RpjAosDASUu6xvm9s/t6O4K1slPhKunHs3BCBovSDVOWm041ODbY6JSQ+gtiW8iJCYQNEhOl
8CviG77K1UbtvvL0IHIcxqoMEDfAxLozjJLZaT1mcF5YhMpioTkB96/yll4uIGYEeFwKyUmGK4fe
WDDa/ejdhxi6Pl59Z45MKP7DMkoagzlPrPl6rNpc5Y9T80857uxtUFbypK8qE6MuGXna2DiSRcL1
Wde8U2o8mRLURNP+FAw0cZfVndjtOZPnBkqvpJNovGJN3/0DmlOJBV0mvz77lKv4DcYMOxHkDVK9
ewdLwujWgifVOm69armkqIThdz16ZEzJLGqRgRMiJMl9ALOj2WXs70yx+S6MesTZs358/QrN2D6B
d3r0pJu1QBAGR6+MPXCuG7bAMwUtTiLviZsqPoM4rUh1/6kIbbXrvpCLFhWQm1M9AZUgogvfAHVa
pfYaVgz1E+3HfV6w9x8DuLw4YLi5F5vYeB7Qob1HZuRjKXuEr995aMZRetYWHh8wLERs4pbwFs7a
sFPwaTSRB6vZbvoDNFYhFKayyUCvwO64WfKze5bNY1kiwWk0nm2kbMX3s/zMuY9JLtKyTVBFsi5r
12668zqgUqlNp0aJr2ppyER5Vqs99xKaGPjDEquh2AsgFpXYxz5Jj3s+bm8za+c6c92ib6H/K3xM
fZkJ8UmrZR+g6+N7Dh4M08NH3l1H3m3Pvr71lgLMXgJvK3zsexD2qrI+ufdZbgbucwha7BToNLnK
Wxap5KpE6gYpmN1/gPwrY5l9G6OGcq8Wkdx2EVChVU4hfFh8udbWGYgZAfHo2ROTGm3poFxqUl2+
U58DPHi0VBtZiAw/WkSBqrVVCbSosw6mmxI13IkmOGudzpzmKo/7qQXsHLL4nyRFtNKzVj2TWAdO
1NWtDCJaQHPJIUEt2zFmiYK9WJutl9Oc6PTla6+6GW7M1cDtvjDK/voqsAoSr0AXFgYMDMH1dSnF
GFD2QVBEZ4hxzk52RAINzxvBXXjI561CPV8faYvcgSki9ixtNCclxb7eDMmJ08Gn3m/Ilmw3aBM3
C9X9qSpQv6iJ5i/SpW95PAhYQcJAHWtvxix+LvfjOYMgdAld4uZBVYHZsH9M9/ISpv7UA6MxTcKC
ZqcICb3ATYmrNK9KV+FijP1JRTSOAV0P31yNOFX1+GKZuDEojQfxewv555js7z0GUPsBhecWiczP
IvsjoPR+qo4m9lFlkX7DpFrmYgMf5vh7wBhHLHtqOxtEtY98Kvh4XpUru0OU1kDwsSMqyKKJnkLI
0rBaeTOY5iZRzMz6bLz15O8qXyumbDsggFpBX/hpNws27iP0CmE31VrnYZ1ZdklZDu5ayAJda2+c
4sQpwmrU/sYRq7E0WBbt7ayvX/pEEiycKkNg6JHFWd1K3zwLwXRw7krneZmow2twUFFaNNMhtgRC
yPGLmIQBlhr7IhGLcsAaUYm81MrGEEsMXwb1Y65Ymxrhe+tKjH6SjY7DGXx/fFltdD1RzN7RRFSj
K0OrCab7V4keBLmRfRnPdRHewxx77d9cPw0zBOJNxcv7BM2zSk9+FueO11B+UVKdCDx609ImjxJf
PTSYOIujWuuuMiqheTRsMJoOhsebI9DhbqOV6jXkNA9DyT0+0PH6p1cRQZSHphzTD56/6edCzvjy
97oJzyJRj7rhgZTW3/5OzW4Ul/wjYTl2HqqTBrt5qcMOZ/C6fJ4ojZVYKldr81Pc6oeOaw7v80cs
xh6Ny1jtawOYaTRNgO5pZx7fvaA4wvJz9p0/pOcUuDe2TSiAKh0xyRxE9eN5RyJT6/tuLsQRLfiI
BJQJvkgRmEUpZSh33XFp8wEYXp995N5k10X5grPhQtgifxfq6Z+gAMYPYnPPIYiPuRVaLMGqprRG
HjQrfbzMn03QiQ55hTDx0qHJ0UMSh8ERzepMWmLWOGNrypvg/9mYWXGU5ATNU32wM7+IUXwtHI5T
eFa73AKF7q0KiDvEoLpaLfRLqCEs05CNJDwglTgI4V79YMlbCwd3losNsZX5yjsJI7anXSBwGYoH
tS5xHK6X3bJp+X7PWDZvy7lcGae7/20ydlJs+Nm7iwhpjCPeHb1PVFP8gy2/TlXlEkTcKjS035hT
2xwWr6hCQvigt73rZqR16POpFP1CP8ILtycEcmfcLwHhnE4zbBz01kQnAW1SeF5OLzzHOyxn/eNo
r3VqxdQgscgH6aybKVwaujSQkUIXL+c6xnBer+AkYknXHFk+0CK+fzdes73K7D2Fge6/icjLJOjt
RJeFyyDH6w6WG47a8rn1+eSA9PQJn6MsUs8Z5mFnljYyietn43zTO/sGq5jSGvqCYIbEwYXS/Q4C
DXqK5/99w9L31Eevgfl/GX6YHatTyusM/WKmRvRulA4gdQjkPHmqsDCHsts80RFVRmmj2Po+/7Ah
3cy7btaNVK+F2hfx8yI2A2uHvUMBfpjBwcjsZQjkym3MiRTPYGAwsE5/KbcL2E91L2BxSIv1/iJq
jvE+KG0/kVbLtwVBexnsDy02qk+5gYNUindp5tWTfCQ5yM8bdNdf4jm2Rz+NCS8cpQkJbDHBs3Pi
FRE77vnmRSCgz8DYKWJxU13r/q22F8+kdlRvWjODHMgfE+EKO0cMzI4uj1lFroa+VgxAdMajoPN7
3HbuA8jyrxAbCPoZJ2tTHjTEueoXeutW0Iiexxz0DsAFoGOUSUCr2s9rgyJ8Doh3UYNt4a3ZC216
Uk8DzdfPTLx7Fukdt3odlD7sc1dIZFwigw+SwaAH38A4MDF5ZJ8t3p2yrnNf4sqPi5TJlQnX1Mjy
3QLYJoQ5IAGrXuGSe+cLycLrZKvoVoHcka0yu6uqQMwrom0iFvdY3s726aGu2uNf0pQVCRfQ9DP6
m/XYEkWiVHkoksGNgl83OTWBkkr3dlnDCQzfw21QXXVzbe0SGfWH/YyzvvQ0uAFWOc3CYDYhOlTG
A0rdbjBHI6V9fVqV1JJdAe+Xs00zwfb8p/Z4sVCcJ5m5izHBUL1JauiZZjhuxb2qXiGiqIpziqr/
Zfa9mbm3A/LU2NuQ2bSfZT8V9BPFdwg5Oq89Zge0sfNM5mA9mw5YpGrVhgttMke16qpB6e1t7jGC
ac0WzIaPmZsOHEiISFE6lriwbiouHreDlaoOh+qC51m6VBu62eiMlIJilClZv2vyYnZ8mTTKxnq5
oD9yIAb0Y6Emnkm4ZofxEXNR6ByyHp/WYDgS2QG+kHyTPoPg8vpPl4KjnW5WiliZYOl7bIzUtG/y
05IFE9D02jIFPVXBzW6WwTomsvkoTyDRTCa0N8CPqj5ktIoeoJoFvl+ac1TX2a6dgg+fnJ3zczH4
l7gBMYdXBEXzPjzilaHUE2TtU1P6i5LLHzwS8KuMnBlHSTCnZu2+pmuHeta5sGtLjzEp6bhm8Dr8
LBiA8VqDA8LMNbWEw7NRqzF8PSsIYStcHW3DmxCBWfl1UX7YFs9AhmzbIbLlhz1pZxbLvD0uwtTz
4phZNuocskJLOIcJ82lrpXrxiLpIUbg/mXoNrE/iZI4usGIesy7qYPsYaBoU6u2r7kWXg9mTHkku
MrBjlM59I40bpjiffhihsa2fqEtE3ulLY3k4CXR98oMCAzWrQNPhg4q/ac7JtGTfW4EAA0DWKsxx
p7wT4BBoKO8bcfPcQuPtdvqJhJRZom/aV/nVjmrfAQTS28kZdWXqUy5EkgA5nwuXs0jHFcr1kJWa
crWOoivDuBJ0GEDt0mStzT4qKBuT9Qp998yyl+wgVYzl6rBal98rcvyZm9lCLm1UqOveEyd1UXBs
neJViC8/i/WIAq+ZDWiHlVQCdNbEKmFc+IgL5cY04Zu0atrhmm86+yiIOnLCmBPTimlb1/P6CeXC
9xpBs6kAlHv+ErtkFq2Ha/9Kl12HgaC/Lgwt+7Qjc2opnYQugjyCa89ez8Bg1rUiwmHCkPoG4c6O
xHiKc/7am6zy9Xk7tuIpH+Z/BcXG9ivFsc5RTM9PXTa3BNIoxJOTtTfAZnRmV3RD7NgD6WsUfjcZ
5Z/w5pICS1WXo5w1tL00iyTk+aMb64v6AdVHEuqb4bmSit4t/3OwCDOrhMYII1nMdt9XZzX/Tvdu
sVzCfWqNBnAtkSSN+xEnA1J+MEhVQfgJOFJJBmK/EKV+nJMFhUKclDaMGnhVvo0EHEnmtQT3xXSI
u8ra3l6SJWKhNCFqEgiDdaLXEjJTR67TNPvEZJuQprIpkMP9spSiC9h0fVdDhi5h0rsT/I4oLP+q
IuMxog8oBR/ZZ5QPpaBVi0i+p/+4c4I0P8swTRuFHDr39yn8wy8HHHvLedMKEb4FnCB/M8ztovIq
cii7+XP2Y60ewhs9y+/sK0hyNFHNIZ1yWPGJsv/B5vYf2U48ctyOoz4ApmIdv2P4xk0E1+QCBVoS
tn2CIzYLdUq/FPmVS0Ymfv67NCeX7ZKFw0um94LLJdwo3iBvoTFiOZCHK4GaaPsBbGExDw++aIWM
+PTQVPQA3D9R4sb3r2zKceXx2/gYjlPLQ2V0O/Hckk9TY0YevAxMMrNZC64OLtVqcax3O47sUjin
yghk+NnYuEMr9gwERilpXtKXgCACqXmrr8Zksh5/6FpowgNc2EVgVmzevOYxREfxDqnQUPsMdaH7
+BPPkRvQ7OAwXP0VMzrX0/4wpwyliNq8etcUIkR/D989yTrtQEgsFMtwyvItwakgdRmpujHfNn/u
DUTytBNqgQjtu5ZkiBcof8u4ZHxV98ojnLDzKY4fflVm9quD3EpSVXKYsnHJhiJh4kAZkpOfS8WV
H+n5ZALuytG64Iil/jqab7HkyqTYuZ71e5mo1Cscotr3+pW6dKJIWUVzh4VqOrvjpg4jykVV5zAF
0VV5swwMCzFP8O2geguLsGReK/IxFqADirpgIP8UbKtW5qRllbo00MLlQyHykNLDb3ySJJhVV3Rm
yVPAu70dSYFgEpoSIvvyVghWEjFt6SEQgpmrASYrxE1QFnHRtpjtIFiIRGRv406CmP7kEA93MVBU
vUO+xrLaEJ1U/sSGnMhjYHqYtytBzTyuJPmMbU84IUDmoiKQhDXcXKM0eEAUM0GiVitxT7cNOV8w
gAtQ0F6XS/DuWkTWV4xg03VsmaplP0sNojeIS9TB9JdJvGsi4EyXMzMRd+EXB4cNb2u0m+6NeMjm
Ea8ItcC7yZSQBGDLYKBVn/IlDQEvcP/ypbCeZ5VakE2nuvl4it7YrBUszn/7KEgjKNUiY56GWl+r
rh+lNbqwSPJsGlpZDthOvTeLXc0xggBpF9/WfcgBvIxUpPczW3BejhX8X4vcNRcausjuLgbM4T1k
noZxwH0E4pnBMHN3Kg1HWHpmRMEOLsu0qiapdjULcyGN30iQ3Sx4Sxl8x8fSIkw1QfDKJiDMzg9I
Dz4sYv4PuOcRom767P2OaEUS8BRKH/rMwRTSKWiZAYVEULoh+I74cETKRUP2+2nQZj60kxBR6f2G
ZeJ508UE4LukBcwqg6zyaTgx4VL4ki+C78L6g/H0k+ePbzyvh15+o/yAemplkAm0FaEAY3fo6wiB
2AdnQn5n+lVAstewMsdl5L1v+06UGlBY6T47oqBKGeldUQ4amAiQpdyt7L4d48vh8P3FZMwFYq0n
R3C+QeHypiOaaF0Dy569MMX0cjJq2llZpMTpvuipaLsrfvzYOq8Wr28tlIa5OnDcnvNmULc8QagE
sznTuIRPSBvKJJK+gNCotrkW/0VnuoMNcX0teLz2hkLoQnuy7cAlmvo8pqT52nn/uFNOb/PbxOOB
fDlIZBkuZcpNobhgbDmwdh53WfQH27KrNcTQfTN5p8G0rplEuJB6IVKsCTgoOneNtyW/Tbp4gkVf
v4Iflon/ZGprwujqzVOMwvGSzG8fbToaRldQeiWVSUoBwOd67P2AOjAjTYCwpHUGYg6Dw2k/uMQQ
EXgpUKhEPFeVNL4a3jem+ABHwq28YHeLObk+aIwrofeUmc6ScA/y7haQkpGK6JK/zSyB88AmMiRK
VHO6Gdr8TE6wiWz7EA/6RIhKq/Q6ktTlcrb2f5KxnmHK71Ptwb1AiizYg7z2kn9cn5BVRvWcsTaV
Yxy/qVc2YfVA/iIBYBf3nCFtYCSGKelPHsFNg8jVP5wmtxEg75DT7EZdPLNUWnuj8JE6xQMuhz68
ckKZf5tSn7bmiSQfmbcoz0/qVFL9zcFal8/aSypu7cfY0rb/JgAxpyRvpbIOuemppF+Yw0aPr1aV
ZXsQE7C7nFELBBcl1y0EPqdcthuktX9JXXPWJ5rhZEO5KVsqIxuiMXQ9PmaGApxxa0F0+K/Q8XyX
ZJlg52C+tAV6HaHzuFyuDchB9w3pnjQlrp5wTNhy2SNIMeSQRqArRyjB6BmXSx7PInFX6qaKX3/3
vVle1iFuUz1MW2YM49x54dVPZpxtT3tr1IS3s0okUWh1UEySRsxOoZPvF5R+eOH9awAMDXhfmXSy
JE/eNpCeaZKoXEeONk3ekonkHRzVEon8XjB5SHv66JV0JMKJEH2aCQu4Cah/D0f+LPPGchYkdWVU
6PagdJ/WQAlouqIGlke3vd5zdxGMl3wiq7R01+UeZXb94xVAs5qwZusmtZipSQtzWywUA/3jXJP3
PPJIcjUdnGSjCVx3sZL/UXp72elYiQXSC2FRNMEtE5DxzSkM7rnDMY5w16DhBCz0ogdzvGbJAPPS
k00Kma7t0rAOIplhn+iNj7tcylkX4FkIYJSgEnNuL6Dw7PPVjIa2+w3D227dpF4eN5r+IQpklsjD
OrL3nWNO2aV+Sypq97nUtSrU7regO0CfivnA03CfNizZZKYQaId7xmH3nEyv73diprzLuYJNzn+R
fqacxDSPTBe/PdYviWam7m0VJC/LdK/XmRCCWh0osVnuoP5hH1g09dG122kvKiPKPBY94XZSc057
NsX0N6ZGZrIyxOu9nFxsUbux93MMb+msxyXHt+gOTM48+GOqqJq8OaC1haYH1HtW3yDpDbHJSfWB
riN1ETSYarwY5tBH/xMQv6RP6skU7I3f2yasCj5+gGCXTwvQLHHdUX6J0aCmjkbmbhuJpNqwkh2B
wGZ6zF2+wHLW7kC7QIrpy/BNQ2Wfp2S90waaZ7grQAtEyrhSRBYzXQ+hH30Vf2IndrKqTNieWPbH
g0h/KL7hw66ieW09tjrr1d0oBp9nlgwIIUJO9EQPT89ujF4QlaYCM8bwDUuCHwW+LkuT6iUodAqP
frv9m9WW6J/b3FFY/oEZLyTFgWlB8EbzvdmAV/7S2U7SJ7r+a2DCeP0ohjX4HcLDlnPyqoVhwKdg
5XcDF/j5h6jiNzY+h20qhAvZBG80/u0ee6q29G1/mPAF1iCgSlto/L+gm8k5kPc3xWrc2W1q5iGh
O45CxJH4+xl/C3s+h0Ng6A/nU3KxNhGWramSnuB7oZHzOl2A3DMhWzGN4La3OyUb0jWSoDQYmwG+
WFvtPGlzEZH/+x+RucoRgkflHAGYUSMSG8cTVgDIhzjlQtCEb+UlC7WsIAQIBjnNtfIWX2MNeKEk
VbxRayCwBl/l1lPKMZazpgn7niFyrvZPTBDMutvUYSWtbWBajbrb3NovQDFd6Yiqt5Pq8+PVi6Py
c/UBQKFKlqOg1nZ1o1q/wZmiP+LavGWecyemS95p5f89XrH/+JiIxjTTh17ic/9nzFM/aLUAvCLp
iWP8oBmvG3M4v3weqzD8st360QjyQ2tYF0IZLRBrCUdFx5EoxOfQiJXJBNyB/OxcLrxjaNH0Lnnr
/v/DQlA2z3aZxw/mnZANLpKdGFI/Pvc/VZJpLz4JCDia+zisaZignqR8Ld2yjdBF5C8EkBpFgCV3
bg6mvmuFwwsGN7Rk4q7RicyhVu44IagnY7fa/Kiij3C0n1X0akQCFquUdjodU0+7XIp/eO2OsmaG
MuA1c6+++OCB4gBVTlfFQj5uW7l1bSTRl3BCFs7TQVqREP2kdFmM/ZqXVC00s2Nmysj5gWGQOXuy
ACObaY46e9NT+ysCexKJTZ/XXtUrXOS4VJIv8+Eep8qL1g9iT/7gorUMbhpZEnXgxLljBTmtdG4r
x0hL121kv+E1FcOF4ywpZCKiJ1yvwWfWA1p8NVR2m3zFEbgmc4KoH7PeJA9lPLnZggB1NSbeCkw+
4DE4+JLtEb22IQKcRPjmKNqcRyKJ8to/i/ej+OwoET6UwYKTxKHOmaOsLUY/ZHcVGR5eMrUTmcjJ
ga7lKP+QnnXTOGpoYcGEFuxZoFTp2mZ+TFRJaCOvzNpogmcQitPRVbJ70BZjwRs2rGLhzNoP9HRA
6HN1p/HMIBDm349jHZY+IghK6DzhFzFlFptxO2jsvj2ak4ENo3I/NnqRBOVv/C+IHDza0PXr8LGo
SfoAuulSNInTSpMoxWd/E2qsp3f8XQpRph6eq1QTQktlEVK8rzE1qDjlD89lQOEZ9Hdp6a7IPzw5
BifyXKiIGnmHqmfW5KYGr4BXSztgyte6LsYwFOVSH/MzkPxRlefOlZTdxEoCxRf5jg+pgSNbtgkR
LKUSBklaVTqC0Qnk4WK0Kue6oy9RCNSbxncwEHosyCpz6RggCw1MQkBkiavsl1ubCZZ9YeY+FYs3
N1LGtmXy26ZDis5dGVmHeCCLTkYV5B7bEvIHjG1QZsFUNQkhtyzhEws3O34hsEQpUhMClIOyUOls
YWbluJUqa+9LQUUSG7wGwLYDpKTO7Ovgw74wwkdVlRDX1UbenLTr63GipnG2Tpm7oLxkenyytnxi
1uJllZe8cESdw/eN70Zo+SDRS24juXSRX8jaL5/Jo+NSbeeoeq5eDnO2bMN+Zf0DlBaCQzSrF7LF
0Vb6ULOBSDhPyj9/8OHU6sNiuHnnVcXiyeknvPPHNfbmbMD7lDsib06KZckFQfy6/MI49wJcRi9H
h6N6dJ6vqc5Z5sqXXFIH5cdlIeH7RWd6n8hUc401Zt4aAG3je6zbTGHxJXa4pA53eYzhDvc/u0Fp
98d/YbS90qPQiRwWBGXAD941Nhw6ueTgY0cFYlk5kR+1SXZ/gJLc6M7CkuZsbVwf0fcw6VLt/duz
T9ZcewrUIm3my101EJSSbGE5WEjMwoNdDs6OL+0afr74CFiPdqON3b/m/uzGNyWLEN3WMXSyLd4i
unTfPzkFQe3wKBqx20wL8S/NfaAzFFGnakgXc6yCdT/6sCdgekWqRNoUUyiheHuqXvR6uctF1XJG
JUXyWtKUNvtE9QzhQTaUt02azbYT6ivZbq4XthapfQ49ARtnlZr/M6o1WwUlOsf2GQ+M0EHySIPp
bmx1nwZrzV62WQKc549y4hnbwXGxLKUNbsnV6Eflc4ln1PDb1UJXzzlystWbwZA/OYkSRZ7gYwVp
DLhorLkOuMguXBhA5zYdRYVNVulb/iq5qxcdsBDjBccXGf8p7MimBWQU+yX+2xQNRhEwtwjn9xgv
YCgC7h6/HnQ0cqaU73aCoY6tMI2Yd1s2wpIOtLiCzrDN2EjAOJGZYWcSb0YwSYIeJQqURDBZMHm4
lwNZBXxywnbalxXejNnjFJMDud87TuNzo5zAgNFthKlUTYtWsE8xwKTFRLR/P7yNOM6cEqbw0g44
s9Ng6+5utDKXYmhOb4+DeK1izr4ra8UEaU7kJt6EskHqdXb869lmsRPQW3jvtF28l1bc1g6wD8/p
hzHPLUURy57En45QTw5Y/T+k6wmzZ7BYR7u42qDZBsuR4YEhpW48k5J0eeQZ+bPNPMhf4ENiIz15
kzAU/+fdp85fmleKNsDvlDPd4d2X7qqi/WvGiTXC0kextLFVSlSlLke2E9MqmrC0ZNi9ICZn8lCf
3KwNa4wl9pAvIfO/1VCFWJ8thoaFZpweuxBQ3lbzOhL9vLqSNGmud8kgURbvC3qU6fUaF8uVU+u1
njped5jTqqb81qmb4NtPEpIkzIRlPJT45c5BRF9H5ekUkjhN7AyFiolpKnLz4q+1qd4GBW43Bc9O
jgdwiF/eZZKqbSTw/vazeLYjXiwyX5gFM60SEkwAByixqKQo5iJT4/pILdvekEeEjFVTSa1kzRbw
F9dCWCuwVNZ2uRPMfnQXVfdeV+uyRCiLQ02WJFWR2YdCTpGKa9KAxuEMZlVOTynFs2ha33PmmxSj
6UMIpPXfnClvEYe5A9fHpnyiOpkf4GzskbMFVfB/lzuK6Q6NVMoItg95CsUL9015dEVmSTgSQ7xn
dfWhVu/d4QTM/vcY3vE0vHfcBd/bnYrZuj8ICCL1kEGkdB2eYhHRZKLfnoIBWu7uYd8JYs063xpa
BUNSvBhreUjJ4cgD/+eJb9PmvHKifbUeD/B5gh85QVt8P9/na9WVxxv1+KMcbrpeq6kHrTPg/ZD3
5LmGqysKC4QcgZzn8svb6+C5RC34xNd126OhunS3mlRioqAiv0I07nw4BPsCzWs0ZZbngu4r9spK
+FNwhCDXf5eMuyL9SDxfV0UArTRrp7WMdghSle9xfSROfnDe5sbLVvG5TPIVkp6vwdTps1vBzfD0
dax5MYn44cTQA+Gme2jfhoVtXC5TJtSz/o8adJ/1eRZadqvBV1nMkRfjKqK+ISXeE8UqmYJUuVy0
LmvTesuIpA6oyFdIEK13AoEYzv6w7FWFZTZ6AasXLcsyjAAV32Bezdj9B83iNSCuFynF9Kq6hLo6
zUdOp9km9BB9Xe0sg/rhhRKsT28vSbqyqpx1tYrEVw82+QajB7JzI73xmW3HDX9L7DVsJv11p41J
ahF3AJKFFSr1mptFgZqLL7eTL7PR/cQQKkchm6AJu4y/9IBpxibJBLQq2FQ4d4dNV90G9eRhxoq9
wTPbMUxR7D7wjb1LBWwF2INX9/EJfWp0Nx/5RUgeuDGGEfgN8lBBG7sN5f0wlmBJ8QQc5rYg0dAS
AC4d0Exudwi6jv6EAj1NJj9rXMSr5dIxgcSOmZB0SNKNF8VCSWt6tBRe1AfW8S98UAPb7bTiCVeI
H60iZ9jgAwFFsqUw0pVFjSlTXdk0cHSnGopPcS1O/Su/DOXVH5mNZZECG2jUGLMd0ZpgcD9oxz3n
lS/0dta6q3EddciIDRaKI2eMzzgVgXZ8Pjml6USqZzDtzfEpWZ7XwKPfg10KrSBNyMZgoXXG2SOu
54CTA3AZyx5KN3jShdtHfb4I8CD4aA19lUgNbTzk1GsDwmkQscirygqDucbC8WV3FnCusIcaxj4f
PhxnV1ZlL+iu4Zz17HthZ7bpbWJDUmsMl2n5cK1Q5cJ5ytOHirw8dn5hHKjNPnrvPCE3B0vUqRNR
zT3NoZ3NU6adq04LzYlw6Sqi2qQustdy+4zQLru9AD0nnm7ieQiAQrAB1gpgedwukPDa6KNhgsrl
WXV5YUON8e3Dh8JAGQHgSOicxV1qV0Xx6whS/m/cEADZuiZkeAZlEBNhadX3L8WSpwBuIEqr0NbA
KLD4KD1H4OA8DfYr2UvZYVoAyRtR80xK5i4CcChMosUDofmj5l+FtDzrTXbq47Lf6xERhYfVn9/m
slBzV9Z6ijyvGU0bCQNpjhQ2DGauXffMmDxhR9NiFcCnCslagnQLj2mXkSyijK4u9o5zHCue/fBb
2Y3+EO/Sx2gLUVQPQvv2kh6EKGAAGCuv9+0YkjxLrzsl4pDFr8Fi3V++e51y1r5aQImbQJEiQ8EY
/ro76lu80See+mpklRloDqZSQP5Rna467fB9usaKbE+rd23w1WX7SeBtAs6Bm+xudi8hAf7W+1lR
9xT16NnpspsOjwPtXnoBmFoSVzqEviqWEolald2Rc0R4dZEgCM87B1UThaO4UDtIoLuj1CkySaOr
7PgC58P7/1Osj8mfmY3gowY7kQ+l0QdEJReMQgz2LvfBpKEg0D6/j7+gZEKrU4hA0slqSqQqvqZB
V4hUIkpoQH1mWymUuxiKdKy9xPYDARUxoEwKSL9C5urjn2mQSesxQJD3gw9QybC794n8uLukblq8
4D+YWUh9izL0rYfHtYx7XsD27ThJ3wguhLaLnIhQ2tcAv7eIrg5iJxVK2ngA4VNjQ7Bt+m5qqQtd
/C8iIdXCHoK5djNPiltLdXj/+fjyZ7O/O2+hqg0i6DCRcCvMsZeT0RDKa62JEW/WekENI0foJBpE
PmwoZp5+MtGgnlsGZ48FIoZpD1zCTrWHmhn+uvrkN9okd0F/1ZAON9AeCLu0JGSZzY1VQV2Ehefv
sbES2xotiyl/r7kzerydxPW+4cT+psTBrO/NCejzyJ5LoTQbWg5mYa1iJSxyVuv9zaVT1tz+Bf8l
s0KTZvq5MWfmh7XHaVcManqqoqw8H+R3DdPBo+2APn8G1Zziunqb5m1CQFYMiyRkmSLB1MZhhOUR
tso9l4WP+WlAg99Pv9ZI62od5dRNvCEz4zzjUuGdKIkOgVt/daNRSttpa9kKl6e0/0mcNgZGaQ6z
mYfITv9A7eIXIfIWfe8YfqiwXmwdbUuA+9E4cmA3rIk/pLw56tNZjYkPjeugXEzGRK5EeGCdx/rj
CkC6ZDx/VRWWAdkRQ3ry64vKYhxN4MvZz93wrlBqFNBbzy9GwqTI6rVPHL2I/HG+KaSsvDoZ+S2K
vAZToj4+Ab+dBmgLEB81T0zZQT3bIt9tpxuWVCD/h9Mi7puqbNmIFOrdQDmuowxa/AA23ZmzHofI
Ov8W9QyfqfXiOxjRK0+wNhugQdJUWq6pyUQ0YWmgjpbjf5naT1KhsbXne1bIvNA7ZLMuOK6XmibE
gFzFibaAwpgQElAsT9+u0mqK9/Hu/q94wjKtic2/DM1AIce6FGwWEXqRQ4nRnDFSmohg7GyaA8Sa
K6iFanNtn99iGfoebV8vkUt6unOUDVK2ywrDq22p9xvAwosu0sbFc3USvup9oB6wH1V+4GY+53TS
tPtQ8hjhd3znKA7OjloOKkFoZeKryUg8HeXWXgk3lSfvRGpwSKfYM+XQLthcKTQi7ao/i2MRwczl
mY1ZNW1FBHgMhejiStpqCTNrAdjGmysdWQgiywIDvtutaxyIT8XoYjsKDuLh2V8qT8XJJnN/pSOF
OK89iL6AclkLyeFwo+FJXZOClDBLhRgn3DfHnGWG7sRvbUPoaJRAzBnZWdNldzpfc4ijJ8LzOHZA
6tsvFHip/ZHsY7QjxajAXxbC5e7xjKuJad4kBf7Gv/hGaro97PMh0twR7V2KHbTebndFQV3s2BVY
c1lSUD0RMvfa26d/kcyqYFhZvQj4i8D33iVsVsT/3fqGLyksAc+w26qKYyeyPWys+i7riClebXGl
ARYfcPiDu944JSBYTX0lfKDrMLKdt1qb/eyWoxDhc+Ij6OEWS3Z90xQvdiFmm1tg+5KEWulGS0jH
XJN0AMdS5mCFzORPWEY2UdYC7E7QFQBgIf9go/PffwAM7X+caMi/BvyUrE/bE548N0dnKJHZP+nE
YayNnn7aK/4AxiHAecLEt4rNo0mEK9we9cVoYEPx5K2zuPLmaqZUCSmUTzVYk2NPKw799ysLmQrA
n8oS0yHdWy9+ZbtTogmyJ3lVM3VvwOmOIf++gHqeXokXE3ibg+6sriS/RuLcAk/CL8R+DeSaGUj+
e1yyXnP0He0pW5BjfsXWj5rSmWHD9Nx1kyp64UHHiWBPDXTWO/sjS9JJ8oT4c97B70hconFROurO
TTQ9Gl997ZNmjwJVd178Djg8cJAu/PTFKB+peUckQ219QKop5670UyxgsFFJPVMifnseXmcz9mFh
yPnfno7r5Uq4WFsSsBwKJblf5Ccd5Lc5xrPwnjTUE6H4NdwbmcwxiLwuB8m7Ot1ekOXbjQSfsXfj
E4bfETHXbxhBU+DXlLFBTZBaTm4kzcrRKmIAgwMEY/ExvodqiQcIM0SiLFL+F9uCzbqMlpsS5u9T
6vGuzlD5puqL8B55+1zG48MKKsR1+WTOzDP8G/YFMU5fyQtHyTyQO0GbTSkgmCc4NMKO7UiO/E1Z
6wDzxIXX03yUD8EY2D8uyvtUdDXPBs1dxrUl14P2E6pxXs9qSJiNRCh6ioW3OhZje5LLHnbB1Okn
hOOhbPae5BhQg4b9soMGFv5ValPWbXEihdOQc1lzPkwb65l7N/b0ai4oDzB6uQwBa5O7m2xrlcHN
47/qdwZIgIN+v/DFmgd4sk7WDoDJ2oKG/zpeVZopX7nwFf/qTggwSwJj3sHmmSOOjZjm6TSHMvb3
bafLGeoY7sPNwRXbQPV8uE76Mz1un7QwJGQ7941s1YxRhkL6wQvC1998fFGaVu0bBqKdyxjaMbBK
kfp0eeD09+lXsK3HlwElfT19idl0FMG5YMA/M58/cDZiJAIzq/+EaDc13J8TPtmsKjqCk/ZVcWPk
uRGkw/7nRU0agahPRd0jLzRASpL4HlYfEK6jFwM4ZxR5VOVJWNpizLBXlRbbN+hAwbLiUt0VYR24
58yZ05HDPLa4uyalzShFJ8ZIYX2WZyHRqWmEQFYnu1HZwgzStSAp6Of2K6zwJIpN/aQZ/OWmK4VE
51H3foHlQcWmNDnrQwSv0/Bcp1RmzA6sp5WTrQ+Lvp2Ov746cjBfVZ6oB4OW8156GcDq0eVkZOQU
+KrxmJqtsIHqpAaMNXa1ooWSfrPrW7XL5IzC0yasEx46/+XbVZWhHAl4SlKP7qjuzQShlcA/70j5
WXNltUK2JVq+lF8w+PzCBjNfcoFugG3EYt6R4fx9mcFiHD1znqbUvi5f0iubX1LNb1tc2juOJEf8
RaZpHxJEyWj8LsvhvrKtOGEaWHfWDp2ZLdAxrFyC/qZPoTcvt/wpkVbt5dm12pJUCu5Jlu1FdkkD
g2uIkCzssErcg37DxRIRJa6eeFUxkV8rI4Y+gx4Wuowy8tWpLazhjktS3coI/jXDVQVpZII3/BsZ
i20z0ZuURFB41cwFP9A5EdCOFCX9x5oW8UQ4KAtDXrS4D4inrnraXgmtlJOSzSgdnxKPhR+Lljd0
X924t8wDMhQ/1vfBsJo5BbGYFSAglxOZaykcxHXLr5Kycm4vAv9fnoiGOGdZkxGMxVXumvKMurXC
IueVGMxXc0S1cNlaolSCwFq1x9OvtNub8kFYjuC74+TBork580rf8NXuDmG8RQQwa5/AMCxUdr6o
iPp5FLKzDpcnZThqIp5VHIBdd6XgWIs0GapGeUJ4rKhFpHIWHBmGgXdgyHwt8Q9ekiPA1eEgLcPC
jpP909XX+HUMO0lFrCWqorOxjskBlDS6O380j/VJ9pgKboHD4PXxILn5o3+nrMUQFmEZQHANcXHr
ZRHpVHV0pz1v8BgP4Yu5KiCqmruGlZAS6S6NjRl8qW1vFUKj0PbzOwpCZ/sGNkz6qY1UU54XXSPK
G0PbuiAlQhtxbCzT1ogbufAiB+jbL5NxE2N+Ybx6/JBhWKWNkfluW/rQnsnibySsjPiIkTBrWe1W
1xtdjtWAOXbs83cxdWAmFGpQ/p92kjNAsizDw2XGD1B35BOXWb3XiRWTQ4/gsM7iVnjiwkrny5Nb
T1WlqJ3hW23KHhq6BJfogUPLsqm2y2pWI0+unwz1BCxcMGtXhy3JVuhtYnORekrWy4ncMMpNvyGa
w20hOtjEXrvkaPvXTenEfzhXjkLOzTQbELF2e36bngZS8i8WKuQ1xgeQ2lYTIydZuJSS7/IuE3un
HKKEfXlfs6L+ueUcTS8EQwoEV/vmx8alMngjWVg5eHEbpzOPzW9Am5h13Q+HGFjJw97nNsBtN8u5
FcytLbkB2xdfztvQLZAnNrww9pGl6yiLcZHi/mdlyeyym/G/pIdgzFrq0c7NFJ0493c+yEqHWKtR
WAWB6iwxYa++1jMcex/lnMD//V/8p72mFM/6T3uWJq45JqCCzzszc/4FvJ5E20CGnXokzVCdbnRE
OncPuV2eul3dEkrDb4qvA2W9kxJ67BQIiQeugpdYqWm5wixA+txGhrSegOQ7NV/pU/LDN7P8LeDF
XehDt0bUxgH9p7mmQvkzpch6O82l1lDze8BlSgaC9KhqpRIp20OxKn53AMmIuo/YXMsnXz+jTY35
HyuM+Ayu5nGpz+qowpCHe0+TRfmHicYYJrWXjyydLJdgOKLKGkMWXyIxYTD1YKwDzWFPfqhyjQjQ
lCaiM841nBEGrHjQ4b2IjJtjJnF4WwVB4pcoYzzdIJTTwUecgSiVd+QorMUkbgMGlGDMrWw8IMD7
IVFfGEZIbkM6bBysfhwrhSStMhq0sUDwyqLijBRV9KOTy9u75QWwNCufhOVO/yyDIaLLm7wZj1C+
1YZM671riAGct/E57i+rpIYQneva+W9ya7F10tmrfaF52awG3fRKldjvCNl4sZPfTx80FKxbLVOa
TlmzVQYEU6eSv4M7cLu275cD7m+433G6bEXKZBsQ3R7/Nn8HA+eQF04/w/OA56vGKpRgIZqRID+o
oLzW9glhDF0IEvZOjccdvKtJ+RgYMe1GwUk6EWLex6EKyKCopSWWUXucXmO+lbxeNkEQdlJPgRuE
8SfHTHHBEIFY1s3xBubCVk568IUatMrm5Lf7NPi8FADxUsHkAmwnRcZw36ObQSbF82cXjeatbFHs
T31/DrLgpSsyKdtN2v/hDb6WDAfYH1WJ+ON7WLHgGBRF0j0mQCy6qO07RIfRQq+gD5rRalA/YwS1
DruR+ninD/l9oMJaO8iaManw4JSBeMkjCPtQh6me0S0pYAfzmhXtb49w95n8rrs7roOxCbXjbBPi
bnFVLb8Ljwg3MzrUGDsqxbjFqKB03DXKDDuHfQU43g0nM4ldpujB3M6hEgSwPjepYfk3XNDX1IMy
q2gLPqFkJ8nJREg/PNXB5ba4Nmmqxo/sRZO7h0Mj1TTyhW8Bq8tghScWJ4fPWdvouKaXP3V6dJ7P
yykMgu/D9ptp/BS5b4n4PwpRaQRKYe8Hy5FQCNS8Uj2LqXqjP+CJOnwx5lYA5jTLY/QbfLIhJEWQ
OcqHz1031CGjvqzhugRI+k60LokGYOq1tGczxJhx/YXm0ljQKosA6tyRGLCAZ/QzNd/teI+AjMjU
s1cde6MpG5aJfIsUU8ddFDaVGD1THR5kNCriBliFm/KUhXcZag7m+HGq3sN/IEkpB4/JlnHAZl2G
U7Q/oTKcV+B5+gca/nXlbNOR1tqyC2xl6RN4WWMJrNelox05zRVteRqz9C0XDVmnSV7t6aMnl8Dw
uVNoapf7gujP/G46bSlLufo+A2FcSGJH+VzgdQ0INQmKr9c8pOKppTXaJVTvMCdk6CrtvSoZ5iSs
0N3/6KGUSwivsJz+sQ7AAjte0RUG3FIYZbpoc2fdLsw4p6k0mqxIYYFPGvSkoUhOdtIRzg54tlVy
d5CznwUks52rqTSBDT9J51ADJ2j1hrifjQqIQk0YVPGmo3lMoaaYLITXawuBFgc8S4UCx6FU8A46
crzKRsJzyPA6tR4f4/o6dKQLFX4JX6uPse5ly8ZbTadYVJNWMlsnRobiA39iBpfkYy7VYJXgz8Z1
3sHvPz3CVv3xaKJr/I/beO5moPgFLszDV3bdmip3hCFveyqNzUD06N+sqiwkybW+dU9jiS1ukNcM
WmV+9rdEd4RNjrsbOhAxIrxuHedxIPH1A9z5+iQkvpTqVd8XZ8o5u1hZMkMI9WFhsTXIfq+jkP1s
n25ojPe5LizUmxmy5d8Wg/uLNN9SeVtqUPXE/piJ8rO0TbtOQVwhEtcIGBl393q1hOalKBloOlyc
Qgc2cxFy0DX/44f1rztfZMHWFl9veZWttCe/GT7AfhVi28WGxxIdvMk0vkeouj33mK7RWaSsrosa
8zo/Lk4g656nLneXIapJtVSqKcDwd9gi2K700Z4GPGnVslcXccHoogTSjZD/cgaKxtYsP1ixE4cr
l4mU44rENgKc0SMh0X78Q4qHOy8qs/LSrp6t6bvJx2AAG9GyiiulS01D9bjCBi2BAdav7ps5qZ00
Jyyfjq+ckL7s1OiHw6QawrQRFeS1wnH11AnfC3fhLZlUj2wNwJnBofjwuGhS8OinrJfLjkIM+167
/AZW9aqiet48rRZB+kApiGGp8kk+JjI8Z246e9P/l0rqSk4Mk5FX8kw93f+2aAu0kjig5XTAeAZk
xHgYguTiOZa/8AGcIuf/T3NhxN9tQJ+g+4S9Eh4/u+EWIX5OJuZJhlUYKuUFht6AxmvhHHacMxOP
+7ZKaQHOZu35J1U9Kk2JvFn7mnCYHDdIcaUeyMIbcl+DWaXn3LdvUZeax1R7CiETQR9l+URvVmO8
D/1uawHTzRJQHfZrxGvk8vwz3/L9fAo+Jsi/ywxyoYioa9yKwET2wz/dt15VM93wc3ZKRc9XMchB
O04plEuRMU/K1K6hCeR6WaVmVvIXfKGbSZZtt++W3/XXcNZuktWqzqVuv5fxIvOw7U3DfW8R/5Oj
cbkiVDY2LYRuOwwvA/Jzdi6U2gMJD6VYVmm6/+gJ6snJUzDdUBPuDNI6jOfUM3SVlq3buan+X36l
vkquKNc/1sbMIlzmn8WsjRIvxpT065o55mGb+I3tMeNxERTY+YJwaRzn5vMF9GPvV+oLYd/xjfcA
+A0nJhhZ8MS1/tQDeOLPW7VUqY2r8QT6rvOoujxuoWt5SRmuDqM7Lp1CTwGprAJnPNgwf+a1SwKv
PggiEBz+aSkdoYSrQXoje5Qw3KGjF0mUPcoJnASY/M+EkgrDPPSO1esc/sUyhZj+Zbx+xHP+kdwJ
5/ATURestDCC6kkv6sgwrtMZvRW/7prJhhDbhh9uPH+gyMdPrT41CLUQhPFmwPWn7+XzZ7XyjOHQ
RnSz1qGm5pSxYQcsfWZQZlVTYutDrmEHndFW4De0gTaC4JZPafps/Fr0osW3o4O4rWLuoiNsPEWH
0ckIVeo5LxgxDgVQGksG2WsfZw+9HVq/Ug0ANcvbgtUbvTZvtdjTJyMxG/XdJj9vwMj89++zXyHg
1MgVsrpkuOhol6igMO2t1AbMOsvXHpLnUCjxKO+S6I4SqHVKOMUfQWLdjojPKmaDfHW99Sx3eZ4t
l4nQoydko9BgLQoYhCJPeSA63vCRn4/lYGDIoqXAew3RgvkHb+1HtL/Nc5LX41NdOSgWPkXqGUBQ
MEcs31AiEWzOM1oS0yqKaAKs0YiCkEgkebNkAcKE5el5egiztCXBCyy3O87XgSTjIY5OoGUUl0Zy
fGo+GjgtSEw5y/S4/SosBU4rtDvI4nPWU89SarniD0GKmFND55H5Q5e53XZwROSTVAzznZOZJBvi
i/EcDWf6WqhBgi8CM2tOMFDgmBpmUrEE0kLqlRjJI1HPOvrT1mCedUlLTKDaIiUhhMc3jdjE0wA/
S1KrvGyJTHwewqU3rCQ5WEvLe+FUUPiTKyL95AW2g2iCuVlxhU+Gv0q2DRT+zX3PURPDfMzsX78q
asSVFxxX5ebNH6h9pWtGym4Zj/ECM+jlYmAzwCyhNIEURPmjAkUe5YupReUDaKpiG3MyVoaQY61U
aEB+4QP/q3mg0jhn4KhDtFcHuTvwXDspYShmaFC9oHlAoTkIErhUKpMgEyDrqvYi+EUZhYPJLeNf
hFZUm9+sfWWRBzOM+/Ag+7TmfFt/FBO2BltdvhnIE+1vbUytge/U6flvRuPaG/YCpTdnDeXLeQSB
Dt2AAaYsEc76nzw4WnyTdb6oCFk1+imLJAI6oPHvb1f715bd7SlAD+BbO78QwtVG7HZxrh3MYYBv
k6ap+/cw6qpcfR00MmflCuhHBPmVoYnaIsub0zr3455qm0uD9lNJhe/z3a+TmGe3D7yG3GGVdbDP
GwEqwt9CmFdQZ5WuFtvWvPXQtQghWlcQ54szvKcG0Vgd224CRHdpRBi476Sa0zVYU6Bn/QWqRgM6
R68TD9l8kPxUpsznP6uzzP2hs8eLxBkMduHb0LGwnC8LsFRex0+yunkfCPsdgssXrrTCzGwVQJir
mcq7bca5C7DIMKaf2wcYT55vz/1dQSZxbA4oTnp1ss8ciYygtYHb2E26HZpz/wQUppleKrR7Nami
Zh4DYS+rOSp1asvdTYKiXOTVdxxZzQGmRapZWkj9MLv/6J8sriSDwHot0oGypxpsYdgcN0YWJjrV
PWTjjAl6WYCwlOf48ZSIBRA/bHTbt2WyYHPn/W7lwwLXz6a4m8r8B+Pzq1RULhdb8pHXe+daNsO/
EmhVykOd6eQLc201eimiCXEU7e3oNssmdgj8ngTua6Z+nY9EepKun++2RDZqaKELXF1PJbbPtVFa
1HGZy3PmWFErEDhEotWg6i65E6J7XPDX8YbSc0HTgmGXXxcwjQYPEeU+JBEeNO2REc/RtOxhMjJB
zQJp73b7ytj9BvQ6hk98AP9WXwBKamSMkHMwm9HcdYAZPC7i6plc/zRB8tBVJEywAR5X8DVgtjER
pT9PL+jVlzgeN2QJ2kSEX71GWnB1oQo0E2rhc/9PsWe2EnoBpmMzOEzh9L9SM+ybPW2q0F2N9R4A
zRjFm4S+vuWu4FS9TYVTcDx+tjW6khNiWeHYqhaNsAH0mjqhblyhqDOpZrCPqmteo/n4fwZ8fKZ9
jmb6tJq1vFOLRstwn7+HP63mJYM5Co8eh3H/wjj9zjjNDP6PVIplKbAJoAWxF6sNrCe+k6jcV7XR
d5EQ4TKk8PQ0k3LMvf0w85n+4a+GuYIFdWISPJ8OV0SJOlSl170R3iuMc1pkM4IFWeqUTTVkTVG8
8C8dN+a33WZIRFS3sXwnTWYRT51yGzkCeFxnt/ziw8oZxs6KqqKJWZY7QLFwZsCF46npoQaKo3Hw
wupOAlXsYmY8h9I4nBFnTsasaLUiDBYtsMPpmeu0CICk8jCDMiECz0+BuV5tHuKYOjmFscGl52fS
qsrAOm/rZQC7N3joLJ0CWDV0J8hBCjy+Zy0m+pIQ9n5dcKMHcVJ43O3GlX8nxeRPj094oCwkIFMZ
f7mLW006jpk843iqQpjnXS5dlJUnilOhYIsiNUshZLwTPhcowtEP2u9bm8kJMo76/cZCWJeTvAV5
vQItLPcHzciIr88QvOlXFasWiloSfiYkBdWe6jF283M8YoDNmbigovctIvfUUphwD/HLcGwdS1ZL
hLXYwdb/BbsQw/PIJD2FudUJdlCz8atpaJxr5TbjaYGnWXMhyQgjsbF1FkmGdza7PT7/u+9nMJ0F
k2Al/vsESG53KbNwP9kh9y6olblGD7em9fQW42kKkBYXGpPjFT3gG/RTy/QulE0mjQxrvSizpVw9
W0l1lc0lQSTm35wLjG1bF7RtNU50Ug9zk5PNAHLReX2ymFzrt6OxManot/Mts+lj09Utw7S+ESKr
qWW8Rw+UYVKmkMNfL4bMWpVqgNufEKuepNzJ7z7owOMNCNI42vWdqKPOzbbFYLAShLHZ4UZvLK5i
YzazdHAEOmkuFZE6GEFMvYiteIu946Jtsv5k7MKQFuqCPwa7dxZK9wzdBZLfLpbuEVkT2grPiKTN
jdQWthvCzGJaUrtLjMhs1q3dmXLP6+C15nmAkznJ2cUH6CQ7PjDR0DpgAkhTdWVA9EmBDnPVtqxq
5t6dNSlyB2mCyRMIqXu1Nx7MDPGye4zC9jrWkA+JonQIDrmsx1D+fhU8RByElNBT8Dq1OZ+0O7ka
XrhZlFRApXULIc2f9WjdVxRc+IPz21uBoWTlJbxufnDMHgSd8EXrLLi9alfSTD27eI0Ge//wAjg+
uSYG/BkqyJ5pXz83bVX+WSic1XPEUZRjiiZLPZk8RwQ5oZ3v8ANTJS0YlL2SpqHYEpqcMffkK6oz
me+ycmBdI/DkwxASPBxnCmo3vii6+hlVv6jzr++FM5ZjWRAweP7QCkrW+Vy3UWV4ddFd2USGBWZ3
pBS/isqZC1G9eVjQbi1EGbohxw8KV6ZyRrtiR68uUbaLV1cQNbEKvOCgst4ey7UoVJGPUz5Do8qQ
/XsNvlR1JU+q7gbVo3E/+ET4pNED+GClLb1HJLr2PWY4qvTtpI4c+5EUOklbkG6FLO69rZBHCMsE
MVXo1k+5Zcq9iAxcXex3sdRTBNZkTO2hcBlq9PNV1FEDhBk2PftUi+gZ/90xKpYFQsj5jeJ5quY9
KBfdZPusw522mZa3aZGng7NIbtG9ZnbelbfN1ndAipJazTX3EQ8sIdttQzgBRhOwZb+pPl7tgmNV
CIIpurMKN7E1Qv2yozznDrO0Ek6FI5q0SoiAfhEdqHzq3/Nlf7+7B7/xxHY+oq+ADffGTldVxqDu
5byM1sj/3O3BAMx35m8L987/VY0ocXlbLw4vR5n3SAB9A3aQzDgq6k7svzrwg7+uXsL7VQo/KCrd
7L1PAjer4XIKJF7W6zhOSSv9vFyBdCTEGHBulJ4hQrJ3HFxYT7m1tUBczEGqfiy42J4lb1E9KCxN
V14HiSxtEPNxKt4y+d1NylC5I5bze7r9/z2t3t2LNnpDbbmiTQMVL9ZWjgkfCGPl/FeDRiMP5htu
oTXblTSfVqG84iLW3L8HRG8B9EVdOyVbin0lap6IBS9/fpVtC4Kp9BDCJ9po/f12ueC90OWQnrpk
c3t2wBabSCSWB7EGqpzF6SaVNxoKn6wr1S2YVCOQzSzmVaveyAhwrhSN8yw4cSTcuHc++9tj/X+i
sTkHA5xysLOI6rzsQVK0/BInvHB65szHcobDVS9zSLBbrReo24eJ9BwrJMTYguvSXFth1mOIJlsm
SP2Pb9iwJD9MJFZOXRh78fvV1QRhxhC4sGXKgLm9AFXiKfFV59Aty8/sGOYONDMZt7CI/itsysqX
IdTbWBdE4aejmBMsuD/leQ5UEZwZlEE5fHzifmca1mRr1esM9rRt7ZWQDGZsIMkYU11+lP2AAzTh
OBTQQ9Xv8o8+vIuZ/C0f7hbnZdbz4ezVrAVlQ7BElYNy29ZjGmdLVeKNisr0DMoiFXSVM4zg+BVW
aSKahyqWkYh/oTRdocNUYnBdhpUEHQ+0+xJBbhtejmaVq/OlSOG/ZMAiSJQ9TpGEtS/HhNk69Vra
id6mUZF7iNaEuslZyGztQD+cC2pqJ+aHj0PnbxMdpyAGz51IeW6UmdEaRjqGG6B7d+8jvxiW6P7S
o6P3Ne97+0bsEGZz71TUtj1NwNKKgQcMGu8q/O7S8b1NxZNDpIiClPqufpxRlChovgV58S/CcHPG
HhgtcN46m15T+pLq/OemxjvvjEyLleqe7730UvQOg1ityRztuXmNN2faO11sN4E/uyNkFIqVSjuc
gBQJ++uhSuegL1MdrcDN2DIEHidkcjpTSda8d/9bvN5cjO/HldkjnYRChk7C6NMkAJfIrPifosPc
Sa8pSSWCBkXsMuiozBGWqty2DSkoQuUX5HInHzQwN1xtCszOXxB49cyl87fqFA03fNVi88Yn5GC+
uHPf1fSzcJLfDFD8dUw8uKgVYF8/I1s+q88KA4+E3U1c/gVUQSYNjm9DD/cucWWZmVZNT6sIGi13
UdqeDuTW1FMKGqjkYARWPgXa48fsQHGFfnDTtQf7Vwp2OaAWsAufmgWMBN+n/R2JSYny5M1Kk+B0
s8rO9RerOvQcWw07bqCd9GgIEDj8r9jJhEIaDurZc+8W3e7yeq7RacaEgEF8XVGfH5YAdn2ZfXky
6JhOZ2mhSUNq83ko/yfidqvXekLx5OYHFXK68HGo3LdJeA12KLHOpPoiMYaKwarnU44bbIhRYJ/B
rfzNZcl7Pgh9v/c1RBpnE37PZ7FBcfstMWDC14tRgz/W5IioPo3ka5idDB7hMsQ6X+vwaQZa2WER
7pmWyix01MA+Jln/Snvv+uIFZXC6Rmog/tvrN+q6QJzzmbg12Hcn21lzY4uaxajWeeqIPWGAJnZv
6nDGUIEUE/KeCQZCYSYGcnkh7mmegTzX/dKp7SyeYvkm/rFJeQEZ5GzKAA4Dx62P/oI7lbxjGdd1
8QOEzkC7OnE/mF4B8zhDfva2/98SuTw6v7dtkAMCNO2jgrHV5Izf/ESWHeZbJM9ddR+Z8mfJnveU
9t9qvxEGY8CzKsK+vLy3eIop3Ks9RXHccmTTJJpgPpZsgdOy1YvE85pY3vO2wVcE4ujpTUenFrLM
WnGHM/xqdXWptUBR4AXTCR/3RFj4fCAcbRb73RY/zLnE7n1K02lEYimCUKLyZQtQ+xXzXubfHQ8Q
OhbnXfScP+SwiCDpNzhFSQEAvYJtunJzrzdxRqusXcAVYpaHFJ8XDFbh+8ctTskbmYLs9f+JDlyu
nKzbyj3dqVzL/8GTZyiAYEe9p7x3yUqlNfzc8rKBHAaANgx3HVzgeotwrNj3n24Pn48hjBBetbWM
faUzQSIjYkrcjXA4l9x4FHX4vc4XSc4s8ALYeRT6+amhIMulLA+hU4POvmUIsFPIWDtIBDU4wZeX
LyFuzbqRgCbFZB1isicZF7j0UlOYlxVS/3NDFvVi23ysj8lOQSaocQeJnNsWpxX1hPmba6/FqXGs
Nmia0UiNJWj0L5XsLHWnu7rbGtrwoTupHRBjx8Ot041WZQmp5sdoP5mIynd+ZvEJmRTvfpklb7Mh
b6fzptqBht6RhrkzXaLlQrolTyHt7fL2+6HYEybAHh2fVhWo5Fa8jE0+QLa01MH7aDmQqQgo4gaQ
YKPWxdCAGqREpaHioF+vyKVS7qdpqMvaMQwHZRlH8JneBqFEYB9w0Jl53v7d8bWYNz7LC41aplE8
1Vt5ltdPT1/XtOKSnZqX7gOFX3sPShaXn/85CgGAFTFFnk65ZvCMTEm4kadMY1LYzMElcXY7VZfW
1zvocZXtkurcahUeXYsn6mHcZrzSQRK+IGeAa0+jhNSKhuGezU6b9IASyQIp2kGc0tfd2nIXgHgb
bZRefgEgf3HaBpPYJWrZR4MBtAEGBgWouAIDNzCAgzLO/J8os1eHf5qkVWTBu4Wajan6BrYByxXM
39Q9ItZq2RAay/yeS7FtXw8ADw8LFQ8ahIMcy2IJunC5k2P70ZSerEsjU7E6U5f1dq3G71XG2HTh
zIu9lGD1IEVoSGe6NUxjaxuvUST9S2zq7qP5RaTJXOWf+H29UXIPZHpCTzCOGEbzqev84xJoPMUG
UMJCWJpILOW6UPKYC9LK1pzuAFosId3kc5RdGONC6QshYHxywae9Yf9eL7mPR59z4zzBaaPRd/VD
LNHO2XGRfr7lgEXtl3FAzdiRsmlW1BaqF5NuU5h0mBzDD17d+ccqjYiCxC0A5JjbeNIvQXkugfDp
q1DbhG6shL4oR+xHOdXYB9KdwEY2QiK5+2TuU2h7VXYAYhb4ky+ZArN2LGpw8fvhGnbbpCrBGANx
xAXIZeIxPTjKux3rVXycb1IxEbzXpjk9aBVSDMlja0dn72SrqwVDYsv1kKYQCHrZIIXnqvgxaxh4
Sszvk4CBYlKIJgCBRy3x7bKUFOxG58MSACD4CAm5jZXkfQsyVH9FstlIvCiGxtSRdSicdsaqePgb
rE5Bwgjh8vJcK+iznQseSQsdLGy0pAnNnzA2z9BwV29s8O2KcKxDtZTR35DnjVkso5Ldtod+FWnW
JiOmq1OQ/su2QxsYZQaXh/u0pxhUlGJb5D3nYVqbwpewM+j0FL/Pe6kO+u7KWC10F4u9JslLJzPv
CLmvFthU7eY7khixUIA2U80a6JJYX6jn0y58znY3vwjhs4eUnWeiPfnjOlmZUU6auNLhFCkMQbAh
e/QwGkGCq/EET/m538pGKbdxW8m1Zno9tvpJ0i3l0qfHum28ALjt87cti6fuVBNmwHurHnqDKgnG
oWZs+E4amm3APGCea3uh5UcGcRRrFk+YPgRY12mMPtAPBAgGYDna4EXLIanc9Dw4jQ/s3s2OSjcf
dy5k2gNUaDPhSHoOBavLwHZzGTvcSgMZDxmZMl+4NNZGBeNzfT9d1KQKwnz+VuffXOf4paNf2fA4
7NcpMmGRUJFqQOoUABc2OJqcjVdGPUxsF+JTzxE5QuUiJJt0+ieVDX7f89TS5WK9HDgt3IlXvhT1
iQuwQgSJi41fJVL83oiUDcrWI0rhevxE6mhstkYqLhVE1G0M/75pUUPHcek4qst/ubr+jUDYnkW9
eKBNN+tkgzJx0buw+blVPNmm+mg24PG6BXtSeygmNZqnwlsS0dK2OplCpjHqrrmtFjEISMLFR7m2
vx9u+my44ds+VvbLl3Px6a4zdHienyAPQwG/Iob8GwOMVpRPBBBKBSAbgj36THgkxIuYlt/q/Dul
qzVXIrf0jtVn2Z47B5XVYoWjf4et1JK+ST8GW5kRrfu3R+LnXXsy8JJfTR6WBPUER2mCbQcQrY7l
xziekR8WP0Nb9YSQ38t8aSrakHW7O8AIuDudofwtd+FyU6htCRDN/5zE7gjsPHZg6h6agn3FoFvj
smApT2SbOlzSqP7/xRSHpz5BBNnj2/wGczn1iNWUm1wLpnz1MmoUj3HTWZ1i6qxrwCjOQ7LIV/7Y
iGUfnbQ+p1S7jh3B1eCYScDNaZoD8Nf9v5YYUMLNQ+YI2vopImuWmr7whaSYNmSNJbNK1T/O3X8B
GKBZcSjMasyy0za0AKhFqckhe7y+LCrA2sqrhFyI18b9qQW8EZsaojwXaoYpCOZSyO9gspi043oV
Nbv2WcB/qheC7EVN9TOJ//ptfpyRICXBTJdb77ZUuA3EXEDlKRn3rp/HWbnLAdXqCB5Z7b0Gom13
t2sMJeJxUkK+3Iqak6bgncbu6NyItkx2RrjDZIMxxpMVWsUR3noU6/o2qQhPkz3tHJZOwvi552nQ
Lv1pc3AJJWw7Pzy0oH+segrgi5QBrAg+PjSuI1+16SaRXgLptro852IMe8ZSCT+HKsItjtU9V69V
uuGIK0oLn18TDsxA7CpGThHER51BapgRD6CRn5i7ZUTWjj0K8BMuLCkxXIOdhVnDWrjwj5IyBKgL
CQ6HY3kAWXFeH+2VOn++6+vCylxKKeubB06kKTU2Dk2+8YRz1TVjuSY9Gd+wHYyA2Cf1lIV39IHX
A3K2S8sBnvmCMNV/L81jE5Sw0A9M45v6hr+YYowGqOIy5IHyeY4gAmM0ybU9G+bl4mpmd2evLDu7
u41Tr/LpBhiDoDOMRneWSmcax/pXl22qrLNxHsnHOP0cngPkSNY2FP0D0i+e2l2ECeY00qLYfgsq
FfCtgTL7/+8XKUDLc8cMt/cmViNROXqyK0SzO/5SaYuHtpS78PItM3jO6XjHMNBNBiTapVvV/Pfp
IzisqBtfoAVf/HKIoX1IMUFmnVv/JTBJudKIGG6DgLAZunV8F1LNftNaSuehXG0IeiXsRBWJWbRe
2AXCzqycTRL3bv3iWj7X1AMjCKLxW16a9XOnm8uieAUiCzAxg5vUjeyiDd+hCWM0MGCwET5Jm5H9
thKHSiCdNswziOfhAEairwoiKhrquRSjoq8o7FtktHPDH+BCq70WazHJ+f1GbSQgm3g2BdqyAAZ5
QSv1xz/iiPgEwDk4e6hcxHPiFsaHnzW44jg4F2M+UmThkbg3Y4a4S5Tp+ojNSrPmPP4KdSfeHWvi
JSB0Yq6uFlDvmUh/vxdMG2FTDbR2wlyNXZgLgx5P4XejdELF6i74PL/42miLZsANk/Hy5ZROGu34
tYjw+nzB3LCgV+wlk2WMfPjMPyRquOGRDxRZ7AJON1ASxyCks9BK2lg2WnV0WKeWVtKobBC3fQPx
RbfvyE8rCR7ivfHXnIljnz9St/H0GPhgmBe3PZDfRHnvUTZJwVWDy6JL9yymBNqVjNhejxjbzbsk
fH+9E/fKkGoQy0ugKCj+NXMik0IzbgOMVLBsW6BwfrJyvzKHG4ZnLUfccDJSo+vdo4feWahWIML4
uUBusgDvEhPYqGVa/ksKSHv2MBiuOciapqM5+MLtR40/Gar7V9SfCjf7vpsKZVOJEdu9fEW3Js7B
SDW3AktGLGud9ER6UGBpkT4JtUFGBQq1Uz8ZaI5lgLUSmXv8Do9ubK7p/eysfvTIQrwmp4Eq01Dj
pMA4tkQ14SQWkD3SkADAbBEo4nmxZCxrtKFlxGfDYyu6l2v2s9wWLiPxzwPgoIu9LhBw9BYAVIzZ
8ErfHWTHG45qLGBMnHgFAtuzonIJ4XmOvbTVW4oWIiodV158NIfwnbJ5a5iPUK7GRxP52XwX6DRx
S1qU1xJmOZv1ksIGuj1GAmCvVq3IFOUBEa+OlzyH3eontN6JMuExzB/9YvKbtUXwlcJ8R2OIKI3l
OFdDPtRaya2EFz7N7HhRaO9U8lY4ECGxi+nSIeXOauGyTXJWO4djeuif26HNXdE/PU2xJgwcpImJ
8aJevRntBa22eS3yR/s6seX01cUp7VnpYvVyxIw9K3o5sCgyj+pkrCvzMQDb7fNlPaSAO27m5fBL
OiqfezuHUtjei3jr0d44vA4tm4WELhAau+cI/+dwrvxGKZG94AouCAQk2b3e53Lyg3+mZloSndaj
xmPG3Vq/DFq/wl/dp+vPLF3pSOid7xS/tb4Bf5QF7lXi8PlEj+D6UFpfTx3jNygYYw2ClBs8cTgs
pugL1UflhoTYqL9fVbCC+pnenudYoKvwERYQJJI8lNpzruzOYpvER1Y/fiN67SNkD8ibhheDx3s3
iL3dHfkZ7cOtuCHiAFBRniXiAI7LSawTCT5IBtczEVPkRfbFlgAEoPzL7C7AKHhy56UwqmtBMiZA
CromPmAykk9jTUXMLBlnaD+/dWsMsRb/D++jER1Xla4McKmPZe09Kbumto4z+AHPPDq9Hslw65Ob
k1g7CMrrZWdcs2lZAD+kMjP84wcu2xoeeX8j/kAe2fSRO2rJwxp/PXIEoEBgA6IrJyKy2kRe5GbG
dThMzIJmxRocEfCy9OzxXOW5nMfkbqU21XvzM3BGUFkLd72gG34JuTDoIUKHAnSPygQPjOBhwWsX
gxK59ZOpmvSLZueUFGsdQGgPaT5JVCSXxF7R4VRJwQqIeYneEXUC38GRNS3VSn0BBKaFrrqE8gjX
Am+V0Do/fTQ/Rt752hZPZ0QvC+hGJUQ7ONvmN4+qW5rcXL5kA5HF1YblI4NvdDoZ0aiqviwkk5Vr
5HhzzNZdrHvaUg4dxK/xvED4v5lmq7a7etP2hYBGvPl2d/o7AVSOfbYgKC8sxJQJL0o2iITUHL1s
uiFKgmVhpC0ADlOTBupfFPotFP4NbmdMiC3emNhEiRSbcu7t9bK6cU7MssUGvpBhEYmrcItqBTiC
8BbAo6PFyaEsF18t63HdJmoRdlFkVVsaj3jydAzTTf7LOCu4BA7RQnUXPrOHW6V3rb4W94Tf7kH3
kKT4/FwamAAAQcSGlktDzFW1xl2MMcfkdHTS4hZq/OlfHw67abfnJSHoIz17uiXOjy5kdMC71/DK
yU7erHjTfhTvsp+ivOf38G3tLPCtAB7elaSBvA4l5TMRx7hjDvXKckOzOLXtdJqJgZV7GzhLvPBl
PJjEtMTK7APEOGDqTa+XfxsykYRYVRns3jnPYh5p40RZcjeh167aRsf3GzmgDhgjZq02aLLQOGj8
UbHrMCN+a8xgIUn5WSxmpCPRZ4+Bi6yEfNiyMJZKVn0oMtNkJX4iD73RiM4bIb3TL4ZCTxv7L1Fb
eMHj3xfoCa+cYljZqJdSEbn95D5Zgif5TtzqOI3yORuuifFBg7/t2b1431ghvx3/RVoSOGdH/F7i
KM4XFqV5xvR4qQPBImeCABWpiINyEjpk17ktTkJLNcIuVhP7NR0hTvDX6wp3gn9x9UV+5XUHKUtl
TkcajswxGDv+C2hMkumQapibDjQiFJnJwfTrI3TwydAW4OLrzU49FD+kagdOL6M8RPPhAOvVEPSX
CtIuSeUMDsSQegwYvk2ZCaogKkI+DIqzUZw7+YxDsJvS+w0huOZHt07sjQ72AUkl3zdYpOf7K4l+
tFmmbEd9XQd1I7cMOa2J7MT3/4Vi85Zj+YFsqIdr/3zHoMJ0v/j2HAMQJwXPXgMjE13dvHuInAq+
vaAYlyZ+aiA1X5BJ7oaOq9R6I1oyMm3bMU8sbdIQ1A8tlJA+i4TxjFsrSiLre1qwPfqGAY0ktGCh
u46Duf5RZcsqBTGuvplOsXwcQMVYLAZoKFoVd8cRlqXIyuPO71J1Dt/sM5ZzsvOuC9ubeF+M7NX5
aqbXhfhAUBjWGm25afkYT+lDrCud7NGNrfLHCjUC3EEW1E49tJKuR2AlY3Ldq4OkvBvh4gG6ZTQk
QdwWY4bxltLqmNmrRR8lnO4IEiltQ6PnV9bUhA74DfOBME5tzCRETJktHloLCdaUOfEeIIIT+UYC
k7C2k7lOEMxsPmWNgdtFQAvb7jJhoPoHOKlegXeCiALlfUvseWekpJ3vGaUboiSScvxS31fUICSN
J4SR/uBt+ydmKf86O5lt7Qd/ZNslWy3xCoOMciFLmZQZxZt52dV2ArMrirAQ2I0wRgQ5Z9/gbwbx
bXCFhw0puCRrBx++VOmPMaM7GsYRGxo0vd2sdfwhB3Wmpn3qNI3307DlJVohbGjTBGDm1/rWgVci
J+cKCwYNuigbXb1141W2rDBBU9Kn8a5mamOUA7GXcKQq0QFBxHtmxoayhycvn1FYR8vx4woGOHwB
2i4ElbJBjgsOttI=
`protect end_protected
