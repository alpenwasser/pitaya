`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BeDk6slWwyJ7dkKWyaZdmI5S1xnQWnB2oiiYkvyYe3ILPohOGwb55RsmeeSbX1QjJu01hxqQuKng
/gQKr+nekw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ASzYKVAZmSO0SmC0FWgRspy8UM6oxvcf3jSUzSQ5aTbQcdQEmkCnyOPWPw5rhfBxgGmpUIes9+yb
Y1HX9gskfNW1iUc9hvj0/7i23Dl3Awuv9PwzU2qkFTur1xa+VTaDhjRdBkmelm1XEmzy0fVWfN3E
JrqrAgqGTQHZ2JkK6Bo=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oJBoHreUf2ZGu1uujJJM+r+7FZbqExapJJyyvy1o9iddxQis4QmRw6/bE0DAY0iOm9OEPedgUYiN
HJiQO008872laIEmtmT/BZsMbhdVL80RK/NlqxNSooHOOtA7Q2ooOW5Qroi6pqh15Of2uGz4EX8r
QzKai9gyZ1nNfMdTAvc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gXcd8sTNtxVLLLKC4rAjsRNsfX1NVlxv5NlbcoCN3RLErB2fm8TB5dri0TbIQGAb+HGHGVOVAHgx
uVooaR3J4n0jcKalCdHupCpw5tdmXAARWsN3+yNMWjktBvDZlREeBk2BplNU4DXuIjpyRlcW28oq
fXURF5uCQelaIUMgDwAyoK4ndypdafocPYsPsbB7ZcLdDX4H5Le9tBCnXO/3QcalHHXgUWKcLkyn
o62h+Ts9twP03kQwoK/zsw/Mj8ubV//CFoyYXoAsGg33zvV6pCpWjHcIR6qmaj3YFStAb9Gwjq47
yV9Y3uGyv5WU5KKhj3xqBA2tQXCqQY863nIZnQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZCOLBlM+DOBMBQ8zvcBqrtqtygwYjI0iydlVEAyokc0UPDasfRQj4taurJsghnxG4bETs5xI8oYV
0HnNJr9QlLNdd6mcJgJqN/c90+zI7I0/hnO/qlv0Pup/OiWbYiiAzYaGPmKRDqi7WYyqSO7I4TS2
AG2Q/zR6LKL+UR1LQcmMcJ4RgLFqPmMasX9iUCz5I9lsv9KntADfsOLwcJl5QoT1i4VZKbohe5Qm
MESQHJetAMfbworTVW5vJr8gNUaDSSpP+4845B0JGNCebeUUC8/1KVkOL2aPgIiLRFtWjAGp0OdP
Hgc1IPHx2d0B9ihxkm+YRP31ignQS302EQYvBw==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NrFXeDUSk0IEdKSAJNgkeyX3IOnuNIcPQAo5W4y9LavsF2f6Nt+rduqEQbagw39p3ash8XtbR/w2
nbOm3koCj/8C0OoRET7PqvN4QJy3y4VTXAZe0/S0IrLxQsNhhv6J/qZfD8QvZ356rQBjqyRt3tes
FKIyW/uL9wD45Iy27+yn385eZ31TEAWa3qUWjlZ4QirRNAT1OkORBDIQDHOOlrRwhcFvBqpmP+bt
dB3NdDgt5niwoonBSPDFf2StNdLHNsQCxz9zmE4Hap77op41g4Avc9CdLgPyKBKRlvYKlsU5dB+X
7VzJf8Jl3UhqXRVBX0i7dzEKJTZE1Bhvb5jelg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1541456)
`protect data_block
YzO9pHxtvhOPxb1qQ4BRxlruOqGMOSQRW2duVXJBnTN5CAa8Hxpw1nBTDkTbSFKIvFMi3V+nKBTj
3kf0Z33eOBMz8BCi63B6SWc9IZ65Gn46U1AbMk/qSPgAcfKtM0/aA3LHDMk60gFomTArxNK4o9T5
PWyhopMGzkEbOU0O6OXrBsQMsYZl6RzpnVz7cucwCZrqvojo/bvp5XktLssOSRdNArsv92U3a1gu
XmtXEm0XrZFiiqiVIcRdozfgQY2itPBFH5SwWIY/GecaAxi1xc1ALbrYc9AF5n9tsoQAWZmfe2zv
5+tPtxOeULJBMeRvGhZmpKxhn71+I4loyI14RjKcnO9rtkjuyoC+aGabKUoPN7mjvqJSiAZQQknS
4ABuDAFSk04QFp6ELm0RPKJP7dCv1RkjpUHsfG/mPnqmD5TtjvKPmR2TLKMnk9/KNQ5zeWbdUKig
4HhteNzhz8dMudMsr5c/1pARjmsLgU+wf09knm8am7o6tPowsU+6WO1oUmMfkZlaE8HqCShyT63Z
h2KBl6luehSdinEgBDRq4gOUCz80MPtRti/lpf/9vm5Ety9QjWOqZyLLo/qO1Ofm8YTVVONifAmV
rXYuY39+LMg7AtdXzcz1lSkbiz3glA2CqmC0Ik7wfus3bPtNjzkyUkqG0+30gtLNxzI7ST4UjNZy
AV8J4FXms9wVWf+d9bafjYNF2+PhprJtarOMG652/jHBVwwfWZ6HDxcnJWAJPMbDD4YnrKILySZd
WTB9zpfgK3tRxj72alTiKW92FovCDfaPJ/RrCyQQDfYwis9JzPVEJb3iGuuOv7r4pfWqIVxoqDqn
uFu5nnqvNU+jCvjif/DhAlg2L7cFjOQiKuiauXmqGn91MuDDCOric/tCIqdWiEJDtEbDZSEE8f2o
KgjYBzO/RSQ9/SVOpmmujdSHCm3kvOdrg/eTnXvLZdddmZTa9x2lIF77SKgzILDFwsgdRIk0CqH8
K2VrR4zweNBf1pi06c+WY3UiZKFT6IezGYgsEVEqpk2lNsiGJJQEideVnhDuHsE7MvESILGQ1DqC
MbHvexYQK1ZErTBXzXnGovVOFtNG8Hk+NYpE/J9+qZsOVgOp4HgFaiySv8rzMEvH5UL1sPVobdUY
Y/I/4Z8GzHo2b15O4BArnm0TzNVZNyCvDMnP1Y5mFLDz2o8V+2THZCwazoB63bn+HS5sq8gMhcsM
A7A3FCW164mO70SYo6xkuAZK1589NlJe6sglkQHtH85g22Vxa++TM7lOTXR5CjLZfh8wUjgruS5P
wiHm4cMG+DqaWoq4knqo0puNRl4gb0O3m0nzxFAYUisL85MJbSAFToZUJdNBe82xvOHGG3CBWGBL
DMXjWMW6PtSMhEd6UJE2A8Q+LFMQ5j/iEXjxKuBiH0Neuc9g5X9+kjPpsW2/VJJcJrC2NMW8FzyJ
URweWrSCZFGgv+w0ArOCde0Zzl8t5xe/oQ3FeS9TLgcHdZAO6DM+eklhR0eHrLeO5jxgRCyqlYqZ
c7JZiiEWyMVePPKsp91Ixe7PLNx3eaCRnwPe0mGYlNGvVoO0/AFPrFjjiFjH4VgVtLgueVM8DkTp
Xs1fN2xR/RvdVFgvd8xcJrwdRLy686XgYgX/+PFdotVAJLSrEiPWWsHPKbP/+pukBH7oeeKTVfM7
N+3NfY99p+I36GFHgEuxBH8fvZ29BVYmOUJS/xwdE8pi2d2KyPCxpTNtGsykR3lzcia04ciayTpR
VmQRpqhL297P5tPKHPi9RqALRD35oXweTcDbzo2h8a4517tiEY6YPhW2tsPzd6XBjCPzvZm+MJBj
LR3bLswivUKmx0taVOTH5PMneHFdECme/68VTtB63esLi2GPKC/ZCWU54mgGjnOhNPags21OLk4u
YyG6uEw2Dcs2XsuqS+Qaxog55t7aDpgHaeoj4TxIX5Zg3xqyN04TUMCcJGNefQWs1wBI/0Cz9OtO
FAiajRz59OhD8nERLnYCBeJdT24iG8jhKs74e7QIepYMMpYQq899f8AyLGqBxxRdFAUPOQkPv6RD
gWk5v3DGfUl3tqu1BG+JdVA1Tywn9BypYdgntPt56YF4j/WlEpejlbgN/3j1Z/KAmh+0PCkbb95U
67dMVeLY4CkYCUTzvZdzhzhhpdC2IkANL0HYCpDm5N04j9/zhj+JWVS9gl310qMVhJgJyGyr0JrT
7VyQY82NetR5fi43VFhK09l62pMQLF8VKPrR6jSSR80VFvbSpeYYRhS2hx7R6GkzlY3Ts1nM/mZc
FWWFmvfOiYzEpD8WyUMwzB2uiSfw3oQTmXaxB7ldTWm5snNUeEnGjDJ/gceychjbW0HDF9D8tDZF
PFHwStl7LwvvXDt98Obh1KQtyfuiTyucAsCa41y1dMxf0ltyTY662r/+JXjF/mBCck/LthMZW2QW
8vhCNP6zhMbHAZ+6z0R9hIGaLTtKiddYp6fjDA4lPiMIPG7SjXLdB4Gj18p5jqru3s20x84tQvpE
EX6+rXjdgab/9OmLSQIO0GUJwYOcBNyGyUdQ7Hgvfnn0R8ABWWw0tKlPmdxf26IPrsW2j6ZARX9A
bEWBRsDDnqWDyYsonSxRjDuZx75lSjCz9H59USmEERw2SmuB3NDI9ihSO1M6Y+sgs5VmczLgb+9w
kIM7FzOex+iZ1bjJQGdakFZ6g9UbdjQ6gUfS/H08cENLIUvBvET4WkbybTAds3fJOYJQ0GUuKWuO
/hE6ff+tpdogMStzv8y/3STj4v4dxWkbb9euDxLuCEperJ5362DGsDRZCrBK9TGBhF9uUY+3MXVJ
l/66w2Jj7IMVY/txsaRT6vC53ejPiSphRRXqcEoQVMzN8rKTJmYqWEvENj1ncSyStRGG4fnvF2SR
F+fqlon0OgZM707aQdkjK5Q4kfapV9w8t84xHeFXTP1FvQKDrxodWwKWOJhIEuDRs+PlHdEubXJG
jwJgydAJxPEDsHwEqM/wvJ65ua8Ldgmb4FpzcI/wlODs7hYXRtoIgOb/F4a/UN1pfZtrg84QnaeL
xsDXEF0mZF2zLqwg1UTGr4JGVdb7ED+i4IiDFEW+B3lW/dzkoAKR/7AmVw+DhjhUtUOGqBCdGkVb
ubPVPTbpD1OoOpR0SMFWpbJFr/3Pb5+S+duCXZCGUwYDnPCAeyLPwIa6h37hlaPR0R3IWvO2pBs0
uScRf3+pWunzjOIvUA16teDa2moLreuytDto8nPzXsxoFB3HIy3wTsp+40ZcTYce+KijxrFGsCvT
O5g3wdiGLEPilCU1th5E/1hOTaXeYEf54n+JbTqzgB4OVTSh9FWLUgeGvHx7/X1JtgNCTh5x0+z3
ssgzhL5nhQHlnEBTR+O4B9NAsI3/hIr6ca2u0oujrmFF2yIFBrJvVojxu+mn6cQj3qNIlr9W+G5s
Lrx4gYfo6WE2z7VmBCo797nTChNZ+yn1SVq5NVk582N48Li22OYExciofmQKA8N3vpqgDjllzaWM
2w79aCvzljA8JrZp1MeaUf+bgJbjNHxARTgebIcg96/12nJrFdiTmRj2jPU38IYMRGF//wz4KrsD
q2Kei6n9TsnZitOjA35aLKWH8nZ4j8L1cHFuHGn5SiM21YKYBT7fGB2myBngpDTY3y6rd1nZikIg
G7K7QEKc51F2PSAktZniLcfA1VYVs21/1ydUN89AORYoOUvqWG/Pg/TmQxHuktlulHU1iC+Tdlb+
kF7xU65zRK5Zk/W5G1edHsVdGevKX0GBxI+IwrXzIAU6ddFJTdduZOasz/e+fHUf4gE3YZksqSZJ
AbzBdEGpmLfJkLS6+GaSm+GGv+UsPHE1pw4g/9Y6XBgMIUsWKpc+rTe/cSDg00bcdZtAd1SUgcD1
E3QbU1VfYBMNT21Ykh/3mfue/lGQWByOgPA3S95Nv68Y143uATHi4grDJ8Rj7i9C7W/obtuxYNP4
P67Pt64PKkJFmSGRn9eeIxyFs1xSDxHkHXNUmPcB8LLYOrl+XMD+spK1xTWaXf5NpAwDsqDmMgrb
GBNZ1vt7IML/57L8tvxbJyOixpQ8gfhLM//eQkD1yig8s7PxPJ8rTY9Jx/KD7mdXCmH4YhHyYnA7
aaaSkvqZbiY9JSjx0CGgKDdK4pLdkUNVdACkhWxfPulvE207GsegQ8+Zshw/LFPsj2FMEJAawemi
aiOTsAlMeUCiV43NPwqAucK/cFkRCQ/qMadOJRW50X6+ToMZLW+RsdiFCgTvBWaAWfP/LM7rjhsG
lZNoxg7SZPQCUniNFZjitd0c2nuL6OQ6p/RqPi3ZJxBEzemgF5BoMmLjN3V1bhfreCZ2SY1t1vsB
9kEEksxlgnGZcoLAFuTw/+H8+Qued3Jf1HefMzpk+fuw4jbMgsVnqZQWp8hfQ6iYz13kgmTer9Uj
Ang+UlOYgSLVZVerq8ASt6szlo0STLKME8NouVgb9bRn8Fg1NU07nYJ87EN5xMnJIIF/GgeSo3+v
3HpCrXs6cvgQ/MfbFrl9GqNJ0DArd0EguGnO/9vZUUcdob6QF0tQSF5JSJ+OPhiKYxlEHk9YnEac
Zqe7gjz1cvBAHe7yK+5KqvxCoAFCqv/vXddGZW+aR8lkBI6hXRn9hCsCo70xJt2sjZuF4+RAyLZH
DLNhI2+jTjqnHIdWyxGTYdPo0Wv83mko59lt/c7b1269Z+B6bC1r5k5WRi2PCPx15aq5QuNUNhNq
5xQHfy20/V/yEJNC1QkHw/cBjq6sepg6d2s5DjBS8QOcu1m6Sxlt/5enVouBaAx8JkNFElhjHAOR
hcxB9jciXrAB8rByNrH04MS1cXkTYdDbI1zGuT3SaM6UT+2hrpbZ1QysIJXHCVsCkkw3efueue0L
J3tBlH1LISxbcnVFeOsh01Pp4pdFPdoaHc9xfHUgS8/G4cZAYjOnF94X+oFqS3HOBU+OEQWHjyyW
QFtoKvW+cIVPJqVvJmwxxFyPlCAkLbBXs/m+5hU7gSKp5HRrbLGLUPY9Mh7zntV+n5nB20qIliDq
uqcmxgu/67THHQfayjpvfFLrXkEebqxHSuxY/m9K4RnJodBViWG3TTRJ2guP2+lGe42yra3MFMER
2s3kVzPd9VitmOeA720A9NI+J3+AgXsDO080j+7BQ7q90sLw/mmzGWUuFKmCi6gs4ssrkOTLyZK6
NJssZ9lXSfXeHnRnTCqGs/OwU+UAVtJsFaJc9ot1FhWKinU9Ocrks5xYToEMopKNHZw26t17zYoZ
hVmXhZk8rrF18z1vpbzMdzY5bRWtmDf14bnzJVX9DkcL+BmuVxMO4r/6+PtMAPVBFd7ivyo9BLej
K7wWoK+JNCAGPZFHl5EZFZwmEbQruYYwEN9fOituLb1LWBJZ1HasmZGrDAd6DS3U1QuVjPdgy53P
Pjkenmn6AafzNH6hNEdYaf526diuQbet9hAFJLVJgolp83HSHVImqQ9UMvzCr0KiJwjWINBw3KO8
ZGVjbQudtpSYtCc8j5tkmSiHK1rJsnHpwjwXkPbRNs7M7PbRVxhZc++ncLw8xQ5R9lzaUSzQaNzj
K0+rL2qM5OkD00KikcfXoBaiNF/jYiCc6qpuA7tlF8tNvKf7nDAILnDVwM4iCVy1VPr5HbIHJ0j+
ahd6sU243cle4zDtIqZRkV5Ssij346Xs4MBoOHI2RZfPrTkLgMzl5m7D7WPJXS5iPgnP2PGsv7Ug
nJof0lq0T96WUci2Kl+FtdqkpkQ2+RAXXkY1u7OkEJkY06pVHkcOUEDfzCtxIWLg02RP7X4KmC+J
5x5SSb9xeR06I8de3qxUAVzLl4iMqFpv7JxqvptHvwX3YymACHjoLkLvumqBUKmkD7sWNyH7BaWH
+er+6iaXKqjH4Gq9kh1CgmQOGtzOR4XqTEf7uBefDwwQd9sK4rdm42wx1XS2DEe/fuVswdxklBsf
dsss+P5TxERSP65ATjvYoncx9oXhZR40QovMlpOOPnFexg3ix0njNB5YTMKJ+F3nZdCNXqGy1w76
CxsfmQnUp9HVNZ/1uzWwnBEypuLgSC7mSRQJcKx7cp9oPtq10GNrr/QxStBX4KgHtkoj8mSOXi+M
4aHaARlmxBiTyFszOG1FVgMcd3wIZU+MxvHBEPNX8vcQl5QXfk0canoSYq6f2jOqFZDX6RLJYns9
49Tjo7zg263D0PK6m2LqOQeRrg61LYc7rc45Yltoif6FLaAacTC1JeFOWC1PNjpPSftSUaRa8Blq
CAtJGsK0b1DcBEbijCpkFyw4At9LEjQMOiVRSqdRr+M1DOuBL0trstSX5aBdLDE/L2YAmqN04hnC
GL+koQJ746Q3oL9mQUNQZMU0TvY8zxEnDyvngHzX/yf1rJ0KQWls0LiyLGIXbmI1Oxlu2/wdzzpV
QjoQ+KpA5fPg2M6OuvcYcpsEZafwx35F2Pvh4Dn8rF6n15ECuDr0uC7Ffguwjdm7Bpw6ThS3OnJb
a8VS0Dm44iq02TyuG1E3KhH+Dl4F75GZh67pgajQrEdA1xt2o0CbPRbR/Up7qT1vNOfPd0Wm0nDs
m2l+5PbJc0Kgkihiy/T8ujNyeIkx0PlqVz9XYMKe1MLnw0BAXpphqgXohK7dzW3VQk7SuYsJT23t
FuzSVubGyAQbljswXmsDtMtG4+Dvp1vfv0On0fwSFGroFgdD2ws21N9QA6sJon7DZcF9W2ObgfgR
YWyoVU2Ia5BuXtEGMwxM9rHbaPd/OIfaqa4Eqq4iQoLSqCP/URvZL7RSK6l0Y56JpHyuEJ/iJo1I
yIrjHu56uQ15RGMS1Y8ztEiZbuvhKqRJqDdVM5lHtWV7o9RuoQR+GePJmtmT1YaW5zcNqlg6Jz3d
GF0BCEZuWiZgUwsT4+qjKct3XYvSn5VBzk2dHmJ8Hkb02I8vwHpcpKK6wKL1McA3LnUza1LoscIy
JiD8k4A0KEu5gev5N1dwPuxfHwYdAGfz/rPrOjWghKvuJjoDCsNaj4FlVrczbWfulpp1Dp5g3+iq
MFr+54A6zM987QgteAT9GwONA/DQT8IWJTT+Q/irHMWuB/KFNWXkrA/P2QXebFwOBQUw/EUrVXBp
QTCx2arO+16UYpKRxmsEVtHSo1cSmOtf8pGAWhD2Ms9Jrwv5aDgXVqvm6EufkBVsnErCcmGJbpz8
8iQj1W4JGdWCDaC3H+DVyRt9L6E7m9Myv+h2DveqqE2gQt+RVPW+Sg/XuMrJ3DVqTrG9O8xBJitu
k70MqozFKuktD2oKo0dhWdPI0G5te3pFzHYNq39mQIkhxuSpsEm8Ip0ZVX9PD3dAE1uy1c17J+97
7yAAqLsEijv9t9FCvidekcCp8L1QxllGIICBiXTMTvQpTaiS8rbneD0w8UlxBD/Uikpn+IA5I34H
F6RAzwnFP46kNtAGCNDqm0bmDx1ScZaTtslYN9NBf1sRWW0wOdEg6yhL2qG0uSyQabckj/Qflqf3
6NXEO6o8xU9epGULXJIGDYfWbLD3/D5BWGJsYB/cuV3vqbgrMLzjJ50jjQVL2713lxLowcBg4NzA
Bk9CTELLKJ/u6MJGJaCJ9onOR2q9O4R2WcHpqLtwKOFWB4hoXLVzQe2ewbCJgJKfwudXVCsPfUf8
FnpGmeH40xw8H7NeaQmptAcxzK9ojlPq9trGamDZK0C762vWA4x3zeWfM41hiz0siY7j9u+hozOo
Kk+MUBbJVF5pgnM6/hvk/nQIb98YL/xG02D3mtG9h0UuEH0uCXDS1VfIHP4VHpgS6o+EuBR7oILM
YL4eDA0vE48ZxHdomrKyi0Nmt+hgX1T/J3nRaVbAKwX8VKEliZx49iFwsFMx9q1A38z92C2g1Pd4
7Po2+cIZB2TTF7oWmQclpd1bKymnLNjurOtA6bmA9R6Z0hGfhQoYvq0U3bbOF9+RcZh+8SlpnIvd
y1MUch6fDkCwpzsk/ZH6gYc4tczwyhDmHVja+87f2yWlnHFRgbiuB4OL/D+GWo2nW8DGM2mytzZI
8fhEAcX6juQIVgjmQVhCc5NWaKmOlRuI+F23wJZh/HyPGLnVFrR3Go905kIWDtHMrBrC47jK/dMg
zCdTUfFlp61i9wctlOqAJoFbyJ7h0YfMbzaRswSq/HAQPbQ6Wo1slIbNz2/D4ZdvrXloSu+9wfQD
AJr1gVombbzr9wt4VRSwclCgzL63saL8qKVNDlF6desCs2aFvp/Mq3YXIgenTj2RJBX1jL1YfU+x
8Nj8nT2vhfdCa8K4E5UIwnt/28DQdLT33IAEwtbNKD7ha2mzqCVCghtBYmswTkji7ZV45tfS5Qm9
wM3zNx4rTHtDboQFbHxCCbrNC4DcOUyOti0C8ScuKq6WOeddVLNs5vMfE0mnrI84k5YNIsJ6mLLf
Ln2OXlZCzAInMoZU0uudiBEN1Fin7is60ZNJsQ/QCQx8wZRXHRMIfZqpSaW2ohWcakBxoOrp50mA
8NlZqrlfK+FnaZvNz6Vlbaane9fkp1Jj88NR45qi/ebBtWmG5fAcuYqAr3/I+0vK7l0EGmSUrZnW
OwlYclCxckzbgWW1BvHAFIaa+/YgeSGDLpD9J9vql7KtPtkRGoq/yQZ9N/HeyOwwIQ3PhZVAzYIu
LGRYIrsqRknvvTXpEl+uroKQFfdc8rPtxUlSho0iPkHZJaPVoZMIw/x3qacwCVdkCXjW042cNeJo
o0su88HSj2SAkiC+7QzvUxSNnmw3AfvvTlp7gpvGHV76X+scA5J8cSxMGE8r21leXJX5Icu3X8Hf
HLDfWlOywDHQJ04tqAVa/75k3orJkbUZwsgIB0ZlxC//z4m+tB0fGLJfBYwWe6LM5gU8ic21Wyxa
K4yOF9gIInHv+WKIMYf6UcrDPMce46tiiJc/mM9gExpB/58sCZKKOpVxPxxaUKdna0xalYMSXKAL
htKSuukdSssRh9c8Z5EzmYMqsWeBQTKDdQH6408IJQbYbTXXQ9OeyCxfO4C6PwSuf+qMATNQNUfc
3hEYwCOqZeU1OICPe0pKcY+3EGH3OiZAES4hLWxOHJyEqzKdS4Ord0MO69+tNQq7uQ4uWG7HnRpO
lRkAUDyrS+rbIjIPslEv447Od7DJgaS3qAEpqPXoV7Oz1hMQsvsRGg6bCLOESype9BSiyd90LyMM
+9irzYwubH5EwI3DGZhi/aII7paQd4WZ/oVfZqIC1rCI4XBPnr6RYN/9fYV1s/nWq8GUhS5Xq/BB
DX4cPPgq98Bd5gzK8aMiC+cGQ2+QHH+pJ98qivGvG3FiHQ2SBCzu0vhaLpxZnuj+sisZuCOTveij
6bLXzOiSOmX3rVKEegJIXEuzKks0FdfkjQWJph0UFJHO+BraM/HhOddb4kiZ8a5cA8cYqhjytluL
XXglN2PYs+xjM5AljBjF5m74JlVCB9B3h+kWc06S7X+sZCXlZgyUAb47s3fSMVZwHmTZ5/Vitfbx
WzvzPNeFrS+LzBBeR3wrjLUItvFOaBEmlZx+MX7HJ8ynRI0/NCvvEsYA2KcYh3nJKE/RZmsR7z4W
sAY23Ro/HTsh0NBo19VMtDJNVeUVLDYlwkWOq9mfjLbMfhJHum2m8b6MCgGtEpRDEq4UAPOIKe7x
8DPWbfp5PeU30csnNd3KnOFZAwzQ4iqMjjrZK8+XssJgv163E6HAR8QHk1hnjHivpwBQXhtuAE7r
3pSpPfrTpev7zb4jI1Ow8SImQ3FKPhqf89GBqTr6yHInFv/fhV8yM40Rb7/UUPLI/5kO7JqPA681
XMFVr5V1QRqHwUHVejCXRhIpQTxBwdmbIn2mb3vZ+dYBLrQAWXDtRClWhcpo2S3bSEvCx9nAziZF
y12CSkeCKfoi1zqDqgqwAOcllSw2P6AwrfkO/XKTfc9Hf9TLjuvshZM8dyRzvSP1if0DPyzNE/yr
lw4t1kei1PsQ0TKIumfmmmytsooYMMWfzeDrTveOghgkdHCjtSR09DBtxUpgJ29FyUMYwWxSW2I1
PLKwGhPAs3k+bmq9z1NRQ1CD/tR4qCsxbZSq/qFtYr1+bQwIqXIvIgjZJm/SbnUtwyHdhQPXWJ7d
wyTD7TPMwwrgtWzhg/lybghA3pfbPnUsFPP5ZJInck8PM8b368YFWsb7/tlmyFuU09BUqoRpLlQl
dwATvu3RD1TKtImkGm735cmItiB8+TxeloQW/nBMiinbo6nZPxW1Ybui3BwDkMUzDOGjYGJC3C4K
fs66Nz0KmZVcIeon3Qs2JlszMrSBHMh/L+taVxf0J7BEnRF8oq0modrToHhIQCTwJrTH9v4w2Jyd
52WUQ/PI/ThCLt+RdctGkOIGkzF79x4XHYCq4QFABS40ZpWB3mofUvR1tBTDpAryYuEeQfGEdnOu
IW8xiZb+wMx0YvBs5TCbQHf5b65tn1bhkXnf4o2hLK8hXiogfHXWpmna8ViABTh0uO4UHoxi0Vx2
qFrAkhaU5HLR03W5Gi62E6bKjGNUha4+yf8s32NA7Pgrzx0KrMhCem6wMAJMc3IDng+gwWYpAPNW
1P9mPjPlPK3u+yC7uvdW7SDgIIDDacPFqhaJOGz+4B95MA1FVXwUpbE+yypLXtpUFhQPebVhhZBc
5uXt4MArok55VXEKH+Uul41xqYAj/4epv4zy7o9gc8YbCgJPKfpJckCvaWQq74RfkjqDXnIgOo2t
YbuvS/gvNMcKtbEp1UPBtUPw95z35MjHrSrjOmXZQilgVZhI07c1olvK6kEbEXlPs4Sryzd2I4MG
aHASHVYoBPdu66BEYxpCPY01TPg9LPyiOzT2sUr+1dvvjVGGl17poXg0bTd9ekLKBSyTGHAV5tm4
qFfK9irJDSem7j0hXhRezU+4U0Hnh/WOHRXTMB6sSyzhIV4BJveCJ2l9OVJYBqfRsnsTrSjAh0I1
PMcLpXCFHyRl9pL8tilYX3JBBtkbRBfHpqQ6zyZXO2QItjkdtu/i5aRI1rp00Jq1WT6vX3Z9wQEP
gs2fW6FSKRuuaiK6jFhuDjhN9MzR8sp/XJOydSzZBNcGFp2oHPGkdvPBzdKqyneydGdEpN0G58yF
9C1MqMm+fkwARqcjPy0nHoMDiV96RPakmcGqYagYXwnWc/+BJz4BAeOGr6XBc3ovjjyB1OKsslzB
t9VB4bIAecTItlQHLOsex759t4deW+96X87YFYOdLCDVOPC9sy4b5GP/VncbrdNJl9zTLF5JP781
rhlqPeZUl420e0ChFGKzKRLNP0NkWOHyvPHrG4T08tSXL+5ZrVCvkPTgne9pvFU3YzklldeHa364
oqASIohvnj1bgqICSqGFakV9kSIVQY2szkC/sAW3pmj5zWOQkWULDmEGVYqFsIYM8wfBLP9plUcT
D06cNHpNKVYKlxkbcB/w1y+0yE2Py4jXow4ikXr5yM0CO+WFI6M0ZYir4STSVMoA66CeX+Bq4OxV
g1KjwOydJn4sXPrvbvoEeN/vZMwlpVUb9vT7T5s6rmcwuqU1gwABbqtz/fp+p2gFeAdRYb3MU66y
m8GfxFyeVcKKugRNlXsnp5XC2rDESLSsDmCe5GPuQWOCjT1OayLF4/8xCcYFXrWyZrbPLJqUJ73h
gN6HwNid1/Om4m3cpDlvxHpdqZazy3WH4dmpgOSGM9/Jvf0kWS9BsHplQVgkZjnLq/B1+inuoqGO
846Ub85Bw/0nHXQBJyi7RKJ8gmRbX/nYMA4dGQo5WnArh4NLUdgavcAY5rlNI+gJ0fPiSp5qrQwJ
X817jUPhOj2n80pyRzz3FdIRkKQhYbGHKNIH5BUh7bjeZ9NKw5AFM8Qkbn7Yyl0MMOIan1GZklNU
7a7KciIGRwQ98DCK4Tk0O5CFC+c7KAapZbMNufFBJ7QVWOz70n9PlFpAe3ImuJlcbXYj73PPtl23
qA12JqnPYJ7T0/hCJy0y736FIKAF+SLKWHiZWBzP0EzCMJkyNwXdNvfH+yYo8sv95nij+cSMzFZl
clzemxWkF4pti2VN451E20Rwsssxv9TDs4ENCQGT0WvIxWtF0I6qC4ZrsZ51t3i8L/7sqptvEVle
ld7x2IloxSa6CyhySLt/T6jK2u9jwIuWGkags3sC8PeIs3SnjGSU/iL/mHEluDZLLpB2AB4U9Znx
5pm5hg5dq3X5lvvJtzwfzNgD7NWRrwugyZKR0Dca+vrutns/6cKduhFhefW7qzB9GhLGv6gE2N7A
Ln9VIxb9EsCec5OOOtpLwKQPXoY7foqu2y447IL+4N36yBwWsBCwgaX7mDpOmYZklKK4TZihslt4
Ucw18T/DngNhycDm3W3B8gz1RA/ADGR73LS2oB7IncjepoztH7lUHgj+Acv5w5dXv7ocbUqgestO
hiJsAaWIuUPNYjxi2XVp2k4/qr2ATsbgG8VmClGW174Ek2UeqeLTq47Pyimg661QWYzLDyHkOO2I
PW6i7rxBnuv0Sb1caPgd7Is+S1tvlwoq2Bo0xtZnoLwrqNdZ4y9ypinwtjs3XB61vONhqh1K6uMm
Ss6Uh3A2jkUfdsD8OaH3ECMo0nx1d5xEAEP82wT5mtFbOc9b+7s3fXrwkqRNzIbRRzYyqCkLlssr
K8JDRRJ+T+9cV03LC2HkxUHZo2LNBhHr/FGVVm4xHpieuzQqt9HlZpZmybVaNp3JQVxJ+HZqqDf6
wCUAwdk0EYg8E+ImjmlNGa6QW4k+jEpcjJ79uK/e+zsravCBMG9jA4TSDEiR9FPbDxMehky0Gdpt
8vEgLW8IVCI3GPkhuGw9WmGulIMPmsSYj+XO1NeD5ikt24Sb1NJnF4AauSboaLxjO6ihRXf3q9i/
qdBctZuwyJoAPGb6Fjjs40vwRRPUontYapUE814jG9s/B1Jm+5f3B/Sn8sTnml3Jvtb9V7F6Or4j
g56lJSYwTK8FhPLOab5UL+vqwQn3j++f9B9RgAZwskkqB2JIY2UMs/ykGi7mrULG6aXIcCK06YAo
LD2s71G+iFgNAo8hhPmg4UZXq/7txHO3jGNkX0MOUGMccLkSXosKxd+ANDEw/XFVUZDr7iHE8maK
011LpU6rQ6YmjHGk5UFa6OGncIOAohIcuvSscIHof20Jv/GRmlYTM1Uul8odls7/HErt6E8/J6gI
Wb7EspkKXXV6MEywu0dQdf+WL5bpgW/V0bR0eUIAjL22QrolPfdXoqb+IBI4Zimjx4sffrztywEv
lbIeCigbKxap+oqtlEurIdjY5DDXfZFAUQQjIZjv9bkgKRlXqRiiFKByEfqBObhlk4Bsxn27+Yzs
9OAOXhE0vr3DM7A6+N22MF33hXR5gCGvk+qwsHegUN4125ZM1j2iOuTe+yNbAC9RHSJjNwAZ4TBH
FE4WB/eECNcop3h0kCvgWXFrmp4AjQrBrU3BvSkDoiGYFYrKb/u0qcUhho4qqIWkePdAjnSPwR8/
CNFo6nYeJqCfVK9j10biDRzS7cezZq/OddF/CFWHpJUGLadofi3zePAGywEo9vWr0eQiqFyTLWsz
SJl1YGES5d7fMuxmKJX+WJ0drCWYTET7QLukK3cHPYW9v59obsRGFUFXbQMJEa4tfAqQEFS9vKlC
bjNfze1tlSucxUo/xcRxNrXkYcuBrw/QqKxX1qVDPPKdFrxsp/ek20UuK8fQn353Z7kkYToa4zHl
q4y3hUHYYHGJxtjU3VW8YjB42LHqO+Ao1VRnJDAV0PQAnzJx6/VR3H+8DhVEMJKTCJ66HN+ukUXZ
pujnMCZm7GM0HiWW49AzQ7LdbrO8aqcJR4hZbE609DQoAo6moeq5vHTP8adLOKltoawVAZXybdLa
ui8SaIcG5agn7kCeEtjSd6lGMbwRzJGZnzpyHdQ3lf2xQ8+Rvkp4000OGVI8FjNMBoAZyFpWw0Kb
hCfANEzSojoUsDov4PU/PYGSceIjV7+AiUWlnydMj1Ko4hpZ2Dxy73pRBK/DbY/mGa9QOBDaejUs
2JCV7qF2RTQEWapLc6AtqMkR+EJNiXSJXCopGuOC/FoG1avxPDnFMYN5GYg9JglZeaEXqj6HsjNF
H/x1RvmXEqpG1wO0smCnEm3tV4z3c0rzegc+6cBIrL+ybdOOBGQtR9K5srVwEZkoefVOzt47hzyq
B7R0S6Pj4BERvD+wUMUVh2dqeQPmcSBY4gHt6YE2Y83x7nd70qlDN8hpkOY09Jww14h4spKyyIbr
4ETYHNS8Tuyh4GSUDI3wuTTNl3WDfSZ326c/r0Cxgr9Db0sUucoYD7HAqpE3GCPMbs7Tto6eVL96
WD0MQAFW4WweTyfzcSQDLckBfImP1aS7hj8HhtGugXi5PFboYZSPYXe84H/88OhQkC6jbhbz0+wN
dJOOyQK9WP7wiqxdsdZnR8biahb45x3CwDaDKGcta2Jqpi2fpNXtu9da1le8ltxqiHMYKjown1zd
GJ1kX8uMwwrloK3GHsj3pCeQ+cTvFpKfM1t8Chv+qyB49se+KTi2BOrYN2oxVgeefOEcu6i84dyU
RuG782O/c84IWknb4HL/UTUZWdbNPlQzadmmyhAi4lha4f/I1BwSYIz9Yr0MyojmtYLcnH+G9apG
YtAMYcwoV5046Fz8lx6eZq7nXfbtdS5fZ3rel11YFPkP5jLUhtJ2YQHmWTxUCJwySAmY/NxeyAPz
4ppEHikjACWL33cA18jVxLjzAeEKbdnYz2g/wDStwIZ3wFddAqSQsqqKU5l117c4VDkZDB0x8Kx+
AkSTf9wCnwBFSiPGonSoXFPt5ENxgCZPTZo405yQ5hs3fZeazsM9LEzo3Bk7dZeXa0k9d3gucrpt
xlseHjaMxKkx42ahQrcuePM5RmrWLr0XJwv4FUwJ5pbZ5HfniH/SUPHhR5WEeZH63n5F5EiXrzAX
kngt35JIAT2gn3kzidAeMVVhECnT/oVQEZDYAXtSuS8PRU/8A7vcUqMADlUTp/wVSbQxya8jjHQl
2pQ1cBdaAkHU0etEg1pDFW1t1vsCSinpwMxUiXxStdXcflXL0wAvv1SBNO1QX2LFDfqfxWN0kJqx
MaFJdH73JM3Nxfx8MPj3QeKBEqi20vvw+Mo91YCfqNxaF8F/XZUCW6yLf9/6JxF5u7GPUZ0ohFxb
T2im5UA6j0F+MR/U15KGnuq4JUhbUxhYLS19jcmkeh269yBUL+tFVTDGH32MHPmY9ZSie40Bv8At
SebzjRtpgTGDbJfl5L/VF5BJ/ceMnxKP6aTqXzz/PrHdPfIx1pyjyFHVtDN8Hrb7VyGWMmNFTIIK
QuuQEzdWwQjegS6N2ceD05N458I3lDfZ3/GpQ+S8e8WFzpr8RiM4KOOpPn5GSOYupkqs8UMhO0Tf
RrAT95zXcxhfbSaY5rZg5B0Th7qTy8nQncqFLjg3IuWpKCFflYWe8fUqD4Wi3LpDISaMEuHO81Hu
P49/VnQCh+x+pRnBt93wn3ZRCamIe1vbyrsENZWT/8wwIgPslkZYMdnOh6PndxpdR1FQjjPpQfNf
CB4/rF1sQN/S5jjvXlz4p2S2R5tXHxhEjBQLxax5KIyo3NiCC08tvZg1alASFv5QJkTSb9yWWoQt
9AQHQt3JtcOqTLGyLpH4Vy4TUKiL19U5l7fUXeocWOvdxoimVF6IFdZJt42w+OkHhHfrK7J0tnLO
7fTVRa0ak322oXCfYx1cph3i+vd8ogeR7HiTEVdxHESgXStabwCB8n6vvPlC5ZUaO84g4Soa7Us/
z94UZc4Ln0kgvEgQrJJZT8M3l67my24xDh7xHu0j22E9O2MWoXH0IPWjZJWQ5Qe2eFhMOlo7LwpK
OPNc1Bnzlh6GIbWfuJyZnY5qPx2mK/6a3zmWtAuC2KCtKuZNYPRjgG+r06qbvOKz82ihxMWJuomY
aBx4YfanwKeuwqHoRRQ6I0xN51y5kV0hXZV6ugxlbiSbSO0yx0p9VcB7zkAwpDdWHySOK6b5H2dh
m/DqUwbf1Jkkxwuh2vNJRa3GqCkSM3x0U/TNCN2GfEc0/yfKrelHaJUPUZ2dds04coSGIw3nyAim
bVcNshneOwRhwUR1snvOtqghcBIPf2bVJPWqDYQy7y9gJ5D0Ru11l626sqo4Aytswpw5u3NvN/TT
OVydOCAhPI7eS7wLB3IQKDbuZlqED/vSyOuXLkxO02jUcVCv4JtSdaJzDctzSbusDfEUncjETs4R
IfQxDJMLpyOyfX0O/vbiwBB3NQjK/GaRSR5+bFONb1QeqV5dTlQOHJixMQfhvbv6cFSXTnDK9wc9
h/75DR/mQuxjXdbEO/Z/aHF3aKSgIWuC7P9IAXQg9XqU25WL7q2JUvvYJ+Pk6bLl13W3WNMMEnMV
nhFbkAAu3ccrAmNeJMtcVFMy/XANP3PM4XZsetjcETpgubbxWH/e8cksRC/kubz82GoedR9mgov4
bMboDVrojWOCJ9MywZvtVwJUFdlFraOSulzx5O//NBZolEB4QX3q/Gg9XN9/vQQLqmxjtQw//48e
9FnKtJE91NSLIilDFYdY1SRjZ30OXhY2GHh43YyhRDn+YAuiohkPufaNIl/uX4Bqs6IzyIRKfAI0
VIFzDMGM9gnLtlkpJ8N3FC+dURQQxaWNQGbix4OQH3LDlr0FX76zf35DmZcDoJCE5TY/mSatOrxm
vhBhxcpThrkDCvPGrAGx6PYBhNdK5Z1g3uuakFuKOYPi4Ile4NAOLKQsakpwjrkCTU7gKf/VNAC9
tk8xfAjv1uds7fURkKh7ZOVEva95Jds4G3VEz6dYOg8uhGEZ4w/61Sxsllsnuwp7FlHD/EtjIYYV
C70BFd9JH834lwv9ugaKuRKBkKGLuzZ57iuzyZD/sN61x8zAJPgwHYIz5x5kjwvE4zVIjDL7cWdW
E0cDAfHcNGOStcSE6u1Dd3vnyud8A+30K8IR7Xq8BL9kePKeY7zAqdWybeY+cpfoD+gvaUwgiqK6
PST4WxsP0jHjkwdoUAIpUSqEVwpCQaRxTG1UnF8TJotwoEWTY9eAtVjbeiHLlOoWCsuHQkhb0UhH
vn5j8aIbESXXztQ/ofr8D4hY72I5u0ibvYbYoC5vhkqg07B+rOWAJUC2oQAF3Do88NrpxKE/1dan
qneBESIeX1nNm+Zob5BnLQeqTd3W1L9tJM5SgaKXdd61S6E8uNFWnjhqPF+SfqDoL4I5Sdu6Pepz
ZHlDD2+dTSYLNVNElrHDy5lPOxy4Ob+A8tzoe939P/x0ET11V/iM36it3gtRTfzh+TqU8WmeL6MP
3BxiJKDWAaevuxMD6SV5f/TkI/bJlFmgMU/5PerCn7EzwbhNWnlhokNM6Ua4mzSf8FKkLF3BgO0Z
sL0N7lypa+3QuIhkaFXglWrGs4pRZeqXz8blmXAVhb4rNasRn5Tv4M9P5CA9AfRkqONG08yNftlF
ys8vRNH93mZb6GRqZSrz2j+BrF46PZ16jLl8+VYV5C3a+mqI8oB9KV3yPrpgepvvUkquWypxNeAC
mr/+Rl8/IT8F6lPYj1eSwh5UeGvpPq7KdChSbEmkomZvIS5VbTcEruOxgcJ5/m+7PDD8OfqAKVFN
0782ztkGMxUE9035puctlI9sRWmqLQObXyV/GIjgezslFnX52C/YVWVwHmUgSj0YoIB+QkmRlE8o
LLdHs9kdc+3L00gJQvSNkOpe+gWXZZYIhmuAubipaWP2uv8cCs7KZkQBoPJ52a0FcUG435Xdh5Ll
1pBRKf5+dxDsBDJSPMOQ3tfLcb9ygEJepGxlgaewNJHeIMUTSE64MQuSAd2HOCrxa8DJsmaZeCFV
chrPliDvq1g7V5v+rctDCZzjVNzOIW6xVIfw7swE844TND6ykuwCNTUaXkazWkIQ5xVHCwW3zc3/
ZhMyuhfwmEFrUZtuV0HcKAyvSLk/n813gcLpG3qaTbv1mSjsFjAUUn9iAwZNSW0oaPOos/ZDf7dj
NqzWDeS1G4qBP5Wr8pbADhYZewihofqY2uUxG7lY3wimoq+moFtNowSIMzGYfEa1BHtEBXI7buRz
SCjLicUp6fBKAoAHCn5j66PrWK36yuhDlN4fGRe14ft5P36i/liFaFKt792ar9+e0bv/A5R110KM
t0Pqh7qhYG8UKADL4GKEDuuXT7WfymMvCWsMMdew03ADXcQUxgUxKO+MTabikU6TwNeVSmI3CJX6
ZsCkO0G6skGZx/Fbk3UvYD7QvBjg8a7+VGec47oUEISKquEbQUpMwxM1Qsfc2kAQgmqS8wzBG1pi
FPw8QMdcrSO7uJcNweFVkn7A3nIF8QziIlZwXkxeqP/Fn/1vcPNhKgtjuykr9HPawSA2ruXWYdUR
mpQxzqGODWjF8sRYQFX1N0cd61je1b73Cr9agqdNhxK/T5e1sUwqX6La1ZeFQk/BP1zmsG3NVNj4
ynxQu99ZYNf1imcCj5QIL1n2VeoeSLdTVc6oqozD2noN0lOwdWEI54DsIGaoKbSgFQtsmINQbHcw
TrGx/hHQEn/YuNfw2xhfmptx+aeT2igR4ErSu21/o4L6cikGhbgd1vC6JDC2TZu5O48yc34CE1sM
iBTh92CEO/8fP8wXfEbUwxhj3zG3gxuDGxHYy6QDgVe8CXZNSvmB+EzM8FaW4PHPfK28h/2yQrvy
+gGNeWYhHNKiDLozxH5Bka6zOeGa3UP9AHjZ9WWCzOY8N4sGrfmD/1d+EoXAAQv0CLp4lHlI7lGh
fpBNl9uzOsZNrBprCzr8QOtlgxFiy6QWsJ9EKw1D7czO1CVnYLn7vcsutk5exSimT0vdn39TRKod
ErGhrHgfVPuL4FJEtWRrlc38wivRFNfajz+f5Ocqyo5AAZ0gc5crkcil0sWN3RePysKMiJ3HA8xU
v/x+KK1/YGS0b+mi/f6kW475htAYFf0YnBkT6MdAv6WreZ27hSmxJD7ByTtosEqKM6RQpcDk1FVC
qt6p1MTLXyktX9koZbjlIhF8tRn/ODugd7/xjTOtIKRY/ljRnqkyD+XOVOhKuBiYwxAtvBfUKb67
YkIl6lpAxbFhqra7JAOmQYsx7eyKW+gFt+MVofbpfL8h/UZJ3bj8W2lgCmYxhg49XNCLc3qdCV+V
YYjsFuNTzm/yP8o+bl3X1uS0PvPFzmwWe1HKBDjl1EAqClyG7JZH3/0aBzY3hC8Yg2ikquaU2aqr
COvCI70CrVZ6cpii98eQbftpR3q+Z4++xers91FC5iXnbjSWjLaBrP36AugThv6oiDtNEOirzx7o
qlvq8FDfud5WUSJmUfhW2DDkfMsc41N6u+1Jqhh/ydHbFe801/9/Zc4ker1Qc3+LE+icoomgCKor
MTT+mfE3RgqqvAn4URjkjyzCmfJv/cD5BWCc1WnaXVixGipTiV/FNSDXDEUXxxCsoHfQOt7m5fau
AJoMglwAagb5PBsAeKDtqkvowERKii6bwt1jlnbqNGbPdcXYBsHo9xs+x6A1aP/t7tFZjeZh4NWD
/bl5m/IkS5xbcLtxiVE9joxpPCnJg4j13I+Dpiu836OxYPNLVfHm6OPh2VD6gNeLDfXxcyD42SiL
X0E+2KUuHGw/LqkdqHKjOt55e4ePLs2Yb74X1RIzXXUeNrTWF2RCIja1t8aCvvc7fBd+WhKQiIwg
HlxCsFIkE0/CV7Xg9yv9Ou9lfoy5P3Cl/p3F4gUgTLUcACY233MYh71mZ1k8UY/ITMXwZA258pcc
DX2G06POepG81QGGKw3W9BOM6HoNNNze83J8+mGs0rdu0W0OlzYMdNo3g9QJJciXscFT9e0dCkj2
A9QVoPqL3BHJ4S0YepfNvQE9O6qt98sjIP81Gtj3E+V/5q87uwt/v1E0QUaZD6V6ET/tJyRN1AjT
LgxqYD9izD6tpti30hgena3fLrgEadY3O/FGsfWHgDG4XvZt6Q9vnSUdrhO2Um8HAEIUc8kMcAio
T0e8FzeKwXMp1C2iyc+emb1OZn9DFAc4VdafW/igOekBT0Ly675gXyevqEBGdId5nCmEqGtKPOt1
03q4SvTIC+5CNgb04qTDaC3rDUTwUEYrtvkLvU2MA2zZFWX5XZXjBTs0SnnkzNEFFLQS3lb1Vyj6
r4DJ8k3U9WH/6L3ObVdNneCtjaiXelS9FWjGPwv4Lxr6D6+2LdWXXbulAlpiG0cvnaa6WzzyzBm/
8mdJbz8IisBEyQVHZe2VWCZ6SPJUreufYiQ0pI9AHIyhSAKK8jY9Mptw3DMtyZbzKjmAGSHSVUIL
LoKOOwIbkVjwF44j4dhJdsPIDvnTG8sNWqZExy20fXTA/jUI2eYoPxmjrQzNvXzPMpT8OmQ5w64w
8xLVDkHima/DRkiJpiBr8ArauPqNd4ayDEAToP+N0cdaQLJd3/+yQvAnuIla1UoRef9QvyHgSV/m
oYEnRwm93oZppHBcM8DCm5Av341OJirDgJ9oUg4q820RP7rDF6SdsZFLaU9EodoM2+IuOl2P390z
tDPp4fCr8ubcw6iUH9luLnxTscViNILAkDXRBBIx9UsWtE0AK4Si3XAvLm40NpPH6xTX4JMtj/0U
eMVLbYkqjVRwTk7lV84bccBC9crWJWe75nVtM2qGILRtAy9Xxp0GIqDm7gCLRDQrOP3VeqcgT5W4
ICv/sd+5GJ+3y4Kd6M49zWt2DB7tOvPdkm9vbhf2fqqNP7ETaIrKYSqFjPCmBK4ADS1o+mAxlltz
daOu9M0AEcB+OHEJICHp/JL5ZbxmkB0wx6m6t5CzkB4Jt5nZfVPBR2jTLJdya1jiw8f5ilDtSUVg
rfvBD06f24b4YHF+/cRE1rJPV0UjnE64MZkd4kb6TKRNyIvDnzVZlUKoDnrbZIXDtdFkun5pTL/I
nz4J5pBofXXQRZOWguZMzM1ekj+7vat6n4scZjhhmLqH68+py9Gd77+jhGGB0PC232zCkd3Od6m7
zpX2Mkhm/+8yD5D01sSYUotkTEYfI4V9JMxC6oCQNUMJ5dGw0tGaNsDEdnQ2a1as8Ts+0rq19Asw
TGAKRigbeBTnnAf6enNhFIgvf6NJfFmUXtzPVFUQLCwcZR0JiLIXPfahRJ/jfgZjhlo9FSLaSkeI
vJT5DQRIxSi4U6C3kDs2Kugr+nFA5/ysf+kt/nr8ZLtL4j2yOSL5PC9Vqj/UmRqeu8tFTl9n7EbP
fKyNYEzSBZEVxVjkygaFydsu4c58zhlzI+b6swzRJf8cyj6ks3xQ/Ir7ETcO/m2g1VCG1Ez9vP7c
4AzHWggr8AsPLbMnEAz1/CmsRupg14Gaz+9gT/f470DRacSj9ysRujz6TRgQvn9RcUXUbqVK8yT3
QqULM4W+Q6mWyEeHgtfGVszkWKVQJ95JT60xtyIy5c57+NFudtAVVT/LNEnJ95RN62Bvke9PWpkz
yP+7wCNFJekBMO6Y2TKr+3E7wjWcz+g1qKcBhzb+A11IAh7mX/XWdbSMQvPKpiUnWMwS5gFwoPgc
qO4tdG/83uFhvOk4xPRtSveG9boluCq0f56UcN+yb7yAalHCgasJapw+mEMC/AjtUKXZx9pqAyM0
HfE3jP5HPO1g0ChPrNMMCTAZjf5dcoatKKrSGhIc2M18ujXLqUqbC9SwClhptShHUD/3AjmQugqD
Qa3OyhIZ8AQJHDB9DF2XjeZPMoXK6GMzj2z/eTwuII+tM9lJSoWtOO5sEfTVeSDOTrtyGSIWBje1
uNCo3xLJLGiderinP94BU03lyIUk+uHUW916PFIjv41k5YYzcbkprKfZtxtS36zgLB7qA0EzAqLT
E9lzTat1EmsPX3WNS9fmBTEdemmwum1ZpOs68UugQ5BoKCjMbHHCQMCrTEUDJXJq7odVfuu4UpHo
nK9D5tHDrf4SOv9IG61g8nkSDTIf+6zUQUI+iKEGk3SSgP6PFNPrsJpv4lktgfeWgmc5ov/7eTe1
d0Y5NN/Bssq/MpaXue8N8COaEYHUjfCO4K2kLKw97w71XIPWA4VRmZSc9D9robMvUJV0oQ/Gqc2B
PlNE0jfJMV++9ZH+fu/YTksWOXsTXTQZZyOhBxZOGZJXZ7hTgxmzP0Np3mG+La4RhJUaOhqqEKsY
eA076B4Hs8+Yjh2h2AxpDUhJlE5YpM+NiaCSIiT5SXa2UeU6/PS5JcG4p3trtd80uqG31G60RLu1
hXnBiNUy6p0ouCx9vO6gXLcexMpZlaY6zjp0mmLJwpZkVhfMNR2BozWjX4pHHwLYHYmBSaG7iPdH
jnib3ORkUXJW+GXuDw5TboAhwPyAZnlhxRbysNaP5xZ8FjCtzdjOrkixuBHrS50umktfL9wRr+5f
XPKWZVFETXlTvbzCvyXB2sGbYNajbAAU2WHWeN73W7hfMsWh5jOM6tX/KqccjGHRUST5hFkNXHxb
MurSHGffLGj5LL+vmXf6ZGrtbjOH0nm6uW+tjdiqNt0d+SoNS1CoJzIpr3SdpHxHUKYRzDOoRX+H
J6fKR9Xaedw/gA7ds6Ta971WuqHOfRRb5W/JudDEtRCAFnch0tbVd7R55BY1Ga48tjT35GCMOSS2
CSqi0srUFt5AwdEfk9Roz/T20m5ns57j6D07DIKTNu59NSPeK1ckdX2EhHFF+2LfQxpgvivWU6r1
Odnu1ZRwwmhaP670ep39zRabtYF8f7TS+3YLlV21SorMIpuw6acDOjWcVo82mhFp5EBy1x6QNG/l
Mbncvajeijd48vvw0bSAlEoClKlsGJIBQAynm3sHqkyyddmoNqOes6nP6YhZF1lu9JwwAsP8YNdJ
3h+iuuVmK3hnrrhmgwinUZfpabtVtDK+tALTqnVPJdcYQK6UKUQcTZrYaJbsxFpwrjgkjRauCgG1
IcY8MTwn0v+AjRgmVJiYs83xB2NtivKFH0dQQVPS49hWVxWquPH4tDqMV2xwzHHmOPuv60OR9iSg
Ag9CUHkRRlTxRQ9RHj7zzR3P+5EtksPWZeOmFGtFmeIPvJt5rkb1H745rNkeJTIcySTJ8+Ero0TP
djLx7DexAydosxwLTWExAB96ft6m08xJxPvrO8yp5tx+tPK0oePwd9Z+qcdjQvhSsKM/c8CZ3ejr
1Xd3xudqpXHwqQuQOhYjkuPQhp5PvlwZ9zPN/8YIKn9TqbvbseRBgC7y51jkECKXEquF8cGdqH5V
aezqxS1S0DiQSaQ89Pf9YmaZUDyb9wWreWE83hgv8MNbZbaxh6nJm2giO+m/ojpnlxbwzGwpHhS2
f1kSG1AY906vGVBcBvogVYXHTDrA6Y1WNqYXkcyGnPOSkl27bWHDzPL6iCm1PHEM+JBKum15Eehi
cnGijVIIWfVt4rSPSOGMj8NCneoeM8UdCx62Fa1DJfn8Uwd3HLxZinh1psNXXUA2bY0niwiCz40i
lClaBg4LXm/sr9Ec37XzbVtkSQ8hS/FlUwQDpZCGtV5zxV65iNr3K4krkY1sUA+6lnnLutUCHcd4
b8eQ9rqkASAz27ofpUO0syEtZDb+nBtxbAq3NUR2LbUaONmzoBblCxUGlJSeIO/803tRys5JnPCs
Wk1sMF+14nszcVh4IRVaVT0UbijRB4629nXYzdoP7F4LtCTNxXjXJxAuoACJZfHzKPUzzb3cxrT2
BbTqRc1RqpIdHiNiKC7LnlpkAw36LUDYewZxIqI+yWS70tK4OX/j6bi2ZpXVHDnKl2+g+3ZCctXa
+wA2Fnc6oq8wOqGUOSEUabdhSYHSM4R47RCCSYPDcgP25zNrdkUvXbiXUVQtEU2BLKKOsxsHu7G0
PQL8VSLbOSqxuScAjFFAvSomoR3WrJoxjahV0KZi+8Q8pE9BkclBkIhZzD/w6ZXgADGtfKtuBoz4
Fh1vkmyxHYkO17dSfvS7tlsSPdrDkz303LtY8JIjVqe0LiT2y9Z184xgGS5adHe90Q97/BmX9saC
MCYb/AvNZnR82Q1L+smR5UFmU1Q2n+mnXWMxfmZKlhoCz7W45UNNZDcwouyx9wdH9JRwEgU801hp
t34vgMu/I/MQppCxgdcTcnkrpJi9R4x8zyed8qw8K9qSSCpNY7/T2iyJwruJ5DB3kyKFP3ltB0oF
PT3kly7KWrsmdT4GimX9sjgNoNzRRlHE+GPxbkzAgNE4oC1rAXq7B+WA0IdiFMrRxB9a76cG5bTF
aFJPj2aliA3LCKq1fDwk/qIK1nfr/NNNjq0vQ75vomIACTSEE3cQxVawZXofFyb6F3ESOt+xx1bE
XwfqCIHosZuemYEYRFwpM4Ts1gB4qAhhb8ka3msaqXQarKQMUrRS0rvP89MyEOtP3bm9gnTL+aoB
7kdnlH+p41Q7N2/baaWIb60NcsjI8R4gUgs81n120XXRhiY7O8jbg3QmAWvz/rPAvJe5UVkfpXzA
V18E1Kyuzx5hX+jU0ZF6wdaaijCZ5bW9hjsiE6ZLDVetoG5qIRpGXWlYOK56k1s5oGxJ9LNwSuKh
wYaOK/e2nWQMBuPHbVPCg/tcELoOWTs+igzdOpp5k7/Ag4m4hd2OSmqvejLs6gmlAZnAXCU1XJUI
nI8EB3oanEaHaqcHi1+MmCea3k4A74qrrmJD9w0eZDqLd8DdM90FinOh0P4DNWLVbEfRiQva4vgU
cQKOOE2V3YQ7gH6dwrfOvYbasdgmAd1Hh9QOClJAsCypEiQQk0srLCJjPsi0Oc4FKnXApM3gqPgC
7vjyMNLAumJx+up/j1pZ74KNwI8xQzJjprjjjYDxyuTnz7jzhialpIo4vvGNq0ghOcCM/z5BZgRs
V66PrDLVbMswWHaN9Xc4R5RXkqtl7UuTZ+hK4SrJ9WDKQNiQ3ybMPPSXIqlfg7wsAPLl+/jNiCtS
QIdu/7+LU7RXvP84+twAIP9Ro7kCCsusw92mPWfd0XMSjf2JCwRx8B2/U6zVWpSx7Vu4LRDohNZY
5rI/+xJ3gD42260XUr9HSwafgdLADvIKaH38/AP6szJwibMfMFShSzgeKhJHHKrOSiqrK4bKWV34
UlUdMbRGUhDwiVR5T72OoM5PRQy6bLS2tVSar2Bcj4WA8ygKJK6fCDaJjz2GJNg+ODOps9RM7KfJ
220Exi8MFvDGIe5TZxKF1JoKwa6Fllsva3pcIfWqzozzq6KkWq1JedOOzbbm6oPTDcVUQn7A5kZs
3Aj9cwtNThxLq92awbdBM3WLAJqrkxVK2mRGKIYPIDyoPl5k/2aY236brTgT21GSQDHlcFERYfhq
5boRS69PSm0kKhTuBE9Rt1R8iPf+8/CkTkWeYK2DvFDEakHCabLT91ti5J00FqZgk60/ZFXknNmt
oQEqDCcBjwTgLq2BKfLpH4emCAvt7yCqzWNZTxk62ybMrmeotXtg6QAEFEWOQ6rQ/6t4nxYTuY9T
DiqKvtQSF7vxe7W97ffN4ETBFraMEjIc55dqDeN44bvrnOPx/Oncqhy5QIoRvvkuqj0womNcwjoN
1YT168LdtRq3uuGj1DItYPotV3ATTvEJ5EgzXh1i0WurKxwzHJQsVJz4H58yB+5Rd72eoa1Ryq74
bNCXrvXpCFhyNCej1Lhc7K28TdAAnSrDdTanO/5wXFtHo2FjT/duzhhnsh5Vmmjg0O4GgeXP+BKJ
or9Zz91a1x047pLwFKo5nMz8naVqorKNLPbP45gbL5NECQtkMkntQdZT4zQFNiML3Zr1mV9fa/ag
PdpTSgyL2VpfDuGiF0zKfuZjRzUWjYDXDZtaY22zPoe6K97OE4v4NbO/9dSqyRxtvDYh1fv9rKz+
LKlc20bXDcaHZQuHE9r06J0r4DeXZjeTqc7RRQOQ4FWsHMhpwad3hRPaEjxXv0EEN9lVsYs5zUKx
Zm+U29W/cldpCHk5uNDCQtw6tNrYKMFxXTlf3GUIQAun3PXb40GrZJ7im03i2b7//7NAlrWyXLMc
xfeh5uE5HYcj7zZ6vX3hiFdcCGw4oyeTdzwbHrW1U1NMdQbvgUconStAdr9El/YIrBsH5/faMgu9
J7VzMFh1gX/zdFhWG8SZ04sRCGTA36JpAFoct8cKWwX490GTFi6v9/CxHaxxNc+F/yLRg5C0qnxV
NHDbzFPEY1RO7FnYLfniVE5BfubsXckoG0Zty28pvD3J/P34Hq28RbWoMo+MJqup1iHCXRjLW2ZN
2XMgG4YAqeeZro3x7qj4mmOZQtChM5YZu2B1V6r2Vf14oCohTT2+0BM23RsOfElHadFz741IMpje
SYBCrPNIeBdIcDCe5JCdVn4yDU6htNjJLvxEacYVGr1KC3RaK0WFxPDRuhU6tyqcE/SifPdTJlo2
xheZVYuve3xqqZbXC33iq0GbWIm+OrP1Hce46y5lrwdqfwlc1XLNg4NYr6mTG6yDriMkB8316d0a
7o2rQsNhmr8NL+FlQ9rE/KYkzJ+30vOyMHcaMExXKXbuqO/cFbenvKNkVpDh6vKJmnf/KJ0Huf+R
s2FlObw8mjp4IryUAWl7WYEZZmm7feGj7O9RUqvB4AOQ2xTJiSwCDhSdVt+TV+/w5g90S11vEMPl
bo7TKfyCtPR1tVqd7JjXa6dNiUSybsoknVA1IfbegpZgDr6qJmFzojl2HWdPTgkq1WgeF397vdmh
+H/LmHztNZ41DzUqVpW91NZAJpe6SRpjSl7wduGPso/Pg3UxOzN9B4+++QNQXrEm74AfvkzSQqTa
81KklBvTldEr4I0bI2/GjD5JAWjuNx2YUTzh5nVMGdVKgwAhdjj953lbuKHX5NZcaYeC5mB0kGzL
wr/s3x2mh3eUiKqQG/gK5ayY1EMyAgYOpL2MqhKbacG6dZ7O+jZ66fYQS5iAMk9I97LWFSlA3qUM
a6uBu2Lm1OjUwuOSyU9HPMsMhHuLUodpBkTzoevRAbTmGQVPhgWNKnfEgmTudQ4VPuBekdTCG46C
ik1mXn50LbqnYDHJbozu/rOH8nEsqLlDdDmJzan6osyYhrdBbODCvzXakUtuXEjxq8ttzEN4EVu7
msmEKb9WzMX6FOx9VJsvODF0p5oPOS4tXPGqHiRBbwNy37DtIfslECwJbSqA0kzRRfRrpiCsTzaQ
4/5Y9pPqxlGA90L2/1VMYo++qHbuoOhX5+2Mesh6KJm4idRp3wd3CRDJ4WkaypQ51FFJAoTXCbM1
xgOedPw5ZLBNXb1VcGwkQkMOmxlIU75i+cFABgPhKdjka3anIUs1FKC9tuEYBPzNOefjYM/kTnRJ
P0OKJAOwUBZCqpH1/3LHGbNiUFPEE9k25QVgvodZuKp0rd4mHWTkEJ7ygU3EmBr9gIkmqBswpVg/
Uxjvu7ACoaDF4htWgFU11A4ILCRGvHXoZ6G9li6e86oc++EieC9A9N0F5k402XXqKbzz1BAupknI
ITHZYzb/nJym8EuHpE8m2gPM94HYbnrDxwrgJ7wt57iFa0KMNEYexEQGDeoeRsRfPWzqrE0Ct6wy
WhAFw1Dki8DfQLM6szBp5ybQXqCe54k+Wrz7ufI8sRL9aFXGD0q+3/5GOmh8vvxI35xEkX8mEGmL
3k44BrIeqv/q+eMVuyFxCYBdg+7QrOzZTs4ewSdXLDX8k8elRBH1ePHdK7M6/5IgH3xwgphU7Paq
AC/34gh/sjKWIr1kN0EhFs3qgQKEvlCcJpkJsmUb1Zak21bYIIkc4ppVVbvfy6OqKzcx8FlcgllH
Cl0lncVie4xgn82H1/fIyKkpQLO8OCHc4/vEThDL6/5giYV51b85jH6zLdh+0zjWD58PWViNGp25
ka090n0LK+9dAV01uWN6XXDUoaJz3VKktXRU19wMHjfnwNUfgm1lQypwXgahNKxbGs+Anx1jMsvM
Q6aQiXJya+ev7NSEYLPZC/BKZRmOcrKeJwdZT1LYE4NicsgMdvTw7hChyDWN1kKnVqUbn7CLiRfd
bs7qhsB6udSIEeO0g4ccXbmIn0Xzka4/n393rAGQukaUkMZbdw39wbNC5MQuPpAq5YcemZU5UYGH
RjwToXu5XBAhrXsXvF86fb063WZtuDQyJsXL4Hx37+vD6aVu5Tm//UafW0VoudzRP2gF/l9hB7hi
vp56tg0gVlrzfvpeeVMgfjurQby0+72lOigYK6Pa9NbrHTdTC7OmOvLnXmaFH+sfNEyJjDobIT2k
EN6mgGwMU8Ob56K7gBu1NHfR5aGXCN1+JCoh4TiO/ZNtpmaR/cSyI3qbbQM2F7x3jBjMflFMDdHq
rUMYzRDgMbZJMhPKqG37QDv6ozezHnCj5z3LgQpXwhU5+0SEY7vCTpejCgZi6M6kLTrG8BawI/Su
ijCloVfsr+bhqMljygVpnPjoScc5Am0wgWiEZaKgCLazvHcJqIkSUNiLnM0l9+HAf13j36KdBzJw
u5yVY0GIH6FAByWCH3/+COjq17ua2aDVJV/34fSFiXCDvcD6kDEsqmhT6X2KlSVa22gmG2YY9psw
3wguo0+Z0tGu/5hNP+/bhjq565j3chra5OIB58vFOeQe5Nhypla/4wjG6cDBtEy1rhs0kjH1+uBF
YTAgcmRpwtK11QiogQJY1CuXsxM/Te8UqzwhzmizID3Tag3erijNi3NRgocaV/6FIgO+kKyT1WtF
S+5qWMDXxvOtsWNjyK68GiHxPKP1vjkMHwXPyT6ZOAF9OoheZ/1BOE87przCW3eGe8N9/jzswbJX
jyokc7cQyZK/ShsLxYUIef2B6fY5MCQMqgHnyrnulxVRIHozF5RBBJnk1Ysz5TZ58HO6bfYbcx1V
EO1z6BYFjwwnciP4MfKd0kGVnffM9TsO87GcFuVlxUVjBVBcehD24mnUP8ZYP2wwxbNV74AdtcHH
auVUzXBRb7eXCf4otH4i1Pl8RRqyQR2yQ7v2n0Ua1Hwb3q7kdu19el/7b3UWxDCQ0D7nC7WP60V2
ekR3CTWUHRdctj2wvmjM5w77DqLQtgLWPOPU3u35B/wtyq3zGoL0oRzc1/51WnlkLp9RVYSP+GYU
AEYhe2WhTZNdQ8ScZlzGwtra1iu5IveX5pdJNBQNF/9GKxSKS5WXkQoCYhAyBUQVNPR3sSW/RGPW
siMIVafNhFthR4q3BNx8UFX5gYcwBYDUPzXHZm3m6EKSncd3DYXtzdzlAwaQ/eSMDu/bVNIEOd2Q
NViY1VhHY/5B28qioTRNq1ec+7178S3e3qCh7Uo+De4qL0Oy4APCNLvG5Mzuaw67nuT5bt+INJCM
9Rpi03DGMQgQ6lyN4Qg/29wE2nTL9tY3DiLltE/FaEJq41HpNBFNyPstNgO423rzh5QLL/P7A23e
opz1nMXtns+diIglYYiPK8O9vg0mOv8ZauC10cEpmJ0FLuFGhQDgDrGw50yTv2Yt6DZ8HTZ3ieD9
H7u99HX73SA3LDN1lzCxk4OdP1xXvBAwBuyD2gNjQ4mINmI8q2B8yJ37lKKQn3BbJdmPtKEMKqng
v/ihq/au0jsFyTRZKavGfWCTCgVXLHSlJtr5uH8hNh1LhYkhaF8sCpBcg2jy5ymF9c4gYU8ZhUhb
Ua/GbunIsVbR4GQ4FgkuLTbi00VZ/QRms+NB3g/29ntwbXsKQjww1nWOG6HP/3QCrijhTIs+PBtS
YF88LsRA64UZoMjeI9RqJS87ZyrZSJqq+ZHQ9CYcNnQ8pqNeDhtFMcG+h1zFSfNIguZ5zZfUCC81
f1RU+Gp0+Jxk3PhpbMkjmaZNXYOUqtseE2I32q1FtIMXOEjXCWew5xPwxlMv6j9FaNj7NUcVX4wo
1/lQoZbRI0hgZwFqjc7mFkNIUue8mmwQUqyVsMSSVc/F4gUS1pHo6Z3L/EiqmEySsqofIuLHdkrz
k7L8kpTUqE0zNh9XSC2HzaYytgIo6JrH082lvoK18athNp5AtFZohP7ORM1NxOnUoSGyXXblc+dy
+G4bEIzBeSVmfHqPoKhZmJCrATD3kHRT2j0ob/jDDhULPp9LaAYf+4MCFYy9WwmrjOZAzVA+F0Nd
XAHQLBM3pdpCpmItjo91KBEHVzoYZiWW9zoQiPzsEsN1jFhNP/PVTJmnvIMjglrhsoFkjC9jvDtj
FuIZW0oLVLtQVFPVZikVlaWurahVki4DEii5Km6Qzo7+o3piZdCpn20/kv5zZeYQ5oYuiLDIDGfv
Fs1PSRN8iyBJDyidbSxPB/BuRNTQ+Eb++6KRvVT4RxL9xZ27BhIgEjNUmiSE16Bhsgui5yxUAEc6
zBq7MmOzMUHg843zPCyQagFYbLVOcHZwnr4qx29C01gYUQEKnSkaGvmHRY5SAKKi9E9h7bAYB+Ru
z8loR8ikqp/PFNio19lwxa0OAauOybdSOX7dICH1D27LYddsTBC9g1bJrUS7PKBPzBg+NPDevjJ7
MW2C5hdH7zDcniZF2BwO2PDXSdQXVA4Kte6ftmpqbWEpXvKl5LZSTxtfhVP16mhrtIx/AucYSdeV
FtmJDSTiR1hWnQkH+MLm/d7d9EXK89rPgJqCN0uwjJi71tbypStnzZ1+CLKZcIV6spEJtpznIHi+
/4J8b5YEMoJI5t63uooVpNHjFgWzxvwU5ha+YN3J1H2wyONh9DvhV5LKBkxSpeEiw050kcZZBwFD
sFVjcH0NvYQv4JJYOPi2BpWzzuPizh5+Ol6Zb58dyEv+pS0aTHFoqVLX758b2FIp6HHvAW8PwYGV
qzW6WbU2KsiTyvewCR8r/6Jz/2dBVxCLoC87FWeetkzgY5ey19EJNbx8Wuy1S5MzAJlq9cCXtF6u
gMf8v7s//LbogafO8fGYOl+vdkoKwGpgHw+2K70UN8CYidE8uQctibTPXKhWO/afaFmoMBbn4ykf
DXAql9+36Y/9ntfxbOG5cQ1gatXwgQxwOb+iaosShw3EklWzEOB9OfCmmIdyyM3lMupl4eV10Fxa
z5L2kdSFHcVR96wHu9vsvs5ns6NBttMKzBKNTrrrFeG2YMCslrnP4LVX7qMwic3QvCkzC/3SR+Qf
1t0ZiWD1mqs8QbqAewNtdGRm81xA5fX1tVnp49fPfkin0dZkggUpV9F2jB7bQpLUHs8PNTZ5V8mT
2ZwYp/NFeBVxUNFjJGJeBm68prRbueIMRSqsFB5zwllyV6OEN2tha50Phx+fPrJTmrFxz2t/Rot9
EBH4XGFspPSVUiaQA7p0fC0Rq4VlmZ4Al9WchosQpq1qHbaF+pWdMiD8T+nAcX9nFSsvPefIwg3l
kWHApnX8O+FVfkijYTwGJvVwslaltjMRDNOxBiri4fCNvXMl/vHe5f6ihs8/67QNvXbxFAT1mQjG
bIwWFT6V8GF1A6klmjGJr9PbOq13LVdG1ryj+vwCMC8WetJUp5iCLf2mewixb4liGEI7DFtrV5H8
7EUA3px7Dsdti231Q6lj0Q4BWvH/iXFeoDHC02CV29iaSCIW8wVzPfcjPXg6EBrVA5HqFsMAKTuy
kMQP/KRjkx8+51Q45TNpbAK+cCcEz5UowssRNgzaGAiyqbxDQ1admUsBRvi2dhmTc7v8Y7tZzHAE
UMXzuN4jhNV2aACxDE9jGHJJen7NoPOm9zLS4glMP9djm/nynJChhO9neLln6uWtJmYBzWtyMgKf
VQvPeIusJVES41lcaZ3ot2qFu8zmX2QZpdnFYNm1EFvQYFd00gvxmf+PmT03p9ePMesMb4DgflM/
X2Dj2GT/cPjNb/Ny6wOvOMnALu2ixaUD97jChVR0aZV+8p3YwvDG+lQ44o+K9xpR+kDpShYAx/qn
/egpy3vr9+fY0EEOWq9/tf4zvKT8AGH26CFYM8d3Gnrk4ss0fXA9h/E02GAe4A1vLrhn47yA+1s/
5YplVjj07jj+rR+EFvlMp+8kGJiVLA1RfvHoIsMj5JH1nimrWyVBPeoYlrWq1CgWBpiIYo4EyaS6
knf+sNLVgpCJzyeoeYvIJUvGI0OWKS+5YxykQx7im/SlJsKJ2bGw6NGDEPKZH7GLUalbjIdR+ziI
bDsbBQize6y2EXcalqMSzemTQxgz1bPQpZvJEP4ppAaJg1scJy/74vRJpiBNk7xkJ09ZudBatvsH
2HXffQjBugn8rH1RstQl6Aowwfa2wXMVwIztRcd1NjppvpmzsUazTDnKbotudYQGkwhpKOZKijU8
B1bcKnFhj9TqUChO2Ixu+2YfjGtaavUgzGKmO6uNsl7u8pNJAhB1dtA/nyzKPh/1lZ0hM6YahKoi
YqTBxJfN3d8FXDDg0EFYu1J/G0uH9TmQQpgK9J2EFcxcB99KoqaaejOkWW6ToF0MmrzzWY2oMom3
tBH0J9jvXDbyM1EU5s2zmn7is8V60bZrpuFNCDNihKFpEgpJWttEDjoG8WfJuVL/rJtRZrdL8TWk
bQsAK8OEp9LGvZpy0bMXfhEA4Zu9wCeYaZw8QVxV3JyLTY3GS2dJS9SM4CIHTIwy/De7SoRnexTX
pMQ76vNjh7Hx5nFBhjZsI3s81RaamTXeNP6jIs5ty880tdOucpsu+PDPwsDnS7IOS8qx7gHGjwMF
KriwnHB8WX65GEvVQMfvnZ7for398CdgwW9r3IVdy0xLFzxIEcF8ulgGnirEvcassyHZdpwGVMpx
P/adKLv4FT6j8aZIRigbuPP9udRD669DTeFZYFwtupTUqkInXsg7c2fs6wOKguMw9AzaP3c33dQ3
Pho6UmAUTC44E1V+eTqC+09PCTfAqzC2aDx1rZrtnz8/xkopmR2EXeil8gQz62KCgugcdaqpdSDo
xlHjm1GHx5Sz/JQkDAP/pW5DNPROq0P9AzdDMdLM5+nZLMLyR3OzPfqbLO7wwesUQ0dfAejRh4SV
UaICU/D1zGs6bHkii6eBisMmY1UWXnCCVnEiIzBZmEBLrU1rBh3biTn/dFfWdPh2X/homUrospU3
USnSZ2FRumwB6JIY+eIi6KaDhEuY8nxi2VBXcRzvx3NahhS3FBWrxYW92/ZWYUoF+gvSDUvEXSeX
LAxn9g7gBM9KhgBcOKUROKs3jPteYYIDml7HmbCY0vo70hjIUsJevzgiy28oCiumQbgQYyVYcvbh
tBQrrqOtODGo8GyMxsKfHV3FFicjOwTZKV4tp7THgSbomtBd+BXSX5PWRzGtpCmmnfaLCV2GkIqq
dozSPHKHyGy3N6GCxmsKNojWM6t4fahj6u79oz0BmitlcYmku2bL23NK2m5YH1Gug60SWO+uqjmd
84iJBTo9uSHf2prXHVJ+2JTsRk7y6oIqqtp19+jQn5Rt5Kp/TCdh5PhNuRonyJI0lX6FmkXkyieX
OQQ3JXRaCKThLh6soWUULBUPttZfnMXY4sFC1OxBM4JAFux5Fxih6vxUJq7I2W9clWU4b4yG+TBx
1jVqihYqt8lr8AJ9gdpVZtvIN7haysDCZfhthYYTych4d5LcU5YcMd4bSOG73hpfy+Cynh/+P3ls
xFyxSqoQkWeMfx1Lxe37601WEvDnnkROorHQBWDwjwrVJ6+HctU3o22bSP1Xp+x3OsxN6u/y99q7
k00+EKInNe7J60U2urbffsBoGdX4BIQsDtA58uEQH2hkeLXkLfU8nHL3UomoIZkgbg/py6iafXTb
Xk4RYYh6uWJ/lNdZW5dNK/FYIXG5ks7R+kQ/zaaVzFHJPn3bHu4lB5cMhKAAVp1kNTZEAl0fP+I5
7pd4xDpiCz8HtJdlGtmp95esoiQqNaP00CoIgBV0ly+CcgJa9cE3HqZjof7KuC+cnH8Sv38z8G+2
81aAJfjEILpAfw4zB+tTWUnPBpH7h30Hgq/oyETycIEJ9M5B0Kwx/tcgj73EbXCznUuDZ5Yw4hze
g3n+NEwedANcvwxIiTogGKE+Xsi9+dAQ72XCKXGW+Dv31SGE6Mg57ECpdLHrwt7/dGACRzIfUvDt
5n3p1Y4wVL4j3d6u33++V7pwjeFI8S/+GQM7irNq+6ugrRCmUMkIhFy97zutaPxeoSdLNslKAHzH
f2Hw80UnauO8Vo35fq6jmw0xy2kDU+5z/OlGAsf3E6hsa/mxPCB2wtrYbC6omPUeu5uc6dd8fhWA
ETaPtSQDOGGYySrHLC5RR3tMSkFOXkO8xqzpRMOSwguS1JALjOD5U0iyR1Z9/LvMEyliaFqqnccP
bzdohpnZewc7CNtWn9tBmiipj2dpOQPJiR3htE/Zn2Opb0Z564Sh8dzIBa+4QTOAzLKuYlpF4bX8
BtN+rHveWlqG7hdORVL+xUMoz0TC04bxGdh/33R0kgkQSpbE5WuIdQ3FZdB4Vg30t6kav99DbkW0
o4f2G5jIRvxOIq1ppajixE53s95/bcHkLA/FaaANY/ZgBPxTl+FDT6zbrXJYPXZB6jD3vQ2Iz97S
ww6bXLRlooze3HIwdHrW5TpNtrJ5u7BduA6bGxmTVn1c7qN+Q0+j+bWTXv/86gZAd43UWgmtsx0+
L2qMmamRCa5lQYDd+OL+zHxPPNGi1mEQk6dLCtLClo/2k4e8sOsMkgCmQXR/FauF10WSqVar025K
0xanClUcCr0KCcypaSp98DoU5YK4y4H2OyRxkewzkBvg2CwCtSoLCP6zf7cqtTUdot3EJ26VqWEK
RqEtwLMRPqxFbv9dqXYJUtc79mwhgkg7FsOE4zcOpmQqEjmLTbJ/IhWqZnh4fjVJsM8M22QXqowE
lCjDy2Ht0TpiclW5POUT4ThSVJJhdJMKlHGqltikpfBJBBNFLr6M6fEm7FHcyrdR9YBw19swFWW+
flZP7Fs9CPWkM0YKNdCn3b8yLb2BfqyPHbQPrXjbaq0jcfi77ZTjQb6wTa+SuP8dmUBOrclRR88l
Zj/8qPzhQ7A+dmgG3gBTfILz+HMrYSRbhjUkh/Hm3tzzg2F7rAaYo3xKPKaTcMC6H8+n8icy53r2
a7MYDLMGP1eanvALEIAfpUIMrYjPlP8reOU6qMkUbGOFNykYwlAOKGD9t+dAmKgoszwsVtR0CE9L
Z9j8fAqlR5Xn2fXvrkaLm1l9vGizxq7mwWxiBr9N5eLhRfkKLVsKGhBGgcHL472FdS3o+/l/+eyL
dbIJr9819HMuRyFKNusIo2XjoL63y1uxkIuk9I1SgnO8sblXcUC82BBxx2/7DenJp0NWZoQr3HQS
L145dXSt/80soBdhacUGawW5qaqvDSFqR0GHcuMlsUmM4nKZuUCRr91LaAol9tQSeD4tQwiwvCIn
XhFHal8u7ATD4rRTJud0VMXcA7a3ZdHaLgGdEESuJmx+sdymZ8yLab/3vICS+Knb+R8/xWAAhXXJ
fo4MjUsTcSchWGOnd4aM9c48AKigMB8cJhU4XWh3ILyIR3T6eughieGYrZPThzdwJWgpWmAT7z7o
kbe0ZoDMWqRmVfmorXYqSzyRo+jZKCIyoPiCtWAQRtA97nXFFQWGV9459DVcahRpqItyp5DbiwMl
TALLgjFkeY2nSS3EeKmx8rpUrDSAxcG1an+sF1rIJDVUpAmM4f9u0eqYrcued0Y/FO6bpRr3w43O
GbP4lucAVYGHsXzlZg4jlppJj7NahjTuNHvXqtQlLoHJLHWSlg2sfRpVBKTOxNyHvAmAiqC5oXil
o0bbds0AQmfKDLSmm0fP5GFtYQ/S2Q/y1ovD9Mpygi7EQcFjT280Zy1pld4naiv07n6hIIQgnvEu
IpdC7pYNRk4cwcWnZeBKu3rt5pIKELWgGABa3/29Hm7qXrVsbrAfidw7LJR1QHdog7iTgiwV4r5j
ODuptMOCcOUoJfJ5KIYslsu+mtxOJkFEvzqVDkdyCaElt4vzkx7q1tqUmu6FUy2JZgRuO85K9MS4
nIacauXk4MBkvcsIm22tHOIQX9P7x90rLemJTOL06Gj9ZXzwaBrljobeRqOByEJxFuUCGbwfFwPH
xel6iYnsC3ashemfe+Rx73YvLr2KA+fpEOQzuqzI4C+ezcowIgfAtcc10VpVx077njylt+QiFwrl
gVgSn2GR9lLaK7pfN0X84qCjIw+FLop5kPDU5Kst6l9LG7MplCf1ACMFz0l0DfJOWf3U8xl7JnqW
HzfrBMk9HakUK5QKPZZSr1vdsqVHtO4HcnDGYhslDgj9TLulnA8h3GvJ2Gm7eYBg9JARzbu69yoU
RPspa1s6Z2CAibdv4HXHPUIqsn7y8fvPi03mExMtTgpQTcsVU7YCN8VkNtJ/LOlepN0t9GKr2a93
ShJcJbTBiI7CPLCN/T2bS/sOGOcZBOLKoxFpEXc/5Aa/zFf2FRoh6NxBgKyOiMTuql8DlWdkfhSn
kX0Pt1tIoSLQRsfslrUTyYuNtlAV8fkgeOOo/TNXnkMEHl/afpFZLV4OAZ77JdSVWSiqrgVIt7EG
+5mULHImmBUL1DyShb7yXbHnOov7o2LV7OfoqwtkeUSFyPBMkjmJMm8eCp71duKdxTmUTErvhKTI
L1S9yAbZdnSrxZ5usDgtVait/gX7jpqbo8PxXuHVThPuBF4kGvx64PBv5tdTmmO/fpZXPY+FtG8U
a/5JkbPZPn2yqzj9d2Br8TyY8ixZ8ASikc6Wbt7hxPEXJKAkAbgE0uwsVvFr5cU46bK8hG43fZ03
gE2+IBDXVL6h7cKL9IAJrSzV72SFkSVCpzIRVjXXv3rVA86x3z0eSCWHKwdHQ7bE8ijnKTBfajsM
Nn3n4gJrilFbm5Lsd7zGhQdNaQZ7l4HRgEz6orSCNNpDfDCDIzxyd8xmmZKFUlCXgF66ud2xqtyg
HEB2I3tIB9QOVsRkVmDfBVKmnyPlrMdiSIOFkjXLDCouvc3BrKGvk3vUi2rZWiMrAHWAg1jBnOPG
h9QYpknVsgkAQg0V5NRNt6FkttsIh9dZLqFvsgPn2BpMcNxRmy8+OVRqZx0ScJ15b8YwFRoKnGV3
+ZK7qjFK/IZ14r5EFps9/g4uMKQXQ5xnoMNaW51KAEOG9g4jsXlG59815k1K8AJ8Z/d/eE0pjRTq
iBW6WK4wLh4Jh/EbGvxh74+0Ao+qmynCKu44r4PRt7V3cXipn26SJfLBOj+rc5vTFeRtmevGC7Q6
VO1kOoZhHJ2iEeF4/LbLyWzAIUtXExsJoGvajedZQB1U4ApoR7/GOegzLUJSa1cx+BTI2SRpC6k7
NeyPVhBL8vQavpfwyUqu36dRKHQVm6SQkJjvy60D2Br9XTyGoSI7oHtxSA6Avpk36OjyuhG8PARY
c3hBtRrv6O1IEc/cgklyDE2ABjPNY4i4/QjzwbjN6Jqp9UklE1SDtO4vsbTWd4K2KjRnIPG+Ha52
XYsTTwyhO8o9wiRiJ/IKJQE4lNNa+JuUV5v+DW6ZXln+gRpxvzuLux++plpkOwZcHn7lwwmcDwPO
A2LXw35Vcr4vYc2ff/PxwGQlqJsSxCa1sWZ0zYsmANN9x903RwKbUSL1lt6xZx84GHuTTTEQmOl/
e1zAXOCbiAH222as3/XgxkGierkGOJTuHRhs2vuyET8GrJk1QRalB2A7lNH2Hbzoo/mldQ/dZSzt
xOUtn5i96szFqdttvaqMWBXud7RKQTfvlQ3YA4/lu2lI4mCo5khd7GbttV1qNRv9wsTt61yDqi+D
Zz2iKwQI4zZlTGbNIPIK5YvGQEuNWXybRlq2L3CoUot09urecS9CLP/VP9Pwyysx4W0HZJDyq0PU
n1TQ5Hy0xuVY9gr9qLCiKvMS/pMsjZuepfrCmJTST50LOkcd/uVX2UjUHeQf1wtSqfPJuvUfRekZ
WT+mittVa6CITDEp43bFXLLOibve4OR7aWbtlGzwNZ67XbJZZCkZBi/se+AIGZK83ypnsUdFkQb/
4Rv+49GiCBKiNRmyZM+9fAiZU4cPgGxy+KmmWsMo6DBv/12AVC8R/S2PW5sHTrJhBXqM2mB5/pun
YHJrT/+Uw0zkIaUUYAP7Jl+FP4os2zXO9UoRBxvgQdyNR/mj2R7BtOcKqNslC8PZncHYEH7TTxJn
yU09M4iz/9tQ5/ny63cEo0FzVcLADsoVGH9UOdn/PahyIQuc1bB8ibwsvCD7CIrVtGglfFM+mE9L
C+fosE7WqbSNEaidz5d9xGmg5u3JWT76EGvRlaiLr5EQ+2WoFK35VHx2532v+66tOElD+X7IjJ+b
Mu62+UFrPavmS1NVaEDJwiOTOivtK5VKLfB4trmZ0YvJ9AEMdWJbrTa+9MWNY9RN0ow+ZTw4qCC7
JrOoChn2yaCT6h5LDBJgDkaLSr8mc8v5qZH9dqZDDE+fIty9MSpl9Z2wZ+x5oiolPOdCtQbFSHHm
tgPMwfCHAEB/xQbV6rUv7qExk9bVeZDss8eDgjwnD4IAJCQ+z+5/a4QK09FeLWfftxJQcgl4jN4e
+Xjd8JJxiwnZHNkXQJ1KlewgjXsg4Qp1PMA0ebYdlBuos5M6WE9fwr6fePJwN7/xI1a7MlQG0Sfs
q514YpCRCj62myYhQf/xahY1I4cKV//rUrfqfkevqDSlHhjlpW6zkK6sSOWdC3pzHWw907HcQ9n6
tZfIBiWTUMpYUut58sq9W7LXyM4EFxqb7CVe08tZv5aTo9LduqEvH6DIVcA8fv1sSakFSulMiyYJ
GlSUr+qpeQh7u5yRGhrs+U25nZNZMgODW0qT68UCbm5VyWVSfGHnAio0W40O9f6Yy2d1xTESAEdp
HwAhZZ4Xs4PsBtMU9sz6vcvKY5OYM7Wsz/qu2SQhVZCho/ME54Dnqe6gkdf02MMFz4t2ID5E+1j1
ic2JcvU/dsQOM3LGlRhALQsBVVM+Tn8yIz/bUmFSGnEgjljobFoxRvJqO0zY4KfqbCuvMHfkE0Gl
3QGXqkjp/GyGCwEPKByhwkNbUT6w0qBmM8SLajSIQsfEhe0RcwargURlklUbAUO/ljfBAoYJSiXG
xKNzEmR8vQE7Atu8HjKct9XT12/RqYd2L1f7BRQ8YJyASijYs6XY6DfwvCkyyLwZnW4+knKJps7Y
x0n60T0MRSHyxOWDB/jcHa+Qpt3lflvx/5fptDzMeC+h24HwaYtiFkGzJFi6wP6OCY5fRnubMsWq
deSGiz0JJhDpVI5leuBwLn42zyKKsUVHku+8ocaG1ItuDvLAOs7bXQGXazs21WcLl1OCV199EQD+
9ir3qrhaTA65d00jG8d8zvr3CvZttfS8/OG+VppDv+VWa8yiL/rSJd/yE78Tp5sEz2STBte3q1Y9
XjLQQrerjOwVJGwB29obwH8A7FKEdRgt+3AD5kjYxMvbNfvWldB9UlRVrkE2KBKD7dpzZxhyQdX0
DJf8F57p7UR4AmH6Z6tHqvQCHu0/BK7HinLpiDs5mCb+VObyqaAh+Fu3mThjmNuLrY7F1oHYQ8qB
QoOrolpKROrCWtIJFezuQ9MUtkBcf33F1w1cKi4rDtnmHHOpFfQSHw0jnSU98D2JD5ZPbeGO1ObR
mN7idi/bCHLDniujR3gBsqV5bWSeScg4q3Q6dbc8KHh6mB5pMxvI0SDee5F2Y5IxYMtw5pOA5mxC
9/Azobyk8Z+9gK/TCe2iFsmbwKqSUwCkZ7FHeEW6GBhGZhPR6U2u/Km3YG5LeyIjimfFBlI5WPA3
h2pWP7+V4iyiWEtTH7qfK/ZYAEk1/yoWhMmyLaVFWcAWtDJo2NEh54apZqBHFl7ctvZDE7IgIX9u
gwWzKj50pPSZTxhzc/RpvHstSG16EOa6bQjIqBNH4cgWlui7aSBmiQtUjBvMXcELB0/QtouOlYuu
4ui9HpXee4yLo/Y4kk7GHhtZC22JNtltQYHM0w/SNhq203EbOumxj3Occ2en2TGJXRP8TrmT8Oos
CbSsjXep40aIER01vUsQg4xz21WSOlYiD0B7gg4u+hgaDAe424ORbCceh4ZEY9TGsHm3efujq0jH
ldgCrbp/5j7YM/f4a6psaHxEYBCS2oXxENKWAEiFAwsSHBfj1E4ILaur8O50QlQmrCcnRo6+WbGe
+w7HXAq/l7mlPrhX8HeAJZduxnjo7Dxb0hVTuOD074SGpjRJ02jKkypWDKa14MlecqwkAJA03hhQ
noaqIi2djb3W4grTpyQw0Dmjze2QiDnF4V527fPCwWG+oCPEIMpGLC2JPGtj1Gt8kxEmy5Tk7Oxa
JT5QvxDl3qlIOvQ03jhGjvHJuKYGs43vNoofPCEpy8SnGriSgaPxxVwHPN3ASdAujomPi8QxvkEf
thGtpzlNQxjaAcXhIaNkp1iaV/DtvQp7rlpejDih1nSbFntnLp7lTum0cRF1THB8k3qWhJFCf5W5
esdqNJNINkDMTQ1hwVG4V2P37ujypNdRXc60P5bVB/3N+WsauuUP4Eze4s3JKWyAwQ9+8KB5OrGC
jE95fn4wYjqahM0Xc+4HAFxeBrn/c6gUnWsDPbrV5BtaMqVmGzHJAbpUBNpcIi23th0nH9EyA5/P
NEHU7X42T0qrKE+BSH0Z7iQtT12kxbFTbCh3PVmJEDzsBI52FwlIU8FfWyDlHob/eiLvSuWCeeFB
LMlMu3XiTuhhaKU6IDgjqIAfO0w+VVSqVbnmFbSRPT1Ic3s6jhvNbDKE+fVXV7xPRktDZINn2299
LP1Uea3MEpsb8H9pYfH0vOGNYWTpw7tNiaatj/A3DlTITFiLTtnG0hdf07aVTOdxdEUr+2yIxiTf
BHRPX75Utj6pyOwJub3zVuHSK0CTBCMeGH0H0vlJJSME2X++nT55D/8lvnC07JzvpWmHgUXbeptm
CjDU8TFDMVHpV8hrqw5o44bEV0S8GuqAEQxd2GGOEjrzEYb5K4Vio82hoSjJy7kpGI3KGJY33BCe
yso9ce1jEG14f+d1JWRu57NLzohnEyb0UsIQ0ZvIqn1kI9BCBkiTbzjcW21b6DSnwS23Cy/FBo49
/ritO6SKlzklNbTstnhZYux87JokSDVs+FNFAj+RBh4qOZq95Fcq8j9SKlWB+qR4xIt7Zy764lDk
NiVXfuVWoJ8PBj4hzJrfxHLnu5n4RGl5OgvV7hpUyugLz93NeJDuTcsVmR9+aZpmltA8B6WW4lD3
fYvxmRtG0kQe3yiQIiimkgmT58O8tMB/wbPXlfZdJhmGtBLp3MBYPm5bchrvq7KEKGOtt+s1O1+k
zsVWTZ73pGkwwTgb2kUqrzA8XO2Wy0SP+vlBEkqme/Aq1+J26Bq5D794VyQWr5cyuJ4oUJ0PD2HR
e8VKmFz1+Yp+neN6bqCnEb+0eZ67Gr1fdciN95VGvx7N2KCzG5DOelevBGIn0yIRz+nlu5iKYeHb
YQXg+SQEHn1vwKwit7hUVRLUTNu/BLSmIj9hEpBhbeLk7/Y4U3+I/K5ZG6XfZ1ilR4h2VJyzJ7qd
4ZxMlTVrGYBsS7RawefxkAIzL5f4rzW9jbVMvuE9mxrKcpOnt+sFiZn/sgo4sqSvQs++hxzZeaOQ
m0F0O3Kwr5/9likWiR0YLin6qtSg030T8AXv8ONH5Prn/61uS2mpVD8BFLwz/HOsX3sVHu40/FrH
dz3Xh9xUDm3d/ed3pBLbvwqvJyaltP+jr8iTCCwpoMu851Gb4lnXllEy6fMKHBimz9krUezqXNuC
RX4gtKO74o96cY+diR6tvAGqm3PjvEmyNYeNg2JicLjJ3CVDPWfVEpHLDjbTdOGbMYR2tr5QuUVf
yB17mCDpmYUrTwmceP0dEzdOSqDn48fcV17oZ8gfmVM3mubd+ZpiwBP4EG5TnOwzQUWRCQ15ygAd
AqCUe/O9CN5cUV20LOh45br3BJ5fRqdYhxJRrxWeusKdv3NfT7WyEvEYCP0lJOn2kY0cBvO44JY3
GHN+ULCSQk8zCxr+zxHSFDN2LJNT8N903eB7fM6HJGIj14CXUo7pLSmwcBWkYb8R+QjqRwHbak+d
iWrItuRJQf8ZP5R/Tulk430jvj5iJtAOZBaKtIkM/PVZUNz2VzGTqoexi9zVeGxFblPwB32VCGq7
FgE0iByW8nFrj4toKfXDblkkCTeuUg6MW22IKxIg5LS9Hmr+Arw7XPqKQk2N3JV8EI5Se2YP+Gz6
UE5aoLaJ1/HOQaARtPlqN3uH/84hZIffLe4PwwCGDjSWBEA9pcgnXqBbsrXXUbhRvQfilyE27oLf
YJWwKV/RB2bpPmBtLJkhI6amavqXPNuwDD0Ny8eBCRNzO6VYpp/vjPPlS/HiteFEqLrHd4em3b+m
bSp4gZ++IvgXdn2tdug+8V1UKvvE0q8VQ39yJuWAN0U2gsKLmkYzArmSNCtB2cHWOpe8eatvb6v2
zBeKU+oFaSb/41gXvi0KWDSM1ky2RscuO0LZBGHBTVycuREQsz5FJSBclfqxsD3BMOrMMsZOLOf+
jZy5/UF13pO8XK+lOQgtCWsRJ+vmjV3VSTThBVUd7uRZig4YpWHwJ6F7xvqh1BT6F2RkFdtcbP7V
c8C3XOgFmSrX513bwVmiX1ir7VYJKpuEn9cJe2zG5xMaoQBW8MZxjVDHAPuNjloc2P4HApzvwDXV
xun2L1zcB2kGytRyG+oeKGgTQ4qcUcyGI809cWfwIw2/29Ya0TuNEA8uvRexiEhkZwVzOmY+12Qk
74hueVUZ3hyyIbmzuXzeuYL/hRE0FVgkeDi6SG7JVH2gCRBvgCmiGVnvsbPYyic6r0upZR5KEGoC
QIxEzeATwGQPbrR+JjOigdVtnzoJhI1UnOxLJviF672DvnESAYMxspw+QNhWvsf5JSjjAD5vUemF
d9MhEZN9XVqNuLGR7NK0QNDpXc67PE/i17wJaBOUdHqnIeE3xkN6ldilWCoGY2GVtDwJG5LoyC5c
H5w7edOJ//bpN83nccG/abQZW0EYEIMx6uzdYn7TzSkC1gh08aZaV+tvaDj2zok9+phkyl4HnJw7
mu9vMtWEB1OXE23qLO67axZLmaJzqcklr+s3sFHcBsJiuGeVmHiKWm5s1/9SepmFpBUXMv80Meq2
3QQu9KeiKEHDFotdPAyjD2dfSg6sw+5N2xVne0yhXU4im2j0087h4WvLWY1MN5cySkvyGhxvR4Fb
KzW62HnZkj2Ui0IZmQ+piHkH2SHAo72lBOPpXShapYUoqLHEiUb+qwgIk4BOQ7okFMXvr1PB9fT5
W3dFvWcigtSdDbxgyE/MIxhHDHOsMjbEh1jLQcvbkM5oculNP66g2iYElHkBSDPmk3DWwFEj+Pqq
hHeNgS/kce8WtwRUBZkjCr+ZcUEh2pk8MXnvMgsNzglse1J+pnTn+pT81JS6sdA+VAL9/NaZaiGS
W0dTsfCKksglUiQtNqle1kwVbzbkA/oAZUlqxNDt0hH4i9ivEq9vgS+xLEDLJ6k9I8eZKB17RW4q
LjtYzm/xSCfbGdXt77jq0EUQuD+sJGhK1DtpSH8xVI58Q09pL36uGtrEJSQj0T4pX1m7+qP4U+Oh
x1hEXVJcNS8im0sjJr8rIOjwitvjd/yjuDfFH3/UqKgWsgr/xdE9h5hl5LRLaB4XsP4n31etdKmH
ySFSv4qlGK+HQyCxvQNhR4IDN/OHCr3phQibivZhuMN/XcCOgBqFA+xATEeqkDVp8UU1TiNGiB6H
+XidWpnJdBfpPCOuy18HNmm6zev7bbCcb0yarwYvLZ1zbCb1LHPGmLk+i1ubViTEeMD3CCYgfuct
v+ZvW59t3sFlBxTcE1Cxiq0ZB+AYLUYGgyu3k3DMViNYcHu4fwyDuDdKkso9s1Ah5+0eAducOAzf
2SXoOc8KHjXLRD659tjgZn+xXreM7KpVhxNCRkHcF9Rqxdtl27fApiQBeIo0NKYEDHL9DlgHto4m
/i6t9AqbcYI8D8ngywsv2WTT64Ip/Eaof0gMLXOLG3q5Q6KIJyS7aQHh9xdwCLMf5nqsOsgbO67Y
9uLWd1BNkg4EUglO7OIQi+TFi13s/skSM6QDmotNvuSruEd4v+vSi7TM1UHm5apWdluJ7iEXEjEH
cnucJ+PTY9iFVWb6nyMY6mHzwlRBObXlrZgbZFAojm5LA0QnOLR4VowWViPp/UQqFBQlWuOZtNQh
Nw7Fttc61eVDF9iXB9oHYdcRt0KlMF0eT1flVwYpSUJlwTGwuG+fP0vZOTnoNHcpzUi5RIHVvHwq
lXND0rzkaLkeWXHWgHawQCtbTivzln50kx6o7i3MzxxD80hMw3tvFfpLfrPVCWiph8m+rWLQiIjs
4OxI9CKvmOcGi4/YyD/Kpj/p5JYFwgoSVB9fBv/Vp5v3JhNpvMBhlAd9w8uiofmq6LQjC4IplV0b
5121E5k4Dp2Uged3Msc74lJDgAUdS6peOK5eDeMiamp8bn3aeYPjLk9rgKgVigXKwKaZB5qcfPmc
EFJ7vbI0zqad36kr/IhFLfMW9wD3a1vI+MTsZ6YS3uAriRHoGGyIjRCH2B10Vkfd+xFuGCeZFcis
0SYY6cGSpkRE++S8rjl7gnyMpepM9ZWmkfOeiVuan4PCkQdaJplBeCypFjJ2UhrvyHlGsBDuP0EO
rEACMaPvSwBBjUSV59aETtlIP/CSzmTjTgffDRlS/kfNg8VFgE1fQRB84VjdXLgjkHzSdQFX7zSP
Ha3Kj0AF/tkCbNlArUyQMkEGccoPocE7rPlNOHULci1/WjaMZ5ZTSK8hIiBwwqLxsr/wAE4vDvAZ
QOt3pZIzKwNhSB7DGzzo7Xvhga8xdsl2mx6gZ2j2sobwBALCHgo14kZ9uxcH1lHX34rESk/a9ZdG
SvNWoAsfwp/6jR6wIwbhSmyMYuKAlNAejCMXZsdOg1ZtoX6kqDfF+ObNQTQP3qtf7iRI9dBzfp4m
k+rOGUw0OGBNRgmUggcmI1bgXIg/Kke4qxsKxNFAmQqcKjME8p5wqzU+qOu1QPJ1wGlkg4cbHL98
PSqK8qBS+5j6vVcrr8OcPKgXgTBVM3LSQ8uCqTrui2nbkJlLxIuA8UICTFxni9DurW2Uv9CC3ub/
RGBiD33jjoGmWUqk4tYN/+dLnHswgzoVKnjpO6Spe5/nZNT/eL/V05vMsh320XxxMSwW17D5bELX
CKM/mpeYbilZqFddRHHTr8tomA1I+MMhpJaMGR6LkegTpDE2Alxb/5RDmS2o3dhfQvCHI2WhO3I5
AyT/8diPmgqlX5lo8elW5RiKw96zRMANG9e5sIa8Kxim6CNHdGHGtqSlJSTOqaYhx8eD8Jw2yLI+
H1s7l3nN9igMUBWTla6vqUfEhd52C1KNNmriq1AjHmfkRckZj+HQkEnzzVaxSEGraAGZtzCTaB4g
RUUFjH7z4h90gTmt74ITuZD13EOq3DEYrl22HkrHak4WL0k919KETrRY00vxYuxURalP7q0mumTL
5aEvswMelz+bXt11BFk3oQtduT3oF+Kj8mgN20flpRNHBSZ5iO1/muiSaXVqbdY5MX+p/tnGll/J
ykgGxpHihjESefq+KAy/1y5n5sXi8EPTEVR6kFrE/PXJbs5gQ0F+qAqysZ5mNnjbZyaSQPWBWp8O
D2BGhh7FgEOo7Jvduw1q341cPg2gmhFp3NzA5l0eNba12TdTNVJMPYTSesWc0D5DNYU+Z1bEtinA
y3hGl7z2/vhR+POogXysPu3ATSeM7eI1TIoD686oyADXWtwcor1/T5tOUl77GM1t6J6xmcYDtjIA
apLLcR8I1wj5mGY8koPy2uy3R3x1uYMjiNPfn2qJpNt5aI5YWSPU6uMo+Fs0Un4SrIxtao8XaUEl
qhGzTUYk9vpfl7efiENY8TUXNmoQxfUSXkrFqSW0m770UEJpEWFYwFy+1qBu7x6A++AmT3CIwGoY
aEWlYe9nsLthI6FtGm1xsBWXZgi3GvyS73/ssspgHlyWz9hKQRz8K6tf3M8Tag3Dx64oodqu/c44
ve2gJcVTnkkt/UtXEhshxdu5JfuPI0sbvAyOVkoeUl693H7L/RIptmBkPvL4+O9b73tovSgs7H/c
FwDLNE6wKuuhh3/USIU1QizZ3GTYYSkAbw2mIeRz4hYD4YzxsHODYM+bRo/N3n1bd882cNlku8ZI
uykiFH6a0dzQvgyMLLzQwBYXXx6iJeTI0XFYniKRgQ+xlXhJS6dt+XHyCdbtqvYE9XjEApCR71ud
iD6ZozAlpGLseEtMqlBk18lhiFmNfXKgjyOyBvTrZBw+/2APABGeWmg8S7OfYrQ2OFZWFFXrQEic
xUmmZnhpsQ6rAf+6H9ABcOhhHi2Xuq/AkOdEPTCYzmfvSXkqy1/A8AVVA+bxb0hR18o41qj9Y7kg
B18ds7ld24HwpvtH0Lh4wQln1ryS+M1j7LRpHa4U81EwspmZvuTFfiHAbN/cxQ1AydtUuN+C7wb2
3DXuoP3Mwav7gxyMcejhUsltz1yRJeK5FmlMDMqtciupyFCsmg5mgRN3mrGP9D3Pr8aqS1h5PcFT
CICV56N0HMtASQBA+RBHyxVpKGnCPgcdLiohbiaTIuLAYX/NCreXYcci+z7VnDQYKlFbERZ/L7If
AHHZoypGXJbmey7ZeEBD8k4dh8sru4khR/uX64o4+e8PgBewOo8IHBPEvOh4FaMK+ldXrJm0fTJR
8+icD2klRni3F3ilYSbqbOWrbZCWg5HalS312OVfxXS8wfKm7NqHiBuiBzOOruPASpoBBv8paZ7t
j/5pxjZfspAD98k8hbQ8q14LStjP1QO2VoJLbgxRYLI+BxERB2x66HXz06NPM7hHORU0Mu0LDPD1
2iFLUbycIMywdHMnkRdZuEy4VstyANLfuA6LLgvrrbiESzHBXWgmentnX8Ud8QTa1fvc3zh74SB7
tlc6mWhw35S7YHatNuEbWt2LQf7c0546pBIO2wRWY85e7kxwNHRK1h4aa+DKF5zAAij5ETV/P6Uh
mosd0+2QA5E1RIKsGiXrU44YUmDum+8pSWktZN8rcYe2IyuihfFuwtNIHg6/h4i5FqInLgh/OH2q
IHx4FRN2bp2kt76+yfLV4suMZFoQngQ8MbrARULvqv0DvsWRSm7SSTXU+owzShuYWZDhZqe/dbnC
avb+ipeGjlpfLE6HPt3HvsKl9koAKvkEkDP87EEITx8Sma1Ag27gKBB3J9/V4kdirOoEHWBmRcc2
lM81MMke1tYygXkuFDsPReNFj3Qv9jkPBWtjhLbFoSvVyU5ELXZpkKl4LGiCdVY2DRRwAr1ki401
3eWXxtZaafleVutUWqbzXR+5MnpUuuxT8yHBI7sOcqTctGQ9zcc8Yl9y7vj/BRqDPkqo+8m1WIw/
Qm14p/i6gt725EutFxUsEeINAfeO9Y1PfIq0rxuDZ/z0Tmj83NXt4NReIh41Ije8ni9P0sDLzMpY
EEseHVeRKdz302MaDUjBKh5H9bZiBjcHZC2JAc/W0ad3B1ZvD4LEARublRFIzXPfMtAxzw4PA8yA
eKtS4trUXmjqN7/qr2Kpk0d07f7grs8F84hwkdfFUhvdZq2Ydvm7jC6e3uU47iGLS4fCsnxKY4a5
I1KyXLYmzFZNQq3x52sDc4u7f/RHAFLxxVhsC8bH3SLMFEmPbt3tF99qcF7pu2V5fWvbb/rUXWct
cmgXjYBTLZC1Qx2gYEkAaOTKZ23tmi4b+flhGoHo4uDcHYtotw3oniKX8Zrfjyyk37MraLvH5TXI
2cX58kzW5whaVQqyWAturR5bDxunqG+6nKpERkOMYERJNsgGUYgU3BKhqfyPz6gNm2mCP8uYUoFt
YO9vsXTH5LnsPLhbhMAz4K05CDGdFfkG4UupnLcHcXWBNMgnGTja651r5h3/0Bn1qRp6pEjBNA6n
f02TFdBLznijP0nZ+xq9hVaoWcP3b1tT60Ho/xX8AdNudA5kDP0wGqdNOv3VCZGSXx34G3pKLdy5
Sk01VzII6w2nCIBVExdRPXXbB6NbTdPB/JYUQyUticBunTmO7ASWaxl2PA4qY6Ufhu+4duJhu2qh
lvz+FtLFM1XRcrKmk5FNfP/jkzFoZsuqmWNwQiPRaq990pPs+Q5i/+oWGoGU9RwqpQB/6Cmmbe7l
T7oeenGrNVhr7c1rC007OQq0fmc4oIfOUh2Piehsd1yVLSYxAEIGDEHbkNA5N3TnFaqXI32Lc5tD
RzPIPimchPEYzpVEtflbfThG59e4unZ8i5W1cRwGBFhGrlDagxCxrukNr/a99PUETpRom8wWVaiX
9ZdlDysLvWI//wh++carBSWs0Xs5SQweZlnbpYxtSHjy2B0Ywkg+ojfyEXubbceD5wvPn2YyPoFe
f9wgDq5XhLPVlmBjOfD7vPhfYU+eHNvtvD0lTaHZz315qYOwleK1OkxXmXeRx80LGjj34IAyfWZ7
xdIlWXqLT100YlO+o80CXYro7XZ+ScLWtTpNdRKPAAnCEAXFOj3+MZ3kOfjHMTxnFVBd3Jcq0FnZ
L4Kyz4aeQ+WqZ7tJ+IsZNtPDhPvJsnGpqcx7iOi0uK2Fk0CfKHLiTBN4JIFOByxprOxzKiBoJiVw
gLty7pfQGDes4OZg0PHE69yILvY4KtdmSFRIm+shOKVb823TXNrYicv0uFNOM80xyiGEXdoCd5F0
kAyP/sZjn+727rEKlBVapQSczdAdzyEKP4lNdPbfKCOKvfLbG1atpeBZnq2yJTnLW5fErL9dsF4a
QpUw7+3HVva41eXTIAb+4a8ZqMxu1SIjk2zMDzCkmMs6vTcME+hhp79xvyFKKhplaOTp2B5mSAWy
WgLxBk+XZnMEaMNh36kAILEazXunPl5ABePtNNacjz4XhfmpWj/CFiizGYG0QAVKlL8Zn+/TwKdH
nDrgZXCNoAP+Fr3EfcNxj2HCTBdhqnTHlCbZNMlB06/egzo9ec5zNQdfZXKJS8BklVQUoWWDO9j5
sJ91FQFI/+RJn/6BY0m5fsDoAmSh6Ir28wUMl3U/HfIBGy6wMy84mXKlw7/xDLNlSn6OyDxuScPQ
EbsfaI+VnpQK378ZroB8QlrTCcIdH7h77KkYp2s+1CCRbkDSOaqUbiyBmMPr3snmIMhrTTlpUqWH
s2cYAqxdZZPqKocAKGgzfBZ+tSG4zZ0x8mq7ovuToBEy6QCmXLeY3AJT8nDF8ki7YtPjYAeHDxzb
DsvKZKaPulwkXopJgfyFpiwZYEJnyQh0FZZ0VDzdcxT5TpRPH4NRRRF6HP2OeNWcozG/O2GvoHV3
+BUnbGlyOC6KTVsO+1iFuJfVmkYOfsmtLBaelL21lUUXN7X/Hfuuv1qVKmv1BLPL33IRTT0x7rSd
LUQRuN40SXLQGJZhclb6cLBf/WdHu/EqzMut1AGyoB0KSIpdqzinV6w1GAvH0abZ9BXe3UXCBZQC
Y2GVyYF0RpHym9gMSzsegIUQ08HIncKmvu6ifjxcyqFad3CKfD176PrrEL2ZNdMx0bIa/SzLyL3T
32i/xpSu2dPY9znnhNQhr8prvRqs6IykDZ8BVCNFAuOAl+sklwJuYcD/JbQq509GTim4gV4Svyj9
NwJqOAQl7cfIbrxXwyZddyy+Jyl079bjKWf3J/MNr87CUK56awUCUKpmIJ/KuhP90Ie5ZTaB9Kb0
G1OPO4YpH7P5O5/qriPhIHCJAQx/Kq0QM02CL7PE3UNfKBBfWKTtC+GABPUOt33rG5VDkSQ1Z9+1
0+8uSWRHAufP25lAK5scIbxJ/MZCjZflT8GT8KGCuD8/FBZnsHN4+VGWs7/oEv5yKyjLslOMGFHJ
RM9qfcpX976fcsUH6TatkRdqY2XOyAg1xznskSqnQAvQJ95YUf17nrJCEQio1RxfON25VCRvFgqW
52qLmrB5YPfmGOjwtevgwVFLm0/yQLjV/ClB8rtr46O/UskjG50SRAZxKo0uE9tHymqf01MzJ3in
tvQGRnJJk9wxkNPjEze6nVXgYziUAPHPtBMImcdfdd1DbfbwC9F05nQdiVGuw9PomhsJ3IclC5nI
LNsBi2XYqAMAHkztM8xBlmBSSK/6RVxVA+m/E10MumV/C4V8McMxbhRa0vkT46UgsMkTmnbaQ4CM
djNdgEvxAYUZ/CYUyKSdxraEguaVJxJXyRPSvLc83cl414KGcJhP0bb1HRa0gL+Pb0EaBYesXe3b
rq+7o6Mt+WreOYY8IoAO8TvWXQZUlUYKdeO7jI3g63NAP6ZvcRoU+Fs7COnuXwsLUapQIBv8VtMy
vEw29Uql4a+kpHFwj0LhpT9uJC8zbHKHO9Ec1/5pTI079BxiVMQFjFhwyPnqvHHduKugY603tZgK
9MXkgz4VOqh1gKMDEcf6EswPvSynAvOdiyzorrL9iSmm90mtp1EtRYzig28q/FjHf9NcBWkt+xmj
vltF3SLFRGwxxrpxl4cg5pGUFrp5qpZ4smFxA8DLhDRUKrGptLDgBVOivff/9OGk9GG8WvKMgqUz
p6GZQ7t4FNPJYeCZJjSze8uqeNdAaStZGZu0plOqBxtsAXG7sdtB6TTBSHm15jum1gr7mPew//k7
XX65798BdXnfCv5u01EFe4byl+oqrpbptIueAYwFW8Ka+8tPSQYyTMmQoiTrCVj51wTIMCWMV8dE
IVMylUfxmjNqRCJVeNJtsEixIDSeXB6D+8OAlp5V91RPMWX2ixUjRYs2G2l/65egGhup6LTFwx6y
mYm5kQHLJ3DsxMDiEeUCIWrISw0OTsF7eR6op+WzdXhjdHTJ+tejyrDDBafTK+VzgBBaIXZtyyV0
tpuHtXPaV5HH/RbOrUVURj5LDR+hJAEIv1jhcA7hwcCc5q4uLIrs7vYcB36UBrf6mVmBtULkkioL
xzWhXxKvyG+bWyX45km723JSCkuyq+TYYoAL7Z6p2D4OBtN4s94hCanasSVpiPxOcbZ4yqwsqW5m
zr3UEYAKNirgISmWrnbrUVBoLUtF5K3t9UCnO/FSnKvIpMqtCYvpACYJZo41CpVgffl5NmY2jPPD
gEwcsBF+FABGU/88vvjc9YES7QtB3a4skkq7KajjqDg7Kj3NBZkJRAndyYsaB8kk0NLBbsl7ujaE
CaGU/bbQaSIaxhkCKuLoBnF/9PWAphzqiVn8u4ES/tojUkaJhq7cTRpOUMbNhBhcD6u23dL8QdO+
bUHPo7qi7nSw99lFYY6457661qnE9ojd9BirPubiUeDGzvTFwQ0Xp51dn2LgWrmCitDqnkNAyBNx
EjgD38+lNYViDtDgYJ72RZZ1+AXga0XYjNKFuQXOT7kFAhm2402hLF+cKalMPZAXuhnlt+tgQOZf
SioL7eso2Npx7YjIXozjXar/f9WjTR3WwTlbAMiuUJklfQNJqDUhlPmDi1KaoUJg02DLS2CYGR0v
mlNxBrXrB93q3l2O9X3RHGxbzOT60onV8jkJW8r2Q+MU72d3Lu6aVj1uL/MWn4uQyQYJAsRkbnDH
yQGVYFUI68LmU97Zk1BMkFisMgQRJkpwstc/6CDzmN0WpaQ2LktOqdrYVbQp4sbBvObr3MHUysxn
/McTlOSl4aHYxkrnOOk0A6knYl5L80s4E71+IF1HAugf7K/aMDoHgXNfOGeuUxeIBIWYhP1uszRZ
QRlqMYi/p/yB7FDGZNaq7LE1LVj3sWQ9qqOAmMdxi4v9mqtiMHBHR6gQk398Fmhb4K49XJNq4PPH
wXRF708KUIU2RccQJIAu/FZIRqLU/6IOx38AAbsWlHv1xN9PMNUInM+XKJtfY7jtQdBtwTXIg/Ki
Tu20WNAVAv8B1Crsuhdc3MMew8FemxpueTKQukbcnXFEdJ0e6+TQNwZ0xp3I+kFH8D4Xr9FinTDo
4acfY8fSLlFGPBykDt+x3McmqnU3x91z1IbeFmDYqnsb0radRX76kpZUWrZFNP4nM2Rh+UlPplqt
NwKwDX4ZSQwsy4HSwUhYpfC2m45Q7v0ZYLaUsmi1MKJJAgJPHFrLBFkJOESLByMXyEVOI0Onm0y7
o56yBhYAsS3HGdbTGNw2Y5vNC33BxcPHiI/bZtJHCE8JnelqnRzcyFPRzn2f0vVtUKx6PYvRKOU7
oueZGDIZj09N9K1H5aflsrpTOaw9fm6ncHyDq2ljUuMlI6+/k7a2waWGiDPv+oP9KpCKOxlBVmoY
tXc38MKLrIWvHTO6zXvj8oOts+RzZvBsCuI9cZPqPGK5wirBgQrMUQ3V+oz8RZSKO+9K1/38Zgcb
fmfV2vapBGKmNtPANYT42PAIRIGYvaReqN3LFm8a3mjeao85wbLQ8H8haA8BybbvN13GoPvJUFGl
CJxxlm6m05VKs/BZVw8GEGvh/zMyAxsabVvQc2LsunsyXJQD04mgO8i1cIDZ2X0SqqEILmikdfvk
KaHPapkPhATiXe7DcSUSA4FQD4Igq3ItWBsRlixqj7YsVBsykiYoVBBwoxIdW5eS3F3iKUPMfKUf
oXKTGSosuDNHDBxSFI+yvVAL0uvhLh8GKKO9BtEjqv9lPJJPOrViCP4QtFmV92uXQ49tlUHEV9rE
MpcubW1Hps6JFmBdVdqRR809Hr0QeHXhnyjKm3A6TvJ+OHzFTz4M8ELO3261qaRwMnyTTAdBD7Mb
gMkha9InBIZ5scTDLe9OgAU83uMeoOueWk2b32g80O7SmkpfBwnpqQU41pH5AzSRWsINSPDILsJH
cOCnrCmcWwcUGSiA8ewgemYjfnPTduzqWsFPi7araet/NIqJcE07yBag9nUB1cCyeM3A3s1tvvEw
0YTDK6rOV9QBoQZKkElNIAuLwJqGA1OxWK/jt1E/4U5J4nsd32Di8FpJeipoA7NfOGM9mOOh1Dh1
WK5JUwlnDil2tU2NUUU9XPk1FZPG85Zlz95jPgcN7sT0SaNtmK53lJWUEOkY+kEn687VKGYihluz
FKoDuSfj4mUhXrHtVJl0W+ns1ys4yn0zjkAefxavmSJ74nYZ0rIxweLY2fL1I/hpjzaDhLHU0004
BhHrS0MAHJLhFb9+I5khOIZ4UnMsqxQSk54/Q24tixomr6qkflntAJneQThAoTHu24OfOPJ0E9aS
pZWqwFXSiBB5JDRi7LKavcyCCbKwWafrlKuWzNJgC0Jn9zGxEbP/ERDFtqRi58QcCaYsky1YLFRU
oikIbphKaH2XVtwEvHSj95TU1VT8alNee9vH9fOOvOANSq5jWpEnBT93TtwZUHhan14xhbqhPdsK
TkZxCaQ7duUJu420/bxd1C7skLfCsiLMKuVPMlItFI9LTYOyi8tZLs2oN3KHRR8iRa85OqFvpEAg
ElvSCHgpPB6MO6qfUmzC4Cud8fBJTVICLFgaaR3SlCBPl9YR5HcpxPoJ5qsIGtgyQ2Dx2n5Iw7Fm
Iv3WkD+sttzEnDw/SAvlIrxAQekz6PbcLtJfX+IAf/i/yg2cD9sux7Fwt2E1pyTR/POImSh4pMYo
oi/Sm2YAlROtkvysj67UuyJwEWjDyoyUbBqRVZwMsx+/LDbPdlq9g7375wixPn3rYzkDyCD+vnWJ
VEOrb2cnlSnl/mt5+v5H6m95ZPCr8vzx9ZC4XRVds4O9HjFkxtQZpI+vEROI90YazXPKvcofsqC+
wZh4ZJC9Kfo75vMd+9R0tQ/dKKVAeOn1fw48MCeqoTW7yElisJEaBBfIQiHzUKexecTPL5VTuPiN
7EmcfgVO2mGNCY4Hi6bkG5W+//+Kq0nm8F6atN5FJZRdQ+NgwHHIvZIU83Jih4StJuRpvbGOnX/b
ImV4wJxeU26EWvYK55t7uAAMTu9dPLAznKkQjgNxws2ULfe/6PtsyDOTXIyURCiq3bNf7HCjsJXp
alKG3wGqDON/QJ0ecp2qj2lJeGrxf4bQWoZaK1ps5d/68nEVj5kw6TusTAtiS9p1e93O1BwBizjZ
nvDUJWTaQmouxXhdo1r3d6Ug87TDbGTnFro5zosmjiE9Tn/opuJ5MT/8rSQytJtn0e8Xn6YDZiVk
MDXxG5YgYJ5GFncLocqjIApNpaV/aIOVBG4fSUfKx+veRXJ448R7vS3AN004THYkpNs9cuEHimlg
VP5IBWHikccqncWSK+AE7nim/M8hpqkQOeIJ9BbcAy9DzmQyq5vJF2oAXrP9gFd02VuroHp7KXpB
cRHOgv0jPvtUTSkFEzlwD5RwM842bMDR9iUqVxg4DOQawsMJmZ9Pw2K64uCvVf2CaaOm9S4Ah41G
v8MYEZxOovmnUHJE8p/3AfAjrxeQkt16fvLo+pXXEj7oEfmzX/LutnXoi2KX5o4ZbS0ZgbKPar82
mOiBSgqYC5LXrlrBfAnnSIaXmufLXMkM5mrLPs13HMJ++RkjhcVIgt2df+f/JZWiPR2XPzQO19RA
ZQ6EuzJVSuv2ctRYnjhvZytIWxcc/0pf76LdwxV98ZUJqZsf0fraOdUcbx9nHHA+yRTmw7gcwsJy
8nfeIQ9BcH4njzLotzr3Bh7HwFcHiY9uA2ZzRb6JW07syMmfSnY+SLP5A0Sutb/ksEqYPlFow5dI
LFOUKfbWzrY+u3dHCn9l9sxtF8iaaHhqL6fLEazuoQnLzMYWZuyH+AjKKww8wQuZlusRGoGuvPBI
qbfsKro+g+TougrFhiIJN+yhGrEMg33V7jlp+bFblaNRmlCoVIrCQwXhwIvgdSSR7QH1OOTAHwO8
ALCKcK5feyPlzBGdr9wZOHpjPDV2kBzvzXuMFj8QN1WCgyaY9COWLNwdjoahblLywuScNzJLtN2J
EkvGuaP3T41pzaURWwSx408j3R45ImCGI/meSjQlWTp/GDzwY8Zb9TyQWpjduh6YeVlLkcU3ivdQ
he7kbNoyNIlFYxqHvFGbLprVrynE08R+5yxeuuZ7ytdu+FnzNae4yR46H3BD0ydoI04FK/s72nU1
iI5y/sisW6XipcqydV4jOI55ttV2dwdTSj1x1rf+hiMS0N8dRZj5wN02sYzNqP6UxO2imwEMrEw8
aJoVxCzEAoSf5klctSCKV0viixLyJ8PJgUVCQmpVvC+g1MYWXdL5dj5U0XjcayrIpbKbyIa+r0GY
JX/WwDvgJ5hyGTvqXVy8ho1Jod+WWjmrYRKenYB3fQJYeYvk1ZKG1N27IdysEv8J0INTWxS+Z74B
MhPMYRvRNmvWmSWdlYhodPVmmZ86c2GVxI/2Y1xC6or65QAuYhD1Y95LNv5gqlBkXMAGu0au4RdK
SDgQ9QUuaxAdcq3QhSSTNj08KIoBWSVmzkPLzKBbV8bBwBv2ZgvxM64Eok/0afXW/3BLIXE6dmeN
BF83a/FN2BwCed4dHbnQf88rstqtgJKkcIf0y9YJC8j4tyNGAuN3ALAnyv8hzSSAkC+Gc2u7Ykhn
lnm5BnWxhmSebIf+UDx3cLLwxXf8KOBBpwV2Z5TZ9oCHaWK42XHK/SbZ1rh3oadnaDaNlKySqlJP
1JVwFVNuPxFStXheTQiK3CMuJbay2ghPp8WeYJxnKfpx2PicQO3jvinfnT6GIlQsNUI5gZX1JHdC
fSADQFxRjtfRe578bbO729vSCCxF3jYqHwm+6pjoigSYEtdq1e0e2oBbfkpnVO7s4QEPGU85tP0B
k1UEVN3W1SjPkT0HrX5b2v7MO/asvFk6tPL0Bx4EHVIqnAxOPYeZdtv9dZb0n2vVGPC3bDXBSZ1W
NzE2JeKo4E7iD95cg/Be12Br/ZEl+ghCQbqWXTkwACx+zi8tgNyRWeJM3icdDZsUm7O9k9wYEmOk
B1IGPSIiVCitRFM/7ctVFE48L3HXfQdroSkZG0H3nbQMsD70ce9odGDUbPMWmV5i4TOogrthiDWI
KCiH5T2+MHGPkv4LvL7ka3o2hZorkSh+WKTtFGAyXhh38EI/aS9wKwFOsqmMrwEyhhKoBkEMwabU
x+PgfVqlbJDWvAzIxuYia5Pj8jfXlJd6XB88qiYs800FxZ4jSxVCLmff8oOmV099BVOcfYeTosLO
IF4vIVKsF0pjULNoxcHOMQvl43CUp6IQl7dlE8CUYEJt1I0eoSMVEdlQGuK5vC43/+2fAxymZ4qf
5MhxAPek5tIq6nAAQ9LHPbPmVR5W36n+OH2CTLYkLm3zOBA1GI6fv88E97HzunNquYr5rB5Q+0va
oqXTQD1kPN6H7zb+yn02TSAQxGSDhIuMn9CPAkdYSNfxP4DXF1fE8TGRg+KgM8pxeTYYdCXiexiy
Tjbf7CRBVGofWWV+l4UG+5TsaBNRqcsgOsqYHfvVX3Az+p93bELxA4J6LUZq3KDayTUjAY/wsrzB
7nWARxUNT1SAwjYRUA9Qrc5V0pD9MQLXDt6P9cmdXMOuZ++aFAhw04twWmsyMH3jghPG3kIOG411
DvJHmMt1Nm583yOzrwBX5UQQlmLHQsFW9aqA7ocD+T+U91cos+6ZNGaCV/cSil9vGxgJUjlQvoQ5
7sUh5jV92jfYtfj6NgBOhMBxf5bJr+lTZWxXebS5IDYG8RTRcnqPP0K7/lIfAKuh9jA4ef/XJ/mM
YprELYFu51lkMbjdVxaublPt7a8Zn9ze+i4DVbSpEXHBiVXf1MnDdOAQ5BQQsQMARe29+RAnUnhY
e9t/odEbVe5cGO4AG+GmBxjW0I3L+nBqRy533KJBizJJ9ysCSPLKf/sZfAYmUa4lWNejqE8WGviB
tkbKhqm/5dUVyQkespG4tmzKfM+WiWg9Gieym+rw81nlpq9PY3YikG7S8hrUd/e3LF3CgVzN8QUv
xGNUlCCffixMuqGzIgb4jH6ssR0OdMZshyDPE0jSWvXU18Z8cLaBgKy+oE9q4RZ5GB1WUKzSDv2c
89mNDCwM+u4oPQ41sdvp1Jr7e2jO3D1yY8+a5W0Ea1AaN2Lz1kCyPSKyXLsUbkBfJaGx40JrQcXs
zgPOrVnIugSefyBRFxuI6Qa69PqX1sz78YY4nxiu0uQJC6ifvhEG+3EZDl678D/aL9TEuCTDfGBy
zQx9RnQi0xPpm7qfIRezcUxt6jF1dKEwj3Cb85SxflfEZo2qILRQeO1eSe9oAr4sV++9BxPInA7y
CGWkG0nC8E2mKgKdaecpOWYbdMKrqr9GeSmVrljNdlUpVCKibavYVDzyqhY1VpknGQvRRN/R9TkR
b7lqn6XqYXm6nxap39MeSifxBSFD1wzNb2dP+7bJPNThOFcJzVGYNwirt9SZMulD1/tZU2xK0Ynb
yYjCcMuosrD2CoYSd8AGCkc+FlZDooXmL7dXI2VjRkD8NPL1Zod7OfALGY67+Jh9xGhwkkAtuJlL
jxGVzw8Zpryl5Hxn3O+o82UZKt3+KARj+CBVwkvjUtYvrf1p+Wp0EDNxrdkGsjeJs639yfEfsEQ1
FesHdIsovugXzSquMcbfGTO9lOoyddlCIvExmYW+HKOr+urBkrwNMRB23fWPxLGh6c3wVN7cgcXX
ttp/iSAbY/bJlRa/FFS9KRBzYo/U9NxNITV/5oefLZMU84s0b03mXecC5EgTw0r7d7THYPF6L5TE
r/ZGC2oyiNTOvoxF6NwWCfoRXwtUT0GjQzt9FH2B5AhxFS3CYaZ+el/Io/Q7ZoHAq5HnViAb11di
5I5k2KYrYF/gvN0hDthp330c72VDloTzUOCa+XdyJj2QjzSmroDgTJlPo+AOWWEFW5R0SVcUqzCy
0bWShdGH4rk0MDyMGvLzPu/sL76cCGw2BvzNWrwl0Y0SyUzJF44qmhd7H3rSKZ3EOHAhbvE0Pe7k
+GpS305vMXF0tengkppSY1ZhQncqrxWDY2jQq2rXmjUo9bvWWZBOxx9IoXG7byuihYv6GDI+8pyG
1Vl8mzgnIYF7AlfiXlIgAp2oJ3X54JHTk+/S/LI4wA/lHZxEcxlafBB8M8bqp+Vufryo4jVUhRKo
tdm9WHebeRkG7Zz50eVqFRcJ8NvXKvXNnlNw/o2yKNiPNesGFaXKfFGK3z8jEPePAUYrpZCEfpAY
GtmRcVzJO+pOUJai0u1JjVaohoRRANdfJsOi7waXppetfrz0l3yEJaUVI/3vSlixqME+aPETCiu9
3zGkWI8V26G9R/exixc4Q6V+pmqg5AOSft/rf/orClYcJF8/6KjQkXR8a6mQBoRusUIWjIwaotP6
AKQ9mFBY22m2lIPI6KKncANNud1/YcYrKLwl/rKytheafqF/e40BIon+v+JRonvUGLVJIjKesxXg
WgCV6F3RtocnlJ9gwizEzKGNRM96RNc/KMnVd26iLJLOSJUv/NctsWMaaUcQf+Lt+acURYzzoR8v
IF7tGUlSdGDhwY4pAK4HIdiuTY9P9R+WgdBvsAjPBUvbUIK347zTEc/zADxxfAFojcGJUFP3vM2T
/Kl/pvTiOz75AofOTruhC+JkR9UQqD/95xm9h4wsX36yOk/UXqL6rnT9SBQfGn4JGLQQ4u7qQNOy
oVYl3iR+sauhWFS8Bc3FYkxn98kqqZDBhJn2utRLug436AgYN3El4YHaaQwzNRH0QJvlbZHXfeNx
XWG0Pg+qUmvjI/P8Uajy+ImPpbkQ6RH97q9Z1Ba9dgZczOF/42Lu+kez8sZ9HyRynienSJkaIPs2
hqVUIyOm24PJyWdFJSscvZCATSXSsnGdOKqSUapCqbwrrLPy2jYPHkRMlRkseuUo/2W3SukyAvQt
I18sdoIktri5aoehy//3LZ4SWoF1m5FQfEBhDAyI2NVvcmh0nx29syPMXMa9fuD1YuHD8cnJJ8uY
Bk/21lV5rUcRAsAsIomKvbH4sBlmsDeLvlWNSJGCtr3VOnQR9CJZse9qvhVZ+IizuZrm5rSgsV9N
DFOcllsrCuamdvdUWrQpbRDcs4jKVp7O/8jf8k2XrJdDHvV002QCSXGoXr1CH9M5TPGXgOzPAidv
UKz9DCTU0eQ1QMNN95Le49eoD6o3FRgLSmeUrZpywsA4wt0gbq+ViNFy9UhHIn7tx4pCBjIbx45P
FyY6aFk8fv+vVF5RTPdKmsYX3BCcgig11qS3l9tno0tBYG515z/P/5eTwvfkR6jy0qo5PFAKKVws
tj3l438k6gekCAdgwjuANpzxipviuiwt6MYgKvfa2PLrNEP4AYWORHUJegef7SLUOeWU0BGCkUDP
3y2xqszr7DrmznpnHuahnYZPSI3UqF2IVZvJB/N4RFbNeQwdusObmxxY4+l3SDoGGiGUM7HNSP+X
lqEG1GVBQU0bzhIz6/obARLHymEps1bCEslYKr8Ni5rC/fwNDQ21m8qTXV3F2OJm4JgvWlWNWDGy
oqEp2vUvgIE6EwYCu+eViKfWB2YqRg6S2D7ND8KrvdJvRfMlNVJEJq0BYVdIr1y/nditYPdUn7qL
RNzh7XAk9kWI6CzHObWSwuBbn2tooeDhNm/O9gVBdE81KaOXPXYyidAzUwb/wQvTK+meKtPxUVag
C2qHHwRCYEE+dJ9Q7XqYSscLqufvUh1HjcmixTTj70RrBAuE+pgobzbdngxEnLHYF5Ux34GmcuTQ
mkufZ2SUsZXv4N7V2GxlRVH54Nektsz8UpxKdHARCGv4NYi52B9i+a3cEyH6CNn+xfHY+tZtT1/T
aiOtB87Q3z5WhHD5F4b1oSL1UXL3jd2RiYiebqRLripo1k8HZ7p327c/O936tEDlrD0NsnOeUmdG
9vBs/QETQa0NBaz7ezD9lq+fExk3SK4LtR0ZODtk5PHYb98up5S7oU6eGILTVXsyRwl2hrovHiqx
iXltv2nv9vhvMZwzMy911cviHbUytmjSnS19pd/u3AgABBILjm8JjCLlW1T1eG91aeLgb1oRcNnT
RNOLwjL5GdAB2z7O05BOCxb2WcUy4rOz6o9E8eRyrdeA2fAePvL6vc1fbdEingbFxKTyYuxaurIT
eT+B59m8Yae1lldjSfIUzRu90plr1N7O4kxrSDkv602LWyhsLzAzHEXqtwQ+qXRZBNynw+ODoxhg
+nv/E5iXiTjl5TohKESgwYXypfhikL18MIRwEUrkDokuQaThBUQSEJ1YoB0H3VVbyHbLFPOIiGKg
ZiR01H1gf59ibzthkFPOXcbSIBSxnze+AOgm+pqbnedB3YcOh3ap+PWl1W7ah20qGFwxt/QdtjCO
pytO+tWBrtLvxijv8So1yy6DlTykKczeZaeo4s0c93YtftZMEcmrgUuAiUnhn2PeG9OnvMSOD380
BUjwfxP6Sp66KXYjSyyCP3B1T+T5GOXrDSNb1oVpMypHuCQVPewqNoUGgtZNgzfvcvQtAFSdvfr0
VqO66GCV0ZMC4lJl2CchTIoBQMwY0OTtQfD6iLzeW1RFMvpfAi2b002dw1N1Cg22kAzh5iaQ1Ufb
JbV8yzUgADRbUwWmb5glWcEDqigw1Jfmkzgxk72PxgDtnhgZkCtocdiqHQvRo6BnTqOCL4X65CTU
K+iYsXf5PP/1UWeUHcssI+fyTrQaidBklGKSbMqJgE+4bcs1vYCsopBytV4Ea3NCJvinQfuKh5FL
VAzBxt5cfEePALxmmfPa78RndCwl0tspfeANVysURWv/d3k60yATH7O6djPOJxGdAmReE9zbhcUm
yeetI+9/oBGsiBovIWGbTB5jzY6QawcfrO/DHDFiWFwjgQHEoEI+HvfS78RCzRKk/M/jReO8sZwH
BzpUO/f5DKDFoqJhsSoKJlVbxZdhj7bYqKH3g5JtqUcfw/kundFqnzLy0ryrM0lpdVtcHXKMPS9c
fJlfBYfh/K25fcVzQeg5rdG6BdAKF1wDKEwZhsN/1ksZ6pOX9pxfBxZr0s+HGSnx8/LoNtNiEjEd
zPwjiefYuRCA65FnqYHxAZ6OYid6z+DM5SLOb1lbnDpFVIMK+rFUhzomkwDsmsORZ6m87Nt4boO1
DXeGmCpkwRgmUDbxKcLS7oV2EPTmLe9inK6M5/yvl88bs5Df1vBkP9XRLoKgS269QfcKOnsqST7Q
pkiR0rfvh3XmmYrkDVTJ5TFHxpvZq9RrOwjlKZr/b5kBrHO4rIiL7iejYmJt/jV26SSYw6wS4YSO
LgE3/d+Ae6LSCC+EjMQihSQA+g01jgxckMtSMK7qCUEry6U3WEL5leXmzQc2NaeWxHhjENoXObdr
Se7Dt7pmefsC4qfPlgEprnYyDTFRTPQeiff4gbi1mdt/GM5ACJHmX86L8c0b52Z+PBcblSCmP+Si
ncgcjLvP8SF35zl5M3+0W0r5L3CfyCv2gVyf7IXhDQ9UOzfIanpARbDk/EmylMtX2OzLjnL+mrog
yZZLQvY2jenVXoLMzLwNLYjvE8gVKtGm9Z2jkEwOD4Gz3okNRopmQzwoRdhMM4+DlU1vIHLCzpY1
b1I+DrAVnytpZXMqLiPEn62+UO82k+JRS6vEIpUC3aw+UyjPOb9k2OWyxZrmgK4tJ1iNHs+ZwuUC
Lc/seUAEi9nFIDxcYgcqqoIRhRamO7q4yfQgL9oD5SYbVc/2OzLF6vO+eMYJHw64ydSU3yOQ4BfH
Y6oLJmZnvOiOAR8cDVim0pF4sRRvlw+H1RNhQYHDjDZpOK+aooe+XubMWAPumzDMscgXfo71o8xo
Tqb5uFjbZ7962zUQW4/TWxhGUa9rkH3EIGRT6sinxH1VOB31eQhiq1heRnbzjGrV3nBIex/evXCL
j8y6cInomGekQaNkGY/1BegtNTt2baLehIVnblwrU9kmDQA0bHatpmKhe7u9XGEXWmarKK8j+RMQ
5dzbhhH7GGc1JFSrePucMwqb1QuWLHnntOuQ7LlB31298LWtMoRMEbSDTCb70ijA2Q6KZSziX1b9
zIUdzJAoDu18NRVr6RKxGvo/d6s5wa70UwNjMr/zq37/yg3m4tTEe40jZ4R3+T7TPllunz0MSv55
xaHuHkusY4P8PC1g+07NdgunvD/vr2MI+LdfR5z8QKNm9XZ4QppTFsjBI8M8upg4ekPqVf4fzL9W
uRCb8qBm2cs/h5KaAMjZ8WYiH6dk0qc8i6OqGs+rb24v8Uub3/ew7p5B2ObXlK/b8wYKh+B9aQnZ
mdojCQ+E+RDZGrwkXCo/y798YzVBIAzdTk254BkWO4OAlb2CIlgrOdTg5Ddou9NW4b6gSxYEHcnt
liqHROyLYC9AHqeNxeBiAZdCv9JLQ2nealtdME/OPCMp0PzHqQH6bqYB1iazjxRkjsSluE2IE5cF
a6p5XgknokPR77WdfroZ1JC/YZr0Avwa6qWDS6sF6ehjHBoMDiC2YPRspMxp0yFSNOYhq0QmKnWJ
6FG3nDbMd1R3GRjz5WLhbfdiElONhwlOP2iCNNnXqIejcjLq6FzJF/Sq/JTePEt1Wgc1yjb6nVUS
01skc7wwjkfCWA4AJlvwn70lhpL9xZi76Fz3vdCQF7w1C9w350sKor+Sa99y4rfan1HfKLq9lH1F
8WQeBiCcBZaVHKUf2c3XIXIEJVWO/0lv4iDuYOeEsWau+p4mhcQobw/MCEbSmXC8fxdGWjGF2AGF
K+QzqsDENbnI/eKVxctgEZGnOXC10hrB80UmI+UBTOVR+z0w99hUs0F7JtH1FzLmGbx1pPMf03if
BxJCq+AQQb+8nOCE0oFJdO9n4IkrsNIfFosl3FpNPGa24GRqexPbnhAHU6ZQL4sBLa/2JtQsDKGF
zg2k3EOKLsQnfi2A8pU/OLlCD++cZrEYbp2D1TEvWBHEqNM0jLvbHYu4perJe9h9sByg9Raq3Lc4
BwiR0qeM6FniOtVcBLxz3Iwu80LsC8PCaE1W28Dcwql/ztBhZ+B2TyH9wi5hSaBtv80KiyCxXb8Q
GNZRH7tZhfAZ19qcW7XaniPVvDZkBh0Yq51aAunI8k+4f+6+U+FTamMU6o/M8RTHnNlEAon5inML
n1vt8ly6od2IZiWepCt8LqLH/m+4tVzgQvtqzX18j4L9xG+8fWcwDWq8eyPyH9V8qYKhz/txDPDi
tgdkYPoemDiS9s/nq8LCMVX7/A9XGWBkFPLtt9//CClyGDps2OUBYt/kGq6yaeXkfxMpWIrJHp+e
b4rvOFAWyT+/FQcpLMXGbqz7oNIL50cwWsiHrMuvTBComZaYciLO9tQkNC35OGGH7rI8jZgx6gAY
kLA4TUA4wl7XS6rfxuBVtbvxFsheLTtP4igthz2ZK54SNsIQ/Lsvah7DmO7nV8tUaD2FRhv/5/9M
z+iZBE2JY4l84qM0nkVxD0qBQrYfZbCfyPByBBEcOlP6hBek3NyDiNt8dDjrktsasIMJtOb7MQGj
a3Xplgqj5pPAziZoUHz9ceVN+Lcy+6bhGfp9pIfQShWv3orY4StbaEqMwfp8E9qVxHmPaVSRQMYR
i8g2sQ4hBBo2ytdCqmOcKRJ+OCZWNnOFHayztxqQhrITr4/MIsrEBYCGylUYZYI4bvppKVvQsmkh
YLEcZltDhV3NjiIsVWHwkrhAj1PAdcbWM/90bZ9RgcRvd9pjcbHnX+bN2HZFzJ+Z2WCaRtC5FLGj
Suca3lSZlP5QyF2kmKL6gkg4Poo/HXQWbBwKYzZ004/EF9fjhb8xucMlIw6mR6hoP5ASim5aOOfX
eQ1gRAv6Sysiw3U3oKpl7FYPXP1I449qU9/E8U+fL+mDZoQ4zF/07p6Vwhzlcbzp6bJTozWEA1T2
3BA+8pVdjEromJX7RmQJWE0J3Yna4ee/m2YuEM6fGZSPFeg7tzQEl4Zj4Ot+K64bLmuAogXk2wAD
LT0akSPoF/p4JIRrY62S6ccpEeoGXDCkickgKErllefIxE9FqJExC4lgQkdThNe9B5ZBz9z5TevN
ACta1WRFAaXkzTZOpvo2Mre6ajgWYyPib42P97Z3ltXwXJAClCiHRMH5PEkcdj3ylJ2IbnyqVr6c
z8ffawgVi8vf1OKUlVF/35/hlDcuWVxUwHb11TEREfyL4ALbiP64LgVGXV522HQ3S9pfPLKw0CWL
o+xtcen+jlSlULQAT+tTkD9au/l0s/3hHdmhBdd/0nAhjE1c/f6BqiGZN2YVAEvzKqS6I91AUPGB
lsZsNRFmCFVov9tPL+7QvR2nguFSyJXHMoYcVrZK42zoIp9ouaosVTmtLndzSrX32yd6M5qhiBlY
04iNuZ7ttwZV7lrNwYkohL9pYCAi+cMWjFNhQMPxSE5XvCaLnd8MfPRBE+vFAyvReLiX7TJ/MWL7
vnpzj4G7BtBCC6fN4j2KwsAnHlDHvmJ/lPlrBzmxxHfPNvrnvFA28Tab0rzhP90dhQIuhVILaKo9
wxiGLsYy4ECcvlJQ1yN3iR3QQYLFtwevS5LwFSAWCc1rrRMT/cS/2aZw4Z+2Ony1OkASWv3pMQWt
UTKMOfRugZpUNvn1+FhMtX29MiYvQGNTT3mwPAzMLKZjFELqeHcHbh6m2i+qzX0ans0id4J+K3BE
p52hdUbMNSuGeZ3XoO5fpxXsx7e6xoBk/L9Z4vWx14uUEao1wuHgfUFBwPm4roNeXcD3luhWRxQ5
4BKJa0tdhkXxjenKVedw6hWncBJSbtrPPlBckHp/2t214gl5f1SoRZIcVGN3Jxn2VifTYeQgBg16
w+TFo2Q51wucY/TJwfTKIg35+2mdxlDYPghyBwIaMEnXwBg7dRzoTnGrPP7tQXdk1SH8PLWG0/S/
CGkmhkDwW62QNiW1zQl8DEZ4YUKUe4XVaBTpLIhvERdTgJRKebaakV1XVEnNi4nsN1EYc9DLryoj
kBRGqIDWiotl8GOOIgvfyULTG9LFZWGE1UUl8ptkvveo/kb4JbEXYSgF+8NRXJXVUK9N3aajC2Q5
jp8grMpgojj4LG8ttX6RP5xnDciX2CVj0R5cXcmh+F6mOL78JX4yPplr108s24Zr+EfpMpELkqjM
rckwqeHSMHClwuV1NuMa/wtk4LDqOT+Qvwn0W61KEsKHoQENDBEj1l1wQkc6BElNJhaUZjEwR7gC
hXZhn3y7u8RI5W6CX167wJS2ExG8HxDbZth64gbgFW86ZI3IAQ1xXJJ+aGkLuiUjQMRyBnrWe34I
Dv3b3M3cfSK4J7/HcsZZQukjjYxZMdcQRaqyo7/mubuh16aDGPtjXoTFy2ep09RG8045IGtHkoQy
0Jq5AyP/Ih/8u9AVCOxwtzAPMpgGgmM5cWgtiTkP5w0FpBq3KPE6adz5kfmtmTLZGpl41P1WYkHV
J9XEe5pzdnCEkpheXKea3BWlxrdZlIirW2trzQ4zlIZDnOzP1afsKuZOwFVlR77oDiJ1GiBIqPNo
7lSjr1QPPJeEsFDgZoafW+mEwn2L6Yqq9F4ZB27N8MxwAVKtjE4Pj7F7ixNR/rj+nf2bMoV7JOgP
z5sWKwNCm+p09DLYNlTj6He39AbcL0pRjgXJWm/EG6yeGnyjMCdxXhbYg9NuRv6Du9nQLH3FLNlN
x6HRZF3XN8zstibjE8kJO4qXhkiVM4AG0RGY9wWbHxjnX0IxntXrBzGLaMH5EfJ+RyPMg0hfd0Gf
TKutF6hW6aIE1GsDXyIMvuQUIfZNQAUuXWpViy7tmzeFfUyicLHtUgCZY0x0cigL1i5+crHVyKfO
JbOeNwagL13VmWbJHkiEgeRkm0TPDBRqtigUk27iFKCOq3wsFiuz5HXXy+LePIARoBQg+dFlXd/r
ESL59qvVIro5YWOasU/dDutmkkDeRBVzhKnp+UeguK3uFTQYzQ0DuPxiDk17gHXf2dBxg5jlBKAR
oX/WaLn25MEkno5bs14HOkuDNnsDgy4aGVLyBRl6pbtACQ/5CqBwpKBVZqjDdZ3FFf27dp6rg6wL
tj7YFqDxouoJOojC95qWy7EIFwxewiwbjqs7uEMVIUEdu1L1Zm4f9cMxIWafF3lxMKwMJ9dDjntq
y5TK9YnDel0wip9tVLO2dmB7ytl4Q0sdhQAehCJJckUMtM38PpNy2gNZAW6Oi++HaOn63VLsqehs
VtyOOu6cvMrW1gBjGXegzIR1VJBzyIbHBJDLkCdZ5lhCW4ZVpSnC9y2ELRl8/yrk6PVzRcQhGHNT
FhU+g2ouuUNq0O0a2rP/2nLIEgB41McUv7Y5cvC7ZPtLNwlnNJRylI5xPMPEUylG6K4jXdqDkYRA
TW1fpEy0Z5w41qm8jvjm9xsbN+jMvDlxPV1maW6MyC7fbwkidyGot10xJFlo1581PM4b1z1yKkbS
7MHUw9MDF48HJi7ORdXkCmJXqAwSzDzkm4/b3nMX+zvBxQRYz7R1Qjl/vpW6n70mAxUHgiUZ4x5r
okS+GUKHpqNWhrFa0U+BqjFcmM9HB3PBLntMPyyjythEJZBmao8G+GJ2o/VNNRh9R+vmxbQvcwoW
l/2Mpfq9GQgiFicDbmBUx6WlcBxGmIb2lRlLmqkU56tZgRXQvEFDf03uL7IvcE4xe+d9IrwASeME
bknKgeXXdn0Zd619ynI4V/wWqlOxn6q5c8D1d8wBma1Hh/S+09tBh2NW/whpg72GP8HVac0i1YtF
BBgtgIXGfZL+JNW//8oyfDJUVXnvM1lKry3+ICVs2XXbStu4IPZOOZYttw9Xx460Ww0V6z94VyPk
JhpWM6jQzgj9BMIqkJKTkNzqxcDHOUgNmozFq8RYcezzZtW/vl8ljMY7uvqHrzTE2sll6zGZHEQC
WIlEAkgWcrNZq7lYmW4m93x2syU7TNX3L8cadGr6TBdvrAyTMlOmOT1MAxahRnmFnsYu82q2PZDu
eqBsBmxgub5yA7dpvRE8sSwHD8XmZtrH6GXKucjIez2sAcGUyizOgi4O84R1Ej0U60Y3q4FMpWy5
I4KmAu5CGpKCqSiwvx68fkedkBrytssrpZLSSmyQ0aEO69xuTXaEvXC/xYGGunpQLYrbSFe2xVSq
4MIDNUOHBljYFIFSD+2m7hw4+BI9Ev3/gPUTGJV9bHD/yuVrKnkXCI/EUl+QY59//H9hlnfSLXlB
YZydoS7YXo7lhywgUogvKnzAxu7fNfhv/wW5uVFuk0tG3/GFNbaM8UamAM40gM0IPcFj0MGKD464
tbY5SuLAsjIGhba580+ajKAyV3jhal3GZl2odSByKWjuF9OzoFvTMk824dgv4I1gdbEKJLjvfMgp
mzeHM+dlcxkiRZIbeCw6owfwTMGUjHGnDGqeDG3VYBgyz7wmuhZu1bLnEDKH8QK/ncVeoADAseeB
HrUjkxi3i9Bgr29YmwnrTkzz2XQogSNqJAvjjsosdElPXFX2mV3IJNCOQdk8LM5OEoikDRFTCNA5
fjfL67bmG8ufNyutmZukTIPyOpPc8xyIyXD8ZhBZtTX68cG3w8VnBF0D2hZhGIFmx8WHsbIehjvd
wSYQrtRHByTNk45IzThT/XSqVOqUwDR28/bATMhalyrd2lzjwzmkV6keLj/EuOAKC7m8Tfo4aGzg
Vau8JGa1klBEuH4ku+DLO5NB65cOEjDf/rDNqstjBAmQ80O18TO2VWELYkeUjY/VEQhtJHCQhcUm
pni0eMDa+7vMBcG19qKmruasHsNuOJg8DwSa35eRlERzaEojG68RaUCJPg3V+pPkwU3KilrNZv3P
1xjic+7Qo8FWALSfD8AiH3QlKE+PsQhCyf56/Fc5tqyy64xZAfDEchsxmwIQa8/v7Vs9CLhWpjws
+a69b5WkboAfv6EfylrJGPaiBz6dsv5Ucc1SrCvDRkjymXBMGkbmalPJstvCIuxMzOGJWiGydLnm
tO3tPJh0C73Tl/u2s243gubOaufZbWbikYhv1sCY8w2xjsyOzQsB4Dd+d7gBRV65Uutg05V/Fbpo
+MIThbC6HCjYLv5PyMowfLisyZ2ImlZRIzmMe7/FY13oM5FgBmNoTWxCMXj7Be8ZD1iQ/EETAQyp
j/FwEu1welxSHJtYqWg0E1T1mNVWt62B3tTcq4bBM6Wu2NnlbcDdbCinZwklHvmJl357nwQw12Ks
VUKF6VS/2X25zpyXRDt1aSHGotj7rmQy425/SRK8fmqzMu65cZTrxd8ssEbeUZHglZxgAGda5r9/
JZ+CgY9Dxnp3OSqYeHb5AEfzjMch1XyxhDriCzkt2/waBqoWxvTXWwmyK+HYFXcwCdDazC0VyZ03
hovH1imoIWjvxLEezlsqQm0q0hscSdtGrHHNTtXZAs4ZGE7tNtRTX14+0DhYRHI1bPgLd8CeRE9o
rMICyp6fU+ej4xfR9Amv/gtKhjHgh5A1AFt3Z2fij5IlzA+HjdHBU085Yt+d4GfIJAL2UKZ5Rs/a
GwfSkFdo3dUE18LY78gDuxdkoTrN6lQmqJPAtHuEoUT+/yvqlgN/Vq/R2KBez9cVoOaTAqNRIkuI
t9Obirqzc2d8mEq5eCoXCMQibs90kukfZtVF9oLsUgzeB4A0OgSKO/bjjRGihS8szTzWyRPFdmQZ
R+thTfrGbJHrdvSrWm0/h4cJEZrVDKIYGiTYVNk3R0LoEdNtAtMmEB21YV0Gb1DqsBP//zLXHs2U
t9i+XsUkIcyBKVX7HGiGoTareF7mDBbN5eq02gSsEAtSOyjZZ8WCxpNP4m+SdzTZclR5kmZzPLnw
FOp5/4RTFa9ylSGMS/4KgIs/HG9bfihkhtd+0SdkvevsDwUADZLZg1gbohvFRyrXAOikxNjLaueb
ZHDffWiHMOjYaoabYsK/3gq6Hcn0ExuaPgQ3vZpkrMoKMYU/5V3fhOI4KX3x8WrOpkvtcgUXKnNp
I5/VwPAixAKw1RN/EEb1SVp/LszXgpBY8urtOTOg2eOacJe1tvkjAH1uDErTQDuUmBgnKbXFRc7I
24ebfrwfgFHnxn1N0pRbkJ4tPAEW/BxuY2g7rscJa7URTMCN6K2VQCNcRs4tqrltaK0nAFrqqt5d
N3/lN+fEmSDN5DvnKCihlobbM3mFkzdi7gwYITbDxVqs9Sk0LkVB0UngDWT0y0xp4HxWE9Zm1FGs
/y/SGRYklyZq7oRValIen08tURf9ioXaE9u1rNDZr8EpeWMf2snCw348LjoS2kjih7FhCQ/Rbvux
hRHPVrEFy63VsW6FJ9I77SDmLflTZSIYClXMt9JtJ3DINtuJHOaEGREGQaKV/AxTQgf9Ju8dqHLW
JDeyxSfiAODaP+fmWxFR4kaktwGIrWo1OXVIM7mywaSqpyRW92W6RWXvO/CH42uQAtLmQym8siwq
+Y9fVdr8gt4WnPq5Ut+tBIooCAleMFKvnMXzMc8+GdTJzsLt9qMJQqx5RCN4BCkxCCOlD8A7v60l
YWiwfMWm3GeD3B0ku7ZEigYL+YTrMxtfSSDWEwgUKCfBfueKRMpdfrhlV5ObfzZWQfIYc/IILvVL
cWwf+Aw60fTCkE2Ue6mD7MTM7o3+g0pwXvVJDywKl5P0Xp9mdnRYP4uQnsHEdk9kPi6g+g90BVv4
ff5+ufshk7EG5VANAx/YGYIXt/lRXBpXyWRG9HGWGQtrv9WhWHrbheFZVJk/cydaqn71d5zB8W6r
OFV0aH8GzgqZX7OSCt3vRMjwE4vKTCgONhJnfmRChm57AQZl64aJyNtlxSRaq/zS5upQZM/37E42
ow6cw6xH7ZeZLmYoyYjdxMwTfL5ms6pHoxkyrbMpiFRidOiWZ6W1J3/Sjd+tiKuSqwk8WwONHPHX
mWi30LeOlCg3DplA2+eQwifp3EuH1+p7LOVTkKnhah4cH6yQEgXqxxf0u3bgxWrmWHUL0eXKsT0m
rKquxM2txGIlzQ2FOu8QXvGyFzV00TrgNEImD1WsAktNkc7rObVZsh+3RhiU5TnvaKN5I4gPIWhk
GOMWnL7+x1hZwpWKEfM5W43BBN6p6DGYZTrAkJvv/nTh7DRuNaNIKwDQRLMheX0cVQ3sTp2/kYWC
kte5g8Av2IitDyupFqetryj6qPujqFDYpFHnEX5bGDwdQBXjXORBua2fQeihU58rCuG/U8N/Ac2h
d6LGTUJZVgzfsImzqKo2nKj+sS0kGKSPy5PEbHiUqYkU7iYHOPR4b9N8WY4tQNztisp0WQ7xXYex
3XWgWSqls7S3dGkLn2vRxcOgIiGNLrkGdkIHnnWUZ7djesnoSkM9HVVeojoqlqCIDyfF9EB4mAaa
17bijYIXwoWo+3oKy//hR28HBXtD3zq6h8RuhDFUapfBR09MSeQUvpln8muqfkHkGv1YnoeFGb6p
/uaI93b/2ioDuE4SJjsGYuj0+5RBbXKNJyJKblx9KU+IDomq2Y3bznszzMFp45r3PFn09bazpU+A
U+YbSLu27Hj8lheT9upfBn9IBAxjogBZVexziAvsPJ+dbi2m1Ctg5PiRRkkkVoK+VJWUOIAb6Kv3
QBqTvQPLkZhsWJzcJ0QhuaGC21yEtmPVkujyS+8i5PndKWtfU9kaKxGefGVyS56yO3x8fW1XK6J8
CfHo4ep5ODpLYdpnzj6z+QeSSjO3jKjbHLoybI/YQYCRoulVasjQfzEKx5nQ8DWAifbaJ3EaG64K
RKVxud6VKLg26dwMStIcTs+glPDxYHzTzz7T88eBRgIqAwyp9XvbYQjTabcSEXtqBuTyTQ2DTyvE
AmQnPQUNFmhjryftTjzC4McNpEc9Hh7Tg8MJBPIGFkjIOW3lfwSqEXVca7WCdTIxi2j46WQ9GZ+1
N8m0qY1HN4yH4dzpeTlLBuXZeyhmbXxXCUSldQ8H/r+dcLmOBqZfVlIsSYl8Nd4Z1ZcYIPUq7AkD
Dp3A3opH9hQFDM8dgxNUzt9y+xH3RmWFLb0d2PIX+LFFkocek8f4POPTWFeVF6+X4JrAfQSeZswd
/eISveTBVmPkxoMt5IpR/GWC/DusJfGc8jAKDOBcYFl/i9XqA5TRPkc39HMvEq3xGN/XT9NQ03X1
Im7au/IKdBdUXrXRMEw/GXjCoHQ37UrdJDFdoSxkbaDvIt5RUHdGhmYaLc6/sRlL/eVthI7/neNf
vBnK1//5C83q+xRXjE0h+UVuB+jiJrKADR/P+rXGczgzoCex9LneNKvkWLoL1xKCCUFKXr/q0cwB
HOwRbhLS0y3kheU8MtSChWmuzxafmzNnBplCPtXG8h2kjdFf6B9H/kzL1Tx+xZOnfKJZM7hxUzms
VSF5MuvJgFFJ1eAEi6C/xvmkDIMTg57wnpLveuT6LooyoaLOjPa9z/n0Twm8MpzzWmthxXsiIRpG
RWf5g3XKcvgeT1VTHHK0U1wT55Yypx0bZn0yOfi0UuLLg93+pMY7Qj7hc2uOer7v1I/FxBwI4n2/
k96YtPN99vUfWOh3pOz5VlsryYZYrBo8r+KIl5Fmb2n9HYoLDIIzYY+ynVaynV9Z9/E65twqESVq
mhFhIwgNr48uDE49FkxgGGFeb7WSjrItBhvxtqhxBpk6fvKR3DaQs+lL1KLimMRyyyzORGqwHqkZ
UHO8oMYcsgkjnsmKm2qUWLlK5QsNyOiahF6o1FJ7COYLyn08p2cNdeRYhNjo1LJqkFlXttxTlGq6
Aq2X5zTn6RhmM5YF4lUyenKfnO2du0+I5waaIzqcKMuSRRg0M1nlsaeM8l5uWw+zaYu1apFm4KOk
WAPY2VmR1Wo3zV0oq/Ncgg/JvxsaTROQP8zgnY8UYwk9aKg2foqsHljQyu1Vo3JxPL+8TwaPTMFb
YDuoVolK39QBKbWQP8V0C5juCq1zoLcM5YP7T4QNgHC9vzSAXJLAZm9cO49eGotNH+ka+E61giGk
b5+vL9D9bonFHivDcinyj+iLX2vv6jFA2Oz4ftQwzkC889HtFpl3Dadytef35sE/EEVfrDL/nZsm
W0hhMz3GZ8vK/48SSqyi4Y8B2TZ4Je1Ae5ad9z7sTUIz8cJa7H3/1FrzmPOWK55X8rDsJV9ctOE0
R9CBOQoJhqhTLEXAy6wcIXL8DOZpNGUx5xF0n2zylA/M2SFFkAI4GR6cfzaqv+W8ukhyQjMQCBYb
zDyMjTBQWfrAUTxYj4N9U94m7+c53igmVfCSUYcLjLQhQkqZNu+iiWqsoidDerYdmlKNKMMtRP+r
b9IvWujremsqriigzSELGwljhhD9bE8BG5J5bzBxI/+MbESIj0tQcCMYq4zF7P8oxKda5lUpc+bo
m/7ZzUdLx3WO6IWIcxrREuVNeBMab8UwppDL7CLroJG0RBXurOxmozFh8BIR0a5nSOx3ZmyQZV2b
2uvVAmBjr2SVS+lO3IGwYt8k9OPzP/EE40lovqOdUAIT4baYfsYmSRoxzWtUpybB2XFzY/MhmvJX
X6ZWeCtSY/G0kMYoao1yIUpIqQNS4IUzYC7aChRhv3gWi3NosTEyXiQox2XBf80xUwbsihnfPRuC
SSqVrldf0oe0WFB4CKfIsULYXuW2yD+pN6wx5UsmHoI3HqwQLYTKJSj9tq16onNeh/WW+AKh6ye1
uS9NiwUhnoosONv6FCru0kTU7X7B2exLngaCqfBhUTlurKPXiKzVeYcGzPxmH+62/zLK8CnECdAV
OKpXzaNInN+bU4+2b+3FD2kJwypMll8YxynUySqAxqa+MzRuXRxY12/F2wudpjaNJweyC6AD8w4n
82GLRW0lH7i2YulnyI7Gzy0Kjhduh4/tgzeL5rdBREbMAZDn7IkpGO+rT9QgQX5W0bpmMheGA5oa
h1jIzPdIeBQAhs65ocK/LCqginpTyvBBQY/QAiOxmJoew6jrSDGnzOBSe+eaqpUcsfjp5esZzxNS
SCqjsXYiJ0E1VuPqmxE0RducBH0SP/4pYD70y1LIffu0D6GyyxylLNT5iv1GP2ZHd5jVP4nAd+62
Nu70m9zwASsUIAecugcyTuMBbpBEtxwMx2bNSoD0TW0lf8WgP0tztpGuCBet/CC9NmvbagZjEtVR
aoIZBXXhw4/2XPX5Cw1hzGNGYkhMGshhfjFvlvVIMy8WQmyozmM3UbmMeU5AVzaRka+CpifaZXpN
iZAT/XPgXkLMCTuhB32dpYHuowc45Iz5P5z66h3Hyw2PXj98gojCII0DPJjNU9drpMmZ/a8TDcH8
AXS3/tRPQZPSvgC+eprU3f1w9hNaWB0wksdpYJvD0md2IzJ94uPHJPiOo0LLAT3oDJr5fzM4vUuF
oyO3iPzumZ63C+pnw9VYSvoRGBtbtlB2BbXTnsoko3Z9PaJSFKQaICXOeQAmkYkMetzTcc+kQgIE
KRdPgZfjSvOCyGQ1pYolktbxkynM4FxNGOQSmbpqiPVzMvCsRfjeFdchPf3rhCNJcK7L1hUEU0LC
LdGTDZncwQZhw3cwKBdPC9LD6trabZgNUajx6/rljjgVxDydFPRz/KsY0Fo4gswBJFc2YZ4PDM5p
T4HD5E5RJ6vwYDhRkBDxQ2MocqxZqDRvOO0+Y+91FmtEppRqjGtqIw2RWZeARmWZnnsa/0cMjz6n
PGj0JDXSuDN6rrMSJWaGkZGSOchUdOH1aUW3vE+YdGkuuVt59uXC/cNAx7rLw5K92DjyK3oLZKnX
/4eja6lwzSJIwzjSJFefmlLa/cUrdQO/Ah4sYfE37YWuqLWr37hVmVd1szHR8ZQBEkWTlliGNA7t
Otyp4+I362qT0Y9mhBfqGDSfBMpn4wu5RMnlh8z1sG6ZQlk/1tpdYjqrnWc9D2pZANzKqD9YxIJA
FIVIwK0vRt3BHKayZ+J+kqE0QiuYem5taweazNg0PpNMgRlJ6y2m6q1I3rKkQb3juzY8zw4Tb3Cv
aH3WXr/5+eIvb87bAV4cvt5pCP/eYhRi23ryixOle74M+ZGHNKt3APxmlNdhadkxpacPS4ygtFor
GSdYbMRvWtTagfIHtdCt1/Y2SS5fExjTRFw7eZl+VedieuLrvfLTgDnkr7DK59VzMYFe63VKNKw+
lEK8AefNz9ynxpDEqUwTni6w3lndxXsWCKojSGd/h51K9mlhOnE8tUm9OkqSDI5v68f5zjwpn/9N
ivWy7bs70R9rd+aXghsu7+tdm2SX5kVsa2eHXnfklSBdnIiHgydI4qOnOe5j9g1zAkJhgEYBD7f2
I6byInphohryhOBB3X34rcYywkQqLXX+7VuBsWzVAZnT4FbNoBk/hqRdNY9XNz2bH29NQwRR/iSF
ADo6E06GxfbUHZPu+Sgen3A690pQEAFdrs1bYaWDYBeLOHuH8sHNsTNA2Jhn41e0PpeteI9UbXq8
K29UrzsoVb0jFLOOoOsXdnQYkMtvcFBRZysmLgxbWmEZM0vs6m12kptbaLiY+ZNkKFebnGhXaTyo
X9vEMWzyrK6YvBulti31SVbSwKoFaJDBKILTf68MIyIsI+BdBxYhEJpFNyDJifuS8PNFUIPAVjHG
Em3kgZDQsx/ye5p2cvQ4EAHhucxqRXWxlbUndLXHmnTmgmmnmX2NsklkoUYRwWNUW97b3gYzjqoc
35Yb4HXraZ1PNIg2gJJ+XYejh3El/brQ4nTlbYto3duFho+zluH0Pdwo7FTa6tnIfKyicZ1u6Swu
+87qE8u/yXJoSnUTglP70hWPcx1fHQKSgtHRaUbApjPxOB4bk57N/2DfZth9bjrSB3NHAaNhIG8f
uec1tIO17IdU8GUWReJHakzO6VCQ/k1lvo7YHxZ73J2NctFp4b0Pqw22i3xWs+xMPsbS7YEsvej0
TgutOkBJUxqbIMyWX12frXjzMbdRP73TnUEcWq1a0ewV3FwtCwwYfZKhHLYVcTr6GH3YG5n2N96l
ErRVGOCkoZ3dOrbBVUreBj9yonkT4/hWnJPX3U0g+Czd6BIrCWDfanKpkDoGAf4K0618r0r7u+2r
CAUamlxam7Pip0sh7dwai+neTXKUMrTK3CL3C7z7Wn6ThB105JVle2P5GVro3Yb0CvxlQFdHz1U+
HgTmG/YiyVr5LiGGEJekGPEpY2uGo0Kdm90Mq1XhtkEnyZrftirfpgVlrhw6+OUgMc9lU+Jlos6w
kfl7f4Ww10XFgve/NsxuMAiCmcmx1kQAOri3PlkEEHStkWk8DAhOIPX86qFTz6+gIZx7l4e0B0II
X6ccTeyOTtyA4bMsjeS9/W8zSqKSl4m2o9gReC3FJqWd9yH/bIrtCHQOim+5KBS5hJLcBfrB/fAD
vFgcaKgamA3m0pKlL2PeekKMadlqcXJG2yuwah3TeEC6xX6aPbEiTelU8gOY6fTtBaMHIRR735gq
NlqmwgraCOWBpS4t3Vj6E+IGLDZJrmSyJMGZkbilifl3fNLbc04EiRHdlpngEefn8ebMMTaoMKFg
UDIpTebWNFPOq/e5oWh67Xr1V5pzogw9wsmpIcYodVwM6b3c/7ZrJoYV3VIvzerHLW8oXCSflG7/
nIOh0CJ1UW1Ud/5ovfEaZ4K/dpT/Y78ygiW/o4ZrguVzu32SucyEj8pzCenkifXfuVZ77fX9AGOT
zmE4q5pCzBp/v7Ev+5RR74hx5QfYFEItDATQzTwQA1/g5aPhj2ephIoRB5K6SFKvKdisn8bUSGkK
2L4H2jyk0/5b0YXMFUqTH8Id9YYXR0h5TGsdhhSplP5QI+YR65TqsA5jyzwh4fTnJSzltMmzOVnT
Rzie3SbgRnLB8xZmfpaNeB2bd6FO/9CqqfkdnLdk4ggBYVABlRl2J9MuPcSTrFY6v+mjVpHCFqWp
ruO63dc/TdD3b4iaAcSWG+4DwstN4wkJuehOWzUSIx57m7XsaTN/ETWTST3rnZwAu7YckIr+6xdT
6PM3/0imhbgiGVaH2pObtomKm/hfXqU9r7sxzGw3EWKCznekLxK286wo/XACNgEFY/ZgfWGy6akr
Nfy9uE0rx5sIdlIM3883H9Mn1tFH9hs/WHpw6y1qxGYVKrBYnWMtu7ayZXJ1yMTLm7CMrBUPjpTy
FUYTtvi7iBvJ9givt6BHzF1wO2g228EKC0QYWLq6rPjvZGrkwoqiSwNP4B0sB/+On7/ohVk+qPql
9VeJfvJgwUp3XZP/uptZwaHVJIc9M59MyiTbBasKgGvZw268LxSxr/JMI4UiMqcaXLgtsBcUiDqI
B0/Bn8IdZZfWJtrqTrE5jFsr/2zgqS5+XZcovTsT3wZpULY2ZH//GspKLf+YFK+JTKqGM/Onf3Fk
dqF80F/KIfGOtqutm4v+jZEQiJZPK31GidQK5S7yYs5hdmk2Y9P08tPepfQwAce4FZGHmd7g8JDx
nv8ujHJ4Bnj5AKcjqrYwFQrqisOrgtEIjUnYs15H8BEBoKLFFGJVKt55Dc3aKOwG/ql5eo6oq/Ze
LIG0DrwXfLuGxOVwd0anRXWaGpicWQ+rUhFThLtk4jqk7zNMScZvN9YF9kOSly03XJf4c3LLgcD/
qcd0zmzS5xRqZm3fX9+1RaKwmdZMtPUx+ltEdF0P5mgyGMY6mwPDqEG3wQ4Rxw8hhnYg9ZHAY2CC
pCJJquUu1a9OPCOgKPN22skKSG0kalIeqliPU6QLOEHRruljK2wjdL84WP/h45PhfiV9xR9U99sy
czlgr18oK6fdsD1qslzBKVxyM1N5X5LksjtI8rg6tR2icAwOzcZ8htnw7tYSCFwMjnRS6r6UQPws
iBhfJajAqsOPpx4BRufwlAaw8TPos0lJs5MAaCLXQ84Yt7aN2/EEDXCAJvkKXXntP1mb+p5F+XSn
TXp46zu0yiBAqpYbremwPyRqI0H5gUGGvyJUfjV94T5cbxoXBZ2LdpVaRvfN7gxf/ZBjMAxv3a+4
1j1AGbUQOxz/HliYwmPa/rdLyT1Q0EB2cl7yw2w1vvvnJAJNCFcUufFCWBZhHmUK/JihUMXW5jU5
+ihkikA+e7PZa71UzJ3CyWbiXsWyyDuDxZHg+I2oofIEn0v5PLh3RRsqz8nHvHGBZH+9VF1NX//t
pW9s3Vdaa5ISKRGY3upwJ4k/0xZnMYYNEgvbKc/cZpmsyN3S+njYYWh+GfeE/lnTn4RMhGHYs8eC
LQqaoqL/74u9QhlwX/XvyuyUxQWBex4kxxehAmjRHIGlX4Tt959yCDgH5tJxp3NuJt7tP4AoSuXw
o6AvYEQJyDHPNiRpe1mocVRF8NNX/mcp079Rp/2BffO1tPJSnqFBErPaEaGfUtFjPNrBuFiytEMv
tlmYebil7G24cDA0Ees2lcmHSI/hKTW608heMfOCbVqAVtQyqgMr7ljpk1XV5s7eDLinZxeZ45UV
Few4IEgP8jw5wgc8iKpe4TKRvlAgiNdHqhb1e6llwyCVzHGcqLTrJ3T4cqQZla3yCGqK4HbJL25p
mYttGmA25cPaJvlHLKVXGyuqj22NVcmx824luamPexWtoX43fFW1AOejLCwMODbstOrYeEarmywy
b3NExSVyG4bD2mzLiE3wGtANnSihcFn3zwCI77lrBzC2Bqy54z7nSmj6YV38ZE/XomqH48v0cXyI
v3YDj29GzXjkp/tTzBMMNR42shVytx+Y6QnNL8RtA5jgeqnMLficbV7Ij3YYeVuMklbLhfj+fw3l
xLESj1FyiRIQNG23Dy39lxNRutZGtEUzLz3DcYUDOuFlukd57QhBaVJOcdMHSN1aDUOKwCHsLjn/
ZibVudrbc0nhfeypRE4UUQpKn8Ud6befQhfyPMirGBwzcLOU5dPzS2+dqUo++ZC/FBAbwg94SF9k
lBMZbrTHyWz1Qzbq7oQ+5wHrPUOa0BuvK/Q4vXGv9EBN6nCWE63kJ9zGG5HxqUHUPT6J6TRrxMcY
zXD85JKlPM08xNWWQuqd1ECm0QmAH93bt7nKGhVHxzPZHYgUyjrdMHcBCif9bW9R+F0BfJTo8JgC
i3af7N5m8DuwUyrD0C8PQrM8jV7x0/9uVbheKXQZiNmi9pK3UfGZR6kd3defbYBktv0arUmU9f/L
uIgHoEOt91ea6bUb4AtZLIPsQvjtW+ErVeL2MnEGR+CyxjikVCFT37QXvzFlFEV7Vuw/gd/ENhbK
RCOR/CGpNx9jv5ElBfsqP7IoMqsM1cSiDRz7H0/iMMRh0HM1q1VJs8xQwO7qJdPRot/y9//6LkFt
Nr49FIF/HIXfqZcWgKLd02OJAaxxqKft8+t41Psf+BdPfDBL2USubO81baehhhNuzVNnhSyJSFq5
GYI9BkJWw73y5IJQUpRl3FMpEqNEFh43JSNqf20SaBv7vIKPY+Y/cTI8lm6ofVnPJvR1fOlSxQkh
h4WA0nuOOtZd+H118fjM6JrvUEunwfIpsC73Ffq/djblXVrYC2qUAX3SKYYAZGX8JS4zFQbcQLco
vIpktaoRmAvghJGP5wkl9hfEhfo+rt0SzWhT0NqX8phtzOvJZNyGm5nqUE2A4QWC/H62CzA9kXe4
lS+nMXBUFH5USNdD6CcIgILR1KcVscTf5WrhxfrCWIG2j2uZs4TDKURYjSLDYea742lotn+nnce6
9pJb2rIdw1Ex9R5e4mAH84xLG4Ck2SB2lWN/DZSFjDagkjCHc2tzm/Ht2fsSRLKy7cfUuphJrF5w
c+cn9KzpAk//jvBI1L4h95B5OtXwoB4KE8pEIpGbCcAFqMqz/JZ9Cw36QY7XlxyP2SgfKLUxEhtS
SFknfV8yOUVWr6/qXfjHL5Gb1lIck9n+YY5sOQxvYoC5fQkH9JxwTyesCXLLhC9SEwmbZNTvDJZU
6Syx2FKpM+Woc/jqplBRv5r1jLukS+2LqEP+L5llhyFQaXXLrvHvYSCmSWwvqJ8P/sYtSG3cUnv7
7igP9ZvZbqSySBPaltuLvTC1mTmhkI1o0o0EREPLSGJf0JoF50peArup6zamOpjjIhGQeJo0dBmG
sCT2GkLHFsYxiyjEcz8ttzSe4QOfcqz431o6+RXj615fprhclAgYpZ1EHW/5rm6SlESdPQoQeXPn
ndKVCmOgXGtbIfP9vhVaUsMKB80Tuca4n+mvMKAihXahxj1JvMUicVyjuneB4PIaEopxe08peVNM
XuSQMFi48BWjC7+QJdgE0PIcC1Seh8aMYUcz+RkXewiGFBpH4ETeKOgiULPBY8QF2Qlw48HyifNG
n2rWaK8TVkNGmvDmB1611sDUBPBfPQ+m5L1SoxLG6tmTXwrnYWVjmcTK60uMCZTAathtOJ27Tmex
/iutXL4mbB04/5xuNtGHRUDLffIc0Hf+3SYlR5GhGx0hBMI3jejudgp09WzZQwxR2goo4nCAf7lx
oWoHLmSjIRhLiqti/HLWRwSvsu4JaNwk6Pmn7vOutMk13Ke152XbLw+mDrGV9Wnb3uHEtFPBn3PG
nZ0s/mJz3fg0zLAEXaFe50QDb+GlbQ3AMeos0JbJp/Pa0MACfeU7xkVZSZPg0lrrfOkacgbajCiq
wdBb1RQZZryp27jzO0YjO+TB+jTDORCLztWGk78Q16JpjBrByQkUT6YX/THGyG/5Vcce6+ZrnnVH
4daP4hsvJPpQsXkFhPexLyXsOHTt0KoG2Okl0T4Pc5yjsNctl1QDnCxeQEt+MvyExA/QPlHZ4exm
5EdMAIg50PJVFFpn273ewktHadnxbYlf/A+e1uVboc8JiUQq5rYkB8u2iUlu8tqVIPplMcSfR0K+
L9qjIXK84D6E0UNxTvG4SEye0qhV+OVmwEuG2iLjFevQ0K+VoHhEnLOUbnyfF1XjGzr/bF/s2JBW
F1sbJkOUklazUEM+C8hdYSIIgvtTKfT4h4WKAk04WZ7lfIOGpq3hq+bdRT8Y/k4gyB8vjhtvj7JD
h/V7/omNkBjOA02D9x0gcJn89PN/47J7J4UtsqdxtET3QjUf8tMuTZ0zG9zEdWpuMd1ZuVmH/+1K
7XNKhUbPBjYxVyOWRSuZNyGBlqWOIRj2aBq08HOlP1UV9KFnSuYkhG7V89v1v+fqPA/LSvlvvRXL
n1Fvwh2yDi9BUezO7snV6BFnSiUafdX+5WQ7br4IcZ28jPmmsdw4zybKHJec8pvncTyqtqv1rI72
cRmpbsE1q6z8FO9goevU8pTMJYb3CHMUiEoij7XGLNJ002z6ImJ0IhwGAUi52usS5WwMKR1PVFIC
vL2z4rBcGNWvDA80uVSG8btvCbyaSlCis1+3TVy9SKRu63Rx67lfVqEiiasdrtxXSEYCIyWMWF+y
zHcjlprRt9VVNzJhPXzMkaEdcEHJfykOXW0e/I3aev/D8ZXvKzMHVEUeKje/mWXr9+2/PExpVfIE
idGCrnBA20TcP03690e/Zut2DUE6ZrpZRQGMu+ts6mfahYMg9UT8kzDCB+peIDZQ9dt0+AcYnHDY
fxuISM1t0qGZsS3+pjn9EySk6x+2ThERQssh6aHZZqAVwr1gWXeLnYDca2wf6WJUiqbbJxZ6ighC
RUPIz5VV9gYcoAakWxz14zrQuRiCTKI41AGQp4S3FO0zYl6P1QkNBO9/poCwQ8HRHoWygJmlshF0
gRtoiloOffWnePU8BAO0b2GBh4XtigYcqGD8WoBT2hI2hDOtYT5RRWX3ZyJX/nFXTljI4go204D7
Kbxd8m5L8SFn5LqLOH8g7xm6EP7MBdoAaDLjAbYtytJTUC2i25pKmlC20Sk4ITnmJU9oxR3WDYLM
YA8NrMgxCmYRs01oQyVux/Mem7IkSmivl0trD7p99OPU/UgVzNop1D5z4BzminF3kLuHoAdjVzbI
UJlHKy3h4XdfOzNJYnXMVxjKwx4NXeA6X+M3GOA6EvUBUTMQAhzbTorG/UWZdchEqI3KBKLpUT0V
vdFWnzeRcGg3PTp1H91+SDyKcq2rPcNCQfasao6SP1J01eV1QUyEWHYz2PSfEFCmzJCpLL0cg/O7
kOUpFsrzoE1+EyhVmL28eSqTV9mydPNvTyoHNmv4XLd+TUIg+FGin7fKRqF8ogEuzUKLSkEeKdyo
bAUpC08mP5ovQE2fQhw9o9jA2DK/RyfcSNHDIZRBkSfJHvJ6b8ARZcc6uK1hDtWUpUxHnSmFlsX0
jC8La+On7E9L797yVRBtsAqmOCYWluZ8Bg4DUboveIm4NDmW6NWybSkYaxRLArMIHrgKhJyPku+t
MY9MByQRB6rAkCLshPVze5rhoU7xFQofDmYAJKBTwn38XB3oswSlkU/yoEpUj13UxohhF4rfuHV8
TUVtgDKDLutd2jTnJVWuKi0Gjccyca0duWAg9C9fAjiG3Wsh7elS9B55lkgpWqVdQELsGUPzoB9k
mFCB5dITukc4UyMCNfgLow9262lpdoPFCbZzCnnYgMdEyB9akj2whKBv6q4szShUhYpU3S1TMNsF
+NLUdu//j1DjgOHJkcqG7Tq6RalZjSYFd1hhLDR+ZqMJmvve2SQ8Uej+kn2L5uUsOdTIb68mxW/S
6Vabc9u0xtH7Do09lQoN25ZuXzhnRMOSKeXjjXGlikRc/mlfigzKjRBfh0voGgBbgUAL9Z0kydU5
67Eu5DLTCS0HzF1P7xdjbXSevrWJtWEf4BNs8OtYnYTOpYDlxnzzXKNLebC6BvmgybBH7XmSZnhe
iyyFP0Y0A8IHkLFXb/viDVWcaqRh3pCwc4lO7q/hP6LryxPLdCCt5eH6MMD0aqikXUiqCozy8U3S
rFxA7DPEBVL0X7/UNQsdcvC+O8W46PEdhyB+99PHetwcJHYlFNyMOoA1F6CGl6lA1xS990ApxetU
USKHji1bQtJ9IYjpvOMhlru4mnt/un/5lAet6sdYQsl4hkt/4hDRG0mhzvwQ26/HP0DeK0v0dT/Y
ViDKkEkFS7QUdMHEAPtG7wCofz9H6rge7j8m4KEEiegawV4OVEktCqKecA6lKjdrWzBe5S/A6zLG
w2uXxu9Yuyl5mhwdDM0pXJBS3Ydto23DXnWx/VV7Ykc7HMqJeSEFeK2NrCxC2+/yejfA5AyX1+p4
TrFItZZZFlODixCNJ0qAp7QiryOohKlFl8KG3vJmY/lV9MTwzdfeu2AQt5H5zHa9lSw49tXxFScu
/6VasfwlKtDpZEZWR0uqTq4y+Oe6+MMB6PTYq1fUdgRhYxlePjZPlWs1eo+qQG7mVpfxNcJrTmVp
V/nY8OClD3+0EdBTVPES0bs/h9KG9VCQMqAeQuMXk80rmfFX0kSWv+G/BsjjME1dQvXadtvMqInG
uoutyOtGZtdKuxG4aqrSPRYR8QdtBznxU5ovn+7hRWo9N9JAPA+29uDmE4vb0g8u83L6SWZvSVrU
wXPOD8J8+SrDhMvpca6+BDpLQKkUIgbucoSPi73KFnH8rJdpjIVUt3u27wJ1UeSlkusch/msArrx
Mw3MWpNac1fjRxhnuW2ineKyGCObNJ13xiYdw0SJveynJuC+37Vj63LoTZ/yEOHhUQ7TtvMy9o1D
JbHLjKx/cJqTqxU4zN1scKK/skFGoA4xsIDUNyJ0VKpe3tOpU0VVtQRAt+6Zf7mFyqA2bHBTWZQ/
bRehs02luD5bNoR05KPYGPqFirbHzPM9e9LMFkkbH2swsnc89kLXwNXHGMMPgMxCaxgSBPFBdHZ5
6Ct1E0Kkxk4DwSxzB/zuFWm/NhCN4T/Pg1rkW8lVE4QYD35ssCziQowtsMa6SFZv2Hw89GGDpZoT
HzoZJ5bVaF+Kmq/UGAfdmM8m0zCJQkbRnsEmC88fm27dLq0GCMYvgrKRSljHGpAizm0g1RUd0hAf
f/h8r0dHsFBGNXLpWUp5zCiLZmgaoWjVIfqMjxglLcfVEIcDykzIRYfO88PAUzjd0ZEOlDdqLnDI
tKp9r+V0Il0r9FwA5ihoaYb9Y3W4uA9P3m+egnawDeSp/77eN2Iez6HbJKGrSP1wJD/kQ4fA++1g
5caJ/eBqYSgREPwBNpfNJ8Qvf9CzNXGRM7Yi0865iXQ+dvtnAVOtcyW2osQAnGXQXO+al676BfTZ
2fkbFTJD1fNZSi/9ujOLpqf4eOASvzyIGfnMC39iMnmriuLPDb7M6NX/Gy0kqc6M5HxIqMwif4eQ
0dQn/tVxcimLzV8nWeys74A/OXTPUIdFjs/ODpBdaeqnlsnA+lGq3LvLYBVa/7emwI1GWMhGq8rC
lVVefgaRBhkJafmmrQ1e/iXyunxir3TpMQq51OPxTSPlHvEJTs20P+w+QoyPuYdhE3KWGE8twh12
PQdp8FIu5egUgfyoyGaKJpZOGGKuqVGI0sqSsCmlzVV1YgfoHnqHfVUdfd+GON/3OluL04/449Ss
Yn9in162E9VAVRSwR1/8amKC0IbMwf4kvoOtfz6IVmvb2L9vbMZT/R+SWQhwqXvRbSB2Y+iey0DF
+SLs2yPS6hCkuqGy9UpwBd3zivcPpSrvcEiFJPwBFTD0z9mcLH4sVH1sNmbFHuY9br65w2ou77eI
veb561m/ZfXep6LE6ore4fS3XOhsU+1bYtvh1JeRqP4uXMsP/0KZFwtcoQ0YFcVLOxkLK7ezQvCw
P9w6TrifViJ7TyD2Zhu4d8nAo2V5+o3iU1Mniwbo36/AV0yldsy6qpgneBc1SNDQhWCnHXRshMS6
d8JiRp+etN7I/+ACwQBpMHtkxShfhp8mQYTe18gal4hzERFEk5sIchxgt2zXkHunihTIbMU5uOvp
W5g8gygcPzgCUB8OEUcw6ybv05k8Ig2WOSO18wU8UUhoifhuojeUDcKLf6kMinaVbkFNH79udubt
eTJiBNA1lxbofBzQjPRXlLeLNklAMi3d8N9SA2XmyotuqcOsBOmhz9rafRBgCMHCJia1HfGWrC9W
A3rVxUGWzIah4yWoa4Q0Sk7vQ8U6WdKxSCMQENZunXdRibwnw44wgkF2q1FFR0D4AuKrCAcqFmLp
+l+a7tNAJknipVMkC8Fcodbbp/tauasTZVaWIifd4XhWi3yxaYJohSitwZ4f0asq0+MfMPw1SmrN
uysYurvlUsMabHda030sI5qbkzdIy5OyoVXvsqGHs2mYTy9/VTyFeDk9/gzxo36nWdPi/RJPiEQ0
TFBRG3O7KM49akjILJK+RMF9vxLDGeKetV8TjmTxL04mLWd8deSUttcL/SN3/3iiUsFirzraFlQE
XXfS/MNrQcvD+41QJwbuwJSAVmYPRPUEUC3dsy4ovOKm8uw6/YF8LVxYX+AUTyIUoOCGQzEXG/4J
vWuvjA2K+M9MRtp2VjfNIBNb/D0YstN7xHmBPaIauwq2sITiPq4OXTua5GCLolqLKYj7GsnrMFIR
NNBEbX1XhM/SzvNLkk69rGUF4xSz6hCbtu2DqkZEXjAxKnHB70bWL9n2hnxnhzHrStYopVeu1zJS
Qnrjmdy5xQ2Nv6A0Xw15AqdJZ33aOWwilJDVHOXWjJTkL/OhJNVZ+Q4wuI/7H1utOyHED0SKZRJA
bJjJCH4BIlSffz4jy8HXo33/2dGuRE9V0X+wthxC4WtHODqPXyCKts87L+BO6fOCxyZVRAnFgeaE
F8ELVw+BnQyLxSTWYzfhOX3oDGiSWksOrnPqafNStsVDM3fO0/MPB4+nfPn6RPQdhSyvy6DWwdco
JnBOLZLlvBAtfOEuny7AtYee6IkawtyXH33YT7zKvNouNkDEGEbjapHoj6x8drmPMXMywIa5WoO+
YDLoT87dUuXn9f180K2a2bb5EH37arBreE+uM7nuP4u2hdE1r8+eeEZaUpiO/Xc75bEwJOoL0Ajf
8HirqKf5rFIuTytzEh61d2ZPKNNTTlz/Uzikpr3neUCSpS8g0GIOD8TX2bH2bYty+sNZAk04Ml9F
EPCjha6hLfQ0daoxks8vr1GFGJqeqkkH/WC+Y6W0tCsDCUoFjybQomOdx3N9sUFDJpwmhOmI65Cb
BcjCQ0MUR2lyvsM37cDbR4TcurgQQfCex7lIAbW7kRQTjirmoa1PDxN8sCGbRDvIe8W22XL2CmJ/
FzRZ2kHg1h68v0V/9ZBDp/hjZItmaOW9w2+eGKpAIDuuVPSSlIHbbfdhNDZvxp6mZ3a3W4Kz68yI
lYjQgzWl99t3628vAINOXkYB7RSCaxRshKnDoCPLOqc7NRB8mziZYp7SBIPqgjWprP2duZ+Ujihr
/m2ckzVTr63tqybxCCapkYB5/K02/kyNN1yx878xPw6sWei0JgpXSMwE4vhfStC1nFBXsrv/HxEz
b5E0FNQqcReDcFACbVd9SuPWQlKc26GIHzPHSryo912uVFrQo6TK8fsFY6Y0/RSMWVVwLR6wcBlD
NFhfSBmHTD676v4rDWoXg11QZ71/JTFl2NURAnYdpM7rRlWZqoN9/4LDPfM4yQ7PNp6beE84bs/D
1jyYczMtvZLpbw0TAraE7T176US1p/tomFcYdBOQstOeZWv0pxGSzt9LXA/AFS3m8ZYVGq2CX2ly
gefUqYO8M05XTsGeOlQCZabTnyVINbU57NR9zsFvWp/IaI3emOEu5qKriqiCcdkd167lLW1kfWFp
fNMCC2t20nq+erzBdZMlcr1FkLkzxBP8rROBoNn3JdaUGXnrhBiRnlBgypV4SagYzFT8HFHVgE5C
OQC8ZxZOoC3LiDAEkGj1RDgulGoMoU0QrV0S4EXKUM8tDdOEVDFSTiOnEuvHEMrbpG6pLKsQB4gX
3a2mEB4j0UZhUfmztpiKby+P5Cqow7PlsJ9eKRzzWx1zk8v7miIp2sx1cWGdC/Ix8eEU+GXy4tXh
u5N16gaRn7n/HDsd+mDnVp5wnFEZmL/A1g+DczeOpgieG5BQ2eGe8y5hr61KXlx7CRAnaW3xFADu
nkb/l0uW/QlCPIF9nkc5EU20ScbIcFpA6XPWJYgG5Y0GWywuUCm2z/5QiGx9eVPK1Jfv+07VNuuB
GU4YtpBePfNo7flhQvTwRTevOb+EhLD1YhP6xcqGgF/GZA8Q59itjwJcT7KmlEFF9VCodwZcDwp4
1cfZy+dTScpXvLiKMas/XI54Sw496xGJafIlfu3HCHS8Ic8NgGjRFDdkVOcU75+zoKietk8i0k24
pfCRVF+trjtrFegn1RvCOQyPYir3YEbkeyZeSnUIriG7XYTiJjJ3QriOpSls5R7MWIHUOLmoBNtG
M8YUuF0VWHcsiqw/w8YIK/ndZ88QkHSIrbxCeT8vD419uUIze65xmfhggBsTbYALYN0KJ2t/TYNv
tC6kAqVRcXGkVAPxWhvj9j0DJwvtVDID9q7dshfwWUdLbRoE2iorUtkpZyLyORzZyQ6/TYKN8EYd
kR/iZ71w1uupUva+5YvCJoNtnnwFob/2gAecPNNa+dKSxCPuMhzXnqYn6dKexZKt5DTg2auMDPYY
B56Y/iRgy9PracGt1lpOAcPMmPRIGDO8ERpLJEYY+x+ZA9rUEu+glSzJQjb1SNj1d3KoI7BrMIEl
/LSKqUu273MSFUZP23q58teXUyes0bwvHsIHzgNCyqcZg+vd4vWY0/bTQgxyRyr2q12HIM8KeRH3
XO7UCEGy1XfjNHS2MqX0Jq3ecGlVOsnQoxozHamxpuVQID5x6MhwzhzSAG5eBAGmVaFVTDFQ9O7O
amQblHi+1Plv9yIf+uIc0zE+TRMUs0nMn7s+RzdIwL+j8bKU5szvYkI08VzSfoStlODekZL9trYE
v6bB+iqY+X4VnM0DjcFVXeDaOkC1KJQQgENPv1bWBPBPI94O3AJ5Lfr9pP2wiAO6yif9dPePFA8h
wMWjZveaC5Msg0LXW1nXCwG6q907HMP5jYOA9dfPFcGdckgGJRkE+qTrUXT/wDsTPFTaOreX8ZzW
End3++53Bzift1L/O81He+um1szl16q77su2s64JA1lqMF7sFuuQlKAPN8sQdMwzSMadZTBmmSM4
Ct7eYIILt/moiHgFePa8DhdZ/r/BPSscw377bQyrOXDRKpEtAfjlYP0EYcDsqbMEh1JMBxF4tqU6
jn7v0oaipaQ1dWn/Dcze9kwXwu+JP8aTvYO8m+4OqHlPcQa2CRp3LH+BR3QbbxCuXPq++w2NjR9q
4RDEqy9V4N1/wGksmIzc+ADmaEueVMRU3/ypGWXqm09xM5YPYqOwk0ztLrts1SJAUUIfiTo62rL1
gELQDz9E72Sy34GcEYul8/d9eotJM4fpeEAEqn7146bVVLZ44DYADolvfYgVsBcbH8wcXnt4SzCd
nFTENXpIaH9K74ZU6EzKt94Gufm3kAG6AsuWWn/F6domKBS5wPbonoYrKIhOat+dtxHHIzzSqzm2
f2UMq5zF8sOeyOVl+d5wrNITUZAiLo0dc/nejqIk0ztsyi1uVHdXnelJ6hpvon+Oq/ILB26KZnLi
EGE3w25hXbP1FhFGdtPtmbVdv7Jx45SmiaWHyfVHOTynaxZPnTdamSpk0g4XV2lKzDDKR0GQp6as
o4A4jREvMlfsGfB+7NWG59mP9+ZuM9SIwqPC6gEyAPz8zm7Sy3qwPAhWuTA8BRG+CpsUb6XufkTz
u8V1hSSFhVXj5RZ1d4B9UYuIfsfLjpDNIlgUKsbae/n7dD3BfsgjekZKI/0eu9mjbY974nTG/NQx
w6ZWbLauDGDfFml8TcwYF5rYwynfBMjXFjGvYTzBB7pVZ76++foie3Wo5JsUItDPGctnyzmtMUrm
LgAZ9eAIHihHV/LSkcTNf03CojDbRSpP8A046AnxB/5VWEFBel6avJOGpqW3MYiznQsSBu2f71li
OSrMRM37nz3z0Kd1lmlRrwOh8WTSF6TyNb+dqahJNvQecSxU3zMcSwkQ+f7LW6iE8pRCLjGo8Nu1
WryNgP0eOkqYlBuS/QU1GzmaVqfH35G2F5KFmsEDFQYRLThx6zY+JfB+dzfmibMz6cjycfax1C+c
F96OjFQqCT4/bcqnlKeiTwHSakbrI5VI1BVt2r+JQQ8Uw4hPtrZQdEfz9E2b0VM/iJ1OEGEh4Tji
SDj4LG+GXDA4U896XFEC+dgmqD2UCHuXBLXdySaJslAhe52sUIPKFhhc+H9p6dvKibGcZ8pFA/Ui
zWFxq3I4aI/zpRE4xv37s9+hF5J7Z1tcEOSZfysxLI33H9SUdDhNqCGO9cax3KEtVSxlJrXi+oQJ
TVLTh1vilcenz13sQTIfZmp3PIyvwzoFXgrS4P7v6xkOohIOEnUFihcRA/rE74sZFvtmlhhsp2Fa
yiCwMmhU9QzZdoeAU/LVXnBbBHI2vrlBuOtlJwgOrhMGodPPbvFvjrUpu7/hwrvo/+MjlNC7DN+a
Achp5OjoIfJuVpzHcLzRnGWNPydqbbFNPGHUv4bau+4IUl8BzQ5htjdqKU+Xh+dKHNcLEftASuSm
6uVoPVhYLY6cjlr1PIn/AQQiNSsgM6Cy+/lbNKpSawFakWwdF5O73pDUFQ1Nc6+7nC03EAieWkcM
lF6jYC5t8XOhKPPKr2uxCFfBzRyS5s1tHcoqkB1FZ0wKViU2LVaa9bAlAsC6nPKbSlPZvu+G0sKY
Xnab1Z6L0uhmWvr8ay4XiZjF/+1Yk87+WgAaKRxFJD0SbDzNXqPxeQjgXce8Pp/VVMd/sqf9AlDP
Kgh4yqz2QGlygQslozWWDlr3sgqHzUb549ZU0eawRXzr8vPAV2f3jQontrN6kbuBF4dcTNKThXSU
DZsTjZtPYA5agg29iIkiT46B90xm8STxeiBYkuE/5Kvb6b77Hn8xkJUPId7T/6kgss3257kGS4lk
L2O/mcS6fYXngbVm4tktkGFug2F1Wx7iuEeC+XSe5iAIsFMXhDybDuKSO1putGSacOYvlOHzBezq
XFdqN9mmPA+66wJDI0e9lixPTb7hyizCdYU6W3SV3N7ezHXJxEsILqUuqvBO0/mQ+yxB6rBaCsqC
HiHbT+2rkD0krIKXhn979wgF41re6vfO//2hPKX5KoPbihkgRRttEfN4ZM1MfTWj8Xs9xE8wEoP4
Asjiwz0tw2gXZsYIeSLJeVjPantAqHxQBAZhQRx+q5As0wj3Am5DLA7PqnEDr5Q5WutlI0QISFkh
0r9NZzAmBLaB5R39svs7b89rXFDO7A6+Yngw7nTJGpb28NHptNkLPVSioBBD/NCV4UMPlbmlv/Ua
3WxrJ+SzCwA3AWacov+3sdFrkG1UmBjBkNpayDhg45Cegz6vAwqvWgYYaxZVhrjWKExCz7osUKL4
R7Lg6BExRjgE7s/voS1CmD48IWBD49mM0VRU3J62alXTBjXN/L4e0Q9IxnHL5NBUOM5uF6mNdHy5
t+WDZqsmj/ggslXcuYsMSVN0LinbAmhPU5Ox6OYZJ0bQwFcErLe3YCJl1mitXrIf8IIVMohIOUg9
hxh/dBCQVhqlZndYHn9t9aVKdFPf1cUFXlZXOKKNQm5CR8DO/vAeiEJLvANUOXR8VbBn0snTH1Fk
wImsezd3S5/FCjwrYNzMYEkPaZOujb/WXYW3cr5O6IlKxTb4ijYMry/PhWgB3E7/Y1EPA7W+qIOr
Sirv9Gp/XiR0E3stBJWyeKjpMwJ+/jLFh5loPc2d2g70Kdn7CWEwa8RWsfAVH5D9OswEz7W5Ll+l
t6Gxn8eAyIRfIz3tY1VIiUXZcmandm8HAlgCjLIzEbGhFVV/RjWrKOpQuo19hPX9a7092vnxsEZZ
TD646e/4IFEO4zn1eq/j3jeTndvcUQBdzXKxHmGwP+FPBpz4buTygz7zLrjy/6lk2e8eIUeTKkVL
HUuqghE2eR8mdgaWqQlD/PD/7HzpQWz3csauOC+z4NLNlFyFTV2jv3hgzkyVm/Tvesrehb9RMUud
V2NVF0TlQljhye+mVSC4GOlP9AJkFnQfhHPXYG4nai5i7RHuvej4dAQqo07eikb6Wdc1INO2ckWu
DFVzPKzTugL4lMrLpdGLaziAEe3BeUozPhhiuaUt1KBFl2ZlNWAq1YQIMR6Wda4iMDhc1Wku6aH7
6U/9CY2TO4QgUIFng54ba867BSx2tOD+bzJFWkbTAv/+Va6P7thzPR++aSuhjCrXzT06aNzIMLQH
uQq/jnCVbqJyxxTxdSeOB6zABoniZnCmOU3Y/KLubAlK3OH2NUIyWPR+oI12WeLpWAh2ntXfdbeI
RpTPPT6X+d1pNs8ura7/V77uSFYCHHWA9u0WnCExBTU7pastMCV7QldkCA8BR1+uOpvQcb3aA2w2
1RrkmWwRSXduLEFlK2R8N4plpKDyS9HNY1Mil787wA9r0a4q/6dalEE5mNrMpPjgBspREkB6JnAs
WUXrAgVD1acG5b4WHknyPkjDCFRCXSL90QO/c7f3D4ysRhAckl4dozS7M9jYXl8KR8WjpMR/UBgc
xwnovcXBW754O9YQFjmRj/7lIN6EYn0I/04TgEAhlUdPk4VRl6t3DVfn2Clspm5+X1bGllbYfZ8Y
tteIprlxdVMBLYHaSzEKiukT703/t5Ls8mSdymQWn8oV+FQkiOtfp7umA2MaQPJxNW3fmlXmavQ8
4giNixJIq6o0qIE6WnL7NofGv7V8CDjL+xbPGB0Y8GRLcPGawZ8O0ntkIOMVEs2UrqDXXkruL/7Q
d+ijTDbrhUFf37v1lfzQ5o8htBc6RBH7EipzJFSy3fSYllA9NMH2q2KyGstZuCpyaCly2qKF3q5W
NSbZo90X6YLX6alkJePB7jXMl51R7jk+CoOxNchGIWnRnI3jmHyUptrUGl2ntF3+KQa16AgVeXH0
xjz96aIn9XXjzd2pWndGLCEUYBJFBa6BdG8/pHdosWxUdYsIwLB5RvJhFTcylvfe6GuZ+IVQTsmU
ukB52Ta9l3MWwvCz3wB2xZWXUgsupmLJGVfbLfFuUoBZL2qjUOr8ELw4yT6rSy0ZQilhdLfK2GEL
CAfQQsZGzCTcUyIo4dM1QGKG0aPRMOIXJ+UNAcKpVqat2YhjX9s7Ki8J1rOOVOUzMazRq7J+ceyW
cEfLTFPMx8MmeZLhRcw6LycditgKnhqV9KVPyAbyxsLKtb6aNP9824HELXgl3CfVyfvTbaewDyzE
eXQSh3h/cWY9D+raowYJxLazQEag4fB8beqJSgRzBJK2i+AlupBevs4oFGMkrJUI4IdxeO+G5ps3
KQQ/TX1XrJ1nl9Zml4Td0EvFR7C+4mg1q/Yp4n1AAOIXBAFQIlg5sdRiAxzUyZvZ33cqxxlfSDqO
8unf5YU1LPcXz+8qqZpuUAoWe/vyt0/GTpXjjT0OhmGJXis9p0mWkvwzTki8+SKhn0j/AEmeRQVO
1p32FctFsA/SLS9ayFuXJ9us7XhBd/kuD3qi7xhZGxf5Ml6y+crjKcqjm65Kau1J1tKWSYNPYKEa
dXmi35K2ZvPLldi8pRUnYHjEEwczK0iwgQn31Dy7Ob8fS8NCnuzLSIH51YE8ZouYy4WQDrbEE45o
K9/60ezo1YRBB8fK7FtjyL8NsrxfNxGPUj43qkzAydkrxCPU8KP/o2/I90Mwt8QyiosnPsNjYC8D
Ib3/Sw3Ld9hZiolJCr/qiTMg5iplxQrz4SmQ1zpGMTP+yx0UkxDQIO0AoqdVpE1uRTnnAYSSTyvF
ETAzmMMTCwgjddGdvV8uWZSG+3TlOUKe+z77jkDj+VkLRXXWRnK57oHsiang+65EV+hh1FGAr9z7
ShGtFxEZ2JjFpluf4SBVrA8sR0/43oXD6YgDfcgbuR6xu7PzVk7wuVcg1FSJvd+G2kZx7r7Ntqd9
5Uy+xyk8kvS4i5zzzsOA1wuffDoxHzwYmmA+lTc1+GX+JA/5qSErKebCD5wMeC4N9SBxCIaKLkHm
kBlA7EEc/S+TW862WOYlNC5pNf7mvN2FvJNEd4LSp6MBgjcwRgFRn1b4D35QraUMmEgSt9F0Pny/
1RgMAad81o2UIhciccP7sRYTpPF4zxBtKodejep3nq+J1pkkAhG18jhY00a4ZjPJNpcw8+aLtJrV
zkUevh/4rEzCcN+VBtpY263DOXQ02cwl/87N/KdZFVeI6ZdycQClxqdSWNHQSGA6X0LILzkIq8Gn
b9JEO8IGhwzYWFu2z/W3mwikIeJRWsQzBEXex7KyhwzCJ3uhRa/94pbHzkrub599oP5iykkTvvuu
YqqP/FmvukoDq0L4DtSF47Pj4BJ17KrEEdXUcHanGiI/G7b6Jo/G6nkGn4YQ+M/6a/Qb0EI5J7RJ
EscHiEiJiLqmTn8R1WHjvpn0Cs/bAQ78Zb0Dp1dzuCDuYqAfjJ4ZcJWwfanNfRjNWDlSaNUG4L1M
XXd2Ajs9b2/TUHH6YF+bmuKDzQ95UW8PanxwEf1Hj5LIvQPWdtniljAvK6XGenAZbQs+IU86Y8DH
Ot7w75Yfw21dFP2Sk4twNNLM0y+dj8EFpeY4zOBQoFLW3Tc2muh8+jSE3/mVIQREclhAobvyFWP5
bTxH2eNq09N8GEKbDhroAKqi7CSezZb0vQpWcmUSZEz3Cp3WGA8h8EB6qDrgyzKRF+XVCuVgOR21
CMYqV4d5u/WZoqZVLQXvdhaNZiArAneSrYqHYBdw8yV7lBAoRXRZ/wqF2IGKHWVMvMX/Ga4WidiQ
IHM1nC4QZLjPP5YHe3XfQYn/KlAkVwQy0v6cxZoIh1k9RI21t32seRjB2jlkHpUJdiMsoXRTrErw
7iQvFAJKoqiyK/S7LQIP+GV2FxJ6aHcy/66fKI2+v7qOmJ1iaHPz3OZkMalAQaxQZ61Wi5EKRMLW
P2zqOMKnm4whT07aD9q0kWE1/8iqobrwY1sdm9oyeYekr7gR3VviIpWxo0Xi4rLEoU4f5aQ8WUNr
H8tFAvox4JkEAMQrRcofpinuhMeVr8mMhemR2pK5nCOenJ0nvxWK+52Xu3c2r0NSmm0CrnIuEI+F
kvF7N99DX8xrWMrfgxqdIKrbdiasIstrZzCS8iglONxmi6ikepVxZldvMjUtR+3BJg5gHcwmdVsz
fGEhbiRUdQLT5LkHqkRlm9vtdL/iPWQjf0GDg2PLBKQrZu5FjdNTWEqC0GPJzcHiHe9C3gH5Wvti
4R3Tma0AwXXoAuptw8fK/JvB/IKbXRBjqhdxQ7Jmve44aOS4LprTqmLbE8qNsMtNrV7bnJreQwAW
YK/SDzR2PuAR58lFft4CkJify67WFIlchAEQX4aVon0YAAC2U2wUjcm2hdpai77O9ir8w0nxA/qN
dnohJWbdjZ1gPVWnbpgJRKT093d9L71jr+PYhryyO96rK8nel+5YLwLF6HYlh4h9bbzc5NafUOVY
VP/OweH45iuxE06Jr6OIROauBn8CRWorSLG2rmj8mCP7O7ZSCfnVO+njoUw6wCqPZcQxhHFfZkhD
vnwTRmaX7Pa+fvvwFyBi81UkimI40drsXvp1XKaS1vi1Xh4mGCnRQ4B4CsiLTkLRPFYd8UqveeSc
UfTNA54fQk5nq8VO8Lk26rgE2Kt/Y1bR8sJgLw0i/a2QRQtDJKgOxnGT3+0ijJZ6QYEKM+JR6SWv
7/FrClfIs/YHgZU18fhxXH9ftJI9FUx7YPpliuxdxW7wuQp+z2Ldwnm/hFXW3xzzWR4XMbKrSVcg
l17j/+4h0ksrtEhnnY3sws615+T/2ZYCcFXKjTVkWURKgXg0z6+BtJZ/jfOPpLfteRTQJFIG+WEq
SEyC5H6rrmpPl5Dn8MBepECL4aeiu/1tsXA9xPMGmGiXjKdOOaavmNr1Iu7ywEbnr1qbcLjEAnLU
jwBehWbYhf6X9t3Y/F0h30VF/QH/etzOHcIIOH2xwKb4Y+s7nlnxYD5WiTN1z94JdtO3uImVpwu9
RTf9rjdy57r71WC7ehSocnhlRBU7jmTJL4KjIHODYs1Y4HbJ6lOO0sUKhPbOeaRDt+/UgCEf7WQK
Sd9aQ9VFDsnTGyY5wgLiMDePzddcpsao1gvdYMcUW7Z3aQLacL6dZeNZoRs5b5yvi2YHwXxMotOu
8Trn0+oEp/yEHYUGDVL4paLLeB6fcqFutbfm1Sv6FINeHlP5Hu+JbMH/o2dpspxh8QyLxaRgozD9
4ECIYOAo2Hi/5Ta//48c/FGWNmKPzbzPWqQkTQ0ssTqDRqzfJtoz/3sc/DNJHjd/SRZFUAp/07A6
YOJ9Ro6u3EJ9JoDM4EIIGNpKzdWGd9Ony69aBY7W8w709gtGnJ6ajzNW5kcKzK8SRj4mJWNdHFJ2
IUEpYgEMWITbKx3XkNK12YIr2YAjeud2j72ZCTXOpu7mnIq5/Rczk5Tt1qciJWWqK3oD9YJ4asFJ
UpZI8mDauYnS43Zcpn4RWVcXmhb2m0I0fjj7peSv/2NZdd6Z3ZyhcUZVrYvpbTvctDKjDnwnkX7V
wkECVByJYniqYgy477ILHfwrHE/Fw/3TFhSi362Fxn1jkTGaLQ24D3bWOqFijf9TxBs9K8FuOP8j
7hVFD6O8fAGwf1HHIONTonMjX9Qko/Jb0K0GlDv8f6S0not3BwjO6zHG4bpSKuRb/rmu1fcVs5gI
7D5OROK6V6i8K7jA65CKfh4H2Yrrt2QKyKagusZYYeAfyaUpVV/dT0OvbSi7cMGY73huvSbhIGdz
4gMHN1xLkZUhtPAM6hcEuWpl6f9S+0WNMvpRMMnFlqritSVgdl6Q0jreGCrcLSOyeSaBDMbGUt+K
oLHzORq/fIXyE1arWreR6w5YLyku1qG21Kw9hPhUKdBUM4iaUuXKrpVKOwkymJP+4pf7P2ooYBYM
KoB2w1Y5utwG6tmzqcg9lfq0QLGgjDISvZAknkBN25aaQgOF5j4lF8/XAx1UfqEotKK4Qa0vqNzY
YIJwVDml5K2lZEDQU3Gv2ZALHQIZT166xFD8r3PygWmCEBbHb5pHK1RwjXN4h8zT1xmALJ30qCLT
JDDxjM3PB/8CHrs2NQAnRAU+EGImrE7C2VTbnr482ZH8h9/XT7blLnVCHPJ7Kr5GjvHu4RUpnjT1
IvAUvdUX5WQA9mgqecBhch2Zu0lUaSPYtmrrNW+PLDB5Om1rvnwhz58EIwUHWLQ0SsCJetqA18GA
pMEH/WmTKGjr7fildb40kBauApZ9lmjoPJTdOtdrRiM3VmAVkoK7aG1XBHymbg3+H7Ubl2hOn/eG
U1+2JzB7+IrZvOn4uQEMtE1qOHNIoz1k5o6WN0imFiNI/YUXZBeUqBPK3SPWFsY7tDwO948/rQZC
aP4sU9tNcRXK//Vk2WhcJWkg2CSWH0TSgNc2t2+9CvPSk4af0YengjP9BIDcL/5jyB+ukQxDWdDj
cgPKUax1pjNwfHBVCrlN48WWfCkimjtbPpuB4U9BbXHkUAnn/3AET0vIjL9K+6oAPyKPLmQw3uth
F79ea3MGB0MOY5Dai4VQjgFGv5ocOqGr5PQVdeBHaOyeufgRRbGBCJss1MoqSQTyjKruN3+NSdAe
jx8/hIbSY5EOfT+oZiBHxIab8XMD0p7zNDwMJIulUHtkTINCQOaqv/P/N2mNUUsNvk6/cFMz6mf1
COiu+cerwsaFqEyiIg7sXJKd/eXTQkg1yuVk2OiUfKEfiUDl2nJsg/e2J/wvsZF6WVbxxcOHYXIG
5B3LvO9QlrMhrVs5W+d9ES8S3cvzVdp0hc6h/mwYWxpTyW1q8po+XjTsmI4i6TXWt2BFTKZcTlE9
Z8BJHAqsyQul2oe4wG/ZSWdvawZiRUiSJXseqoy7ohKovSVn5T0F0uMDAFl1qowFOHUoxP9VdMDb
wBeBv1HQM/vCPkL//KfoSNEdxiQQSPZTrg2xsyrkVQepHLT3n/b2RhivLWOB3qBXIP4gCMhNZfDX
friPzA2xp8JZF9eM0fxXyyUzSvtA2l8cvZptMgjbSFOpO/SLFWU5lwjNc3Vfh+N6h4bHjplgzS2m
nJCkjK+Cm2eQeQc1njGdgZa5GPMbTfJBq6TyZtRCvZP6U41h/jxbuBejdLMglKpHsm7IzZBz3Fxo
DJFtaRS6nfIoPfnp59UEYoXhvo2QbI85+NMCJBIKgsq5c5VNZqj8xtnola8o6R+2MFejyy5mmO6Y
9s3X4nuEKH/rFDIrpmYkcn3Op04pN9YOiWfqXlacPjB2TrKAb4/WYQlUr3TLg+JDptukoVDAg15b
Tez7wpfnMapeScw1MhRFmgnti/lXBmWkXlV9a10A6AyeusgXdiLpm6AVsb45aUla3Gf9ZYAJorUQ
8PvL2WZogO86cTu9FmfO9Mtgs5MnwnyEpre4r/XXECgu6tFmEsqZ03AFVVb/D47PmJZzBuaLO6vb
hKMlqSL1b7SdO5NxJWhrdQQ0A39CBbFukOZFZB2GXYM5eGIkOccmWz8LQt2FHHQJhO4uBezgM5s7
wI+cs1BrWri9pxTMGlsgOUrMAISbULvTq6FBh4yzXTadc9XfwAlkQgZyzsyA0FjJ850cQc8LGFtC
ZzYGl+hhBjUZpGuEEM/obPydmDCPH0iCCZ5gZe2X8SapMRfVRQEgrDKFnUZXMMyoBODLjtS/Ip39
hwSqQKajnoAMXFoRk3Ixp3nO5AacXoJw132hje6BxYPQcCuzHvkq3Pe2A5d6LE+/z11lsdupZC1K
76UYpsHUEO8q5H06m+ZYyGODSziQQ2lJST44pwi9XVHo03gRLMa8A4x/9JZPwhEXUvuzuBFwNpzY
Z26vZ6KSdw/y5OuHjlyE1/3OdJOVxPCBpwKJ8bYy/cQbsRUTC3OFCDiApgD11sUyXluX4nGhBgOG
dPGppDosR3yCwBHys3YCjqavrVRf6nRbB2KfTyB1iIGcqIayyYbxp0TzFXa9CnYCesx64vVuhE53
EKRKINGHHJ3HzmnCVu0JfxOh+v3ElF9ZvNee3LucO3A2RujmPy9PFs17NlMDNT90fvzC0OtXx+F9
wkQs9k9kTBuySuro9VouDNgqn0YyS5Dd1Rh5VgwZ8Ln/MpMn2aJo7Z1YUGH3OVCCRYjqX8fdSVz/
QwCMCezyq+qt7uWpkQwci3zFT0LtLWYPCnzv4keNeLIcQJsF13eFpcbX0nWEgn3Cjf9DM4BD9XaG
/d6uPMM1DMUKNjfcVrCwBpuPF9vZMvnh46+XVLb8qbLJcVbjXuIfvLRhftW3rxIwcyyvFkV/ckMr
4SkU29BTv9NRzWdgOEF5Cn42r3ymd7ZeWYVmsGpeP2nf/P0S/ESKBCtln96hO2KxvG0BJBUo9v2n
zJK6xiCW2b2nF8Asmc3/WLpsaNQNfjT/vgtzbu3kYNQTjdOBsc0a472rJgchq9L61Ff2IkdKat3g
UvICRmcZxnpTqt/f/hOIAZMcabaw36XT9goyC/5dPNUZLREiB7sViCmvZUjMb1cSWb2qB8wzM3dy
FYMU9nnh5we7DMAvscEariOK3AKztEbAbeFVznKoWel9VJ/FqEEiDjkIpdmGE7LX7PYZfWTlf/gN
cjXj4yYRlt6Sh1tCKqCwd2WjggHqz8esjVxulSAT0gNm74ZZovdL0/0UhsINAvB9GCkfN8Y9S2Iq
+Fq712XBM1jO5pBLN7/gH6n9QdCOYZtFSubDcSvoH2kF/xfAKgYIhLPiL2gJRflb17I5kw8UumDl
uhI4y13mydPIfK4+V7VeVQm9SWPJoNQ6AHIUtAvrwlDAfKAXzQhvnTY0zzviW0GTQ4h2zuzK6qKG
6IfuM0EeijJrR+SffIifw4y8xHBHgjgirQ2F59A3xPl0SPpaMuHCkhEGfprxz4OxoESTiL9B3HHI
SuuLq35eyMZk8321ZfBesSIV6IH+Q57jm/17BDUk2WUVsNPrPnZhZGVtORCZ+eRwLGnmni2uKsEB
SYI30GXJEojIpnKRNUsVeBRgG5l+YCKXsMdN3Yv4ivdpKObESUtlU4jp8IGtCiUObFbEkwXlUXlL
NzxzqlwVCoJCSfcCJ7Dn9S2yuDzeJuLEtxy5b0B8hlNjLayOCLMVxrIewdynbTgV5rAkgqgX8d7j
zuvl1AcSRWmY0DZqmuk+qKmdjRAHWP3DD3ufCwZfr5YEODwAHqJAJa9bJIdKizFF9d2Z/h8hrRax
9Vy+/JxHsb4K/tUxqwczQZwqOT3dLE2NvzL1U3l3DdVfqIkxF+I9lJBK5tyIOWkW2IQeQA4GTP/i
dOZWGuNzJyz8GUZtCSlA7H9cvze9w2pEb8MVgCwcuQgrELQdocxEe+7kgD83dAuNqYjluMzm0ZEa
ZFVdS76uACSI8ZnaEpPv1X3QLl28+w8+3ae3HpmNzKjiFzcuvkVumLfI0PRQ5prPPCTqEW/wFWZB
sRN3q5UUVKvWBqFmG+KZ36goDd3/RvROj0KtKUMhWNDE1Fe28dGt/lLSd7I2RNdiR1FyNYoSMwsY
ZoSLrf8gZUqKxkMDB84jXVrcnhmsVxpstWs5xwBEyaAcvZdIxTBy/9IszrduWCtrceas9GfJw448
mlGlVNzmnye8UIW3DwKeaANn6xBfm6ITLoUrpmUy0W7OsEJh0xxUXVJY59EtZstF6eWxPwz72QFT
hSkDre+NQNBvwhCF1jWX/WBeHLDAGK0kZa4vhhzfukuWhIuFFpO5Yv06X71FDoFT0sOwIevVWgn7
3vZ5vYk1A1BokvzGRatsEmCJo99Ipm22AxuLzegPE0b4YwXJRsEzUUhltPwVR29vyfwWR0wN36gj
YM7e9Wvxf07vpP4UYkhrTUQCRJwr/H5sIp8o5pN0+f7JzTcvfh/7aB6kVAY4DiSVA5yNiyKaKsfb
Xbp62TaOe0+X/K+NgBOct3WxcAxjLYaBSUZMgH9+wdUyLg4rp41Dy3zwtXtQZlwY2jvI4i36220q
3WlMHLbcjcdR/q1T2d1fS80C+iC/ZHlPYAbH49r9Gh9o4GngrpNGiyR8FekkwgpNxMNpzTzSBuNR
eKU+tGnfOPcJJpWYNDSJLg5n16C4dDmUX3U1Dpjf1lUF2cHyLRschvcSN3YdAa6vLgFUnUSThM5G
wJCJm7+ueZtEd09t9AhHG3VT/aTBwtYJq02Yv/FDR+wYQV/zCJVH8ijZoIsZATosZCwVtlML8lpX
GLplXoIzoz1Nv+rnW9F0PvN++1VBe7x4JcAKN/CyM473uZXdfNhoqrApt8moJVkHYOlptCMukShk
RUbY9vFyOaF/EDyAM9OIR+sJ0WsIoq+UB4bYKxZqLpsa687D/T4L3KinOq3kzSbynJ3dB8gpxWDG
ai+1fudVh0SmuOuEDJgJDzdA5GBwRmv7e2DYHjlEQH5auoKMfCAoaiTa+h4uJE0qnnYTZbaI98St
84gNhLzG117rGI8cjjrxqb+XGhJpojgFBG3+KxF2A8AK+bN1tuaSNDpviyPtmKJ+zvm+jn2RFe4G
wBcsMjKJD2PDrNQJFZYpPfQEsCG5d/KycWkwRzkkVfrdCioSjzwEMbIFNtFlnj6AjV6B8WU0erz6
nfUiQ2QyzH5Ky+DRvbs8EqVuk1yaEj9d6dIrGYvS+AgjnOw8DuJuS5pm+PnYPD0T+CtTJYMid4yE
2oZZeXHUPs8Y+ke0nOcklCAIRlitysZiyMeRBY9MIjOBqiKncaMBiTboeca/SyDhU8fiLa685vqu
mIB3Yz8v5gTFW06Nz3rmCwsxWHBV2Ojo/L0E+DdpSg1qAL5rjfC10RrhWFxQXdzoVHHNq3/F+Kh8
xFRNBzhd5wYiVf8GLRDTodtAOMDXoy4zFuN8mc25cs2zQUD/rZwG5aeYsH9VJ2QSX0CqbEgq9lns
7ZeeX40yWBWUTsl4PNHqNYp5Ju8Ubyu7UURBtuFTiD1nPOkQhbiJrW288W117g58elyAq/iGjssh
waPcFEsWHjXTiiL9CJgfNjY+DJba906GTd0PBsZNmS/1BLUWVr+gv9e4b9wJa47GbjlBXTPeVc+r
c+CBKnQs9I7zviyG2zDYdM88kvwC3exFmiuaKnPcLVkzdeopjislIkKyoS1BfgURNHJUzLs1ISZ6
4YUKHyI7K5uNjthcTDJOdOqYj20iCQhG6kiCQ4HU14B7vTycBz22Df7P01Ie63vu5BNEeVtlIIrT
bJd/LlHd8GrWLyDIbezI3jMYZlcum4mPB/5g0k47plX/2a5fdoLhrt3bn1Dh7SEQLbRNgU2Mu6He
DPAQGczb300V1ibViOwI4s9GT4n5cV68JNGS30iCzg+ZGBm7m+p4MOGrykpDdWdg7pqii9c20lli
u1cWkJxEG3EKwfRZR//BHGTROt6qSPyDUlbUwPs273ZK4G+T1S6nry4fjOuX/857923D+BNiunOy
P9UXaY4m4u+4S+6CIrLZMHxgWh52NdHdF5Pq6D86naSfZiunryp//LFu6IwmeOi8CEB7AIly9zQo
y5hB/F/YPi605bD1i1FnQ3ScVMCYhuQ8VlO1qIIVqO0wARpzlouLkC/++tvJHCPpRx3Ibf+JQ/Nn
Ghv1jEAHcSKamBIRY8HyPnwmDQ+WsR1uH+GMgdlbxxODSh4AQnLLWHo0g50wdhOUhSrG8x2FDzv8
tozQ3ieJu3d5Uws+1rWEzsPFV+RZlObA/EU7aD7oi4M/9CtsyRNOgojYtkUyPDO3sN+bjpu1RESJ
iyMSqYjAxMXG8bDOApqjjv/IYscVuLfqY419ndzuVH/73MqHH0GovoKJGdBvtTeO7hqezWObLK+R
CdiQpWSPDjPkpTsYzDVPxZ4Iz/qmiJQHeevKdMg+uEjB8uiDs8lDuRh10gS86fCmOzSmEHlDxkGx
PsN2qmXvdw5eDLWthsIRiQAJIhtD6qo1K12foooJVCiPMSXiWtnQVsrpeqGWHKUTKW3jkX8gnJVz
dci1KHG9FmZ2jhSjS2HwieGbbJV0ebChXKM5n28V5/hqoQmBXQ+4+rJHfr/4OUVZYxvt5JNsU/Cg
Ogv0X20lo0T8NL18CNElIKzAIEjZnLQ0yJyg1qdfEfkY8KVhG6VT7aOHrOOja8+WdtPMqB3+fwBO
0YDGZqkO+tY9mo9RoZRGIXbk4L9N5YjT+znTkhT1Uh0OFoYrZt9EljZlN1c4ZOFJpeU+No6GU4+3
kltmijCaE8Nm2fBFKzGl5k0V62Hbht0giZRV3sdZKogar46e343QQkRK++zHLdOfoiq62ZlF2I5+
rcK0Z6Z99NY0FA2ZEzpTOQorWvAnHPYbn+uAJfvUx/xMP1jq2MZOajlOo1UnDJUXtavTGEM6KM55
ho3+VtgEAbAwCBj36vDxOQ3GsV/D64BF7Ak5LIc9v209bqADrIB7xiMTjuZnchW+QWh7Mndp7Xv3
t9byeEY7fLpS3D65P3fTD56Zg7h+LSnzgEOSQibwIyP/G93APVnBFazFP+vavGdaEqjvIUeKsDNd
aX3CVlsQiubb5woiyli1vb1fsDg68lBHwQ8Z+4McweP2JMtRC2mIrRsuFi+KrsYqkyjavV4gFHwY
EE78gWkywDK915r/zTZ0LKxwD61MmbhD9qCEgcHtCnexiBze76xnZbvM3SmuFXbNazydLPivZISA
Y3uMOkgK/cYMyTSE0Gl1mWHaILt4dUB49f1uwn9VcRY/E5pJtDmvFghK4ZTl8juhwFWIxF1EDE6N
f8eTd7pY8JUMdKc3r2XjkcI2L8Nzkm88u0scYZn61XeNMOzNqBtUPQjH40ipZ2+PiXLKYiCd/1yA
ObmvWNjrgKm0z5Qyw9cGMXSZiHeDTlLINOdPw7vOTwJT5yxTyduLuYypAJuPvP5z5Z10t+D+Woxw
i2gL1Z1NiRAwzTT/l4WgT6IhWae3G26Pr0oUl9ma712oNiIJLu6H9VMYTIeDeThaMYVmNNZum/ny
I2dBNe5CwBvVrbmk57PTltUv2srmXVykOkB7Lsd8HujGZ6AxO02uM//35gCHgMwqbgY3X4oCp6JG
UgbDVcUQiMY64kzz9IwXdQWhDBzCP2pnJtM7dZniAxJ2sTdi1TSt3DRaZiUf7FwtYabzeC1ieBBW
Y4zBYbyahDUBBBQuWevit3WFLIbWCZEuRH4mhbcVxNwR3tNy47DrNkX1/hvs/tD4MSA15ANr8Pl1
2LhkvNxi6v6+VUECkWOZX9+vg+z5DLbe4xiEKEZDlcKSl5HkJEeN6IjngJ9KOV3EEMfVX+XL08vF
qdxSFNs4Y8O6kVnBrdWtPPs9Uy8Gp3iPWOqHzTI9p6Hs+RS/5j4uuPoIpygZr207pZTOuZntVPAL
U7zYACNpMPj8w/VN77pkObVx5J3/2bweFlVDv4cMusAPXAjV8h2QlE1XW4McaGeFfw/2E0cnXFu7
p2n46XR9Y7BL3qBP8FBG5nhN4leXLygUFEtM6KF1Yh7hu2K9QQ59AOgMVP0gspy+3LRr2rn/EpUz
BUR6EPs2U8Wvd3aUXRdeDoQxfJcVjZU058UgpLmOru/TXTs7mKmNUFZ9/dpCFt4iP4H6euTKNL/t
ACTOD85PCp7ma5PdWpOaO+HuznVXZjypKOUdg4IL1qDgp8e/z8v9KUquG6GGyOcbSKw5/WyxzTaa
vyksoDivZzcuDPAxSXaGP+3e7bCTFtd/Unu2Omimr/AXqM8nQPGPUSJOk+fJGVXYoqAjdnrPIUMK
h7FPhtSbE1UtwB7kbAe28+aZ8iIoBF0Tks42Ek1qjCdlUd8W5guhECzqHWClVdOxs2y+QpXQ3ef8
UrzDqHV6DyQvMmlxmwIJM8Gcy2iHNDo3Oc8qEFwMsYzxP+3jhq+vNAj7pwBwFgCQJ+7jvQiTrDlK
taBpQSJ789Qs8y/OW13WbrgyweOrdBjDNdQzfzNhWPLZoMaTOpnny3FCGKLOXd1U/4veJF4Bxycr
gI8pb4gXvG0JrtO0gBCbmn3lBtAiq8T4+dJxXD6lBGnKoXeOg3qC2RE3qkaWvTMGhL4PygYD3oK1
zjcewNsCgutWUVf7jkjFrWb/LKi7aQM/h93aEnNoxxNwOeG45q90ejHST52iuuwRiDnUWxGHFzzu
eX4Jwo5mMwltwVYBwk7RSVo5H1iHW9mJE/jpIR5X36NMU/R32nIWztxCnpr1xx5rvI11rKVl782I
Afderw5ZJ/sOVom1TUtCa/fHjvyqajwl3bbD0ckpcvLDJNQr/hQjcktY9TzWAWW+MKIg8XmS3dhl
jR4QZId5q64MCV02ww0yuGjAgsNfB9pYTdC9t6jbg8ipGcpEdRJR9PxsjpjVBXRTdovnm6Bx6FLy
SO8Ap5t6q6wfBjBdKHFndIQQZwIFOECOycy+yo6X8scjzLbgSRG9z9/P5RAyMlW6hnQNfUhwiFcF
UAwdo/12oaEwlpIG/dxBEWgrYYfiPO/q7wvEhpPku4fqIpqu6odNiCSYTjAUjH6C+qQbXkhxy9tb
nZYBiAwgkM7Xjv2b7sQ4PTHiEpTjqzj9/EU+7ycM7TCEFGB+vHlWCx22B0mMKHLfCF68gKzH9HTv
x3vnULXq72O6wGeqDppS9ysBTcM1WUqCCWuNKPQwPWlMJd9W+3KxA/Wd0cc3spGqeTL1gT0BPHXf
9B07siRptMyTCQqbMenhsUCDTH8r2w67gYg+MAkNr50DMUIOK4otuU1v3slCuy+y3RgizsMPXRPh
knRsfICHwh7TMqc0gn/qDM/GtEgyPEjyWF8hEDqx4nLI3g0WaNBN/rKdUJUt4GdAt6hVlukg/K9Y
D6fiDg2zY3LDmuDVKMIjTwtLyqTImXKTKtVQXL66huZJuf0xvF+8Ep1zj+xnNIBjuVqK5YrA+ar5
A5cGSQXFJ8UDXtLLOJJ2WwUT6cSqh6C39Lds5pBMfo9DHv8dzPOK1XGpCGjGOgupn5lfkHIsnaYg
xj0eXt+c5H1JV0R+lnB7bLnmt/vPkYrK0JNGIcReoFVnnecKsUhussB8ry7V53YGuSSl6SLQHLM3
cKSiXTuhO4tVBXVrXpznW20RjC0i9duBD0soH8gJRVHfDtruT0RAxT029LqaxGGzgMvi6DC8W1qd
FPeJGg1E5tx8aO3I2Zyfh+l8JAWrst+Ijit9i+0GwMAo4DYfgQknf7Ggnt/NmRvLXF1fEPGepay8
WXbelTb06Df5J3toLEbaRON5N54VFKqQ7Wb1tF4Ernipa76QYH7ydipI6vtRMC+icFExpQcRIxvd
g0u4I6P8Io2QgJuDuugbCdo5Ti3DcttYcfAZH9YNYkNo7TGG0MsLigGVRzBlEAX8FK4OnjQJhUYh
UxIHLIS8dkrZbFfG8Ev5u61jQx6RKGRw9nSCXPchK221edAZ+ke9B4UG8It4KN8c7TbX61MLCYpb
ZxhsQ6Y0/i2xdaHJ6SFQBr0EhSQdatdTZ/mJy9GDUHXLgnnNJHWkVv8rdxcJrzhc10zUYKKFZYG3
A/xz1xMCT7VRSowkxkkufjZzISYJPhDaiAYNVK9NpEr1dh8D27qgkEEqhI92ywwLVuZesjsI31h1
1yeFiDB1FaFbsjBcfaw8ofHa66Cl7srvcQPyxP4IdZJz7aAIo15XVbF4sYzqggDDSJqKnbJoWMbm
waqHX/0j5UDAMjxRCjxYhUqFo9y7ScGxA8Q/dyUl9YJlPNFu4IYMr2+7P+FOfkW/04qH7DYDP52y
1cHtpWzxTPAzxAkQnKLSsqfNFbUHbWtrb5QOXLiQNZgvTTgplFjnSL84c2FmoL9pP9/aaMv8sS+J
wRzoV9V0gjbRaqTbnEl+KqTdEl/cvo5auzt+TkXXU96yjPtDTlatGdrv2Zrfuk4OADdwlpdgQ/5l
wKfz2J6x/fC0zMlXiYLk1UDTI6nA2+dyP50yCuuvspED0cy+uMvM1OlLyU2Uk1+MIprazwKK0DdG
LBeBo0eDTbCkM39F8S3d2w9Itt3ubeCMHe8k0QBpYxCqiYKME6VE405M1prHZfOSIxBQDlPY2yjO
+yzxE0OUDO86oT2C6DNF4etKmFiSR6ELwPvsENUZS0XRWfGds5QFiQRnagJLdSm0xPclhSkelR3F
qdTjgKpfxtgLTbUfJADbzWtKpm7GB4PTB3+Vtxev/P31I5Q4KMp3FH0KtoIVFw0mXCzWEIX5x5sT
lDQfFZurrJNjRh91nsOuT/HykjAAM+unhWLxqi76U78eaDHJVBbwX6mDxvLR+rlON+AdsPbIfToY
DcXp7DQEZUrZOtKF6DBmKRweg3cXRUWjydBkjdwtrUQvov+txHc349NHQXRaqZcH/YmCuPyedJsx
30S2P4UGRRTkQ2xWFZyn699jCOER5aCoZCsAob38l9eRRzox17vNeBED9nNSLcQKT+CbWmyA1689
RBm9Pk5ygfdBxgSxspqoF4orZZsuWd0IYoI0aWC5D53QwK+XetVEcsOt2+G1brS33VlAHf+YCOml
ORAsbYjWUhCzfqsLY4MH1ehOt/ciyNDays/icwnN1PkmuLylyP1IkQO3SI8CjQ5B1Pm8RaOMtr/B
liMeomstk6zTH8kDP1e7EabjhaM3HrVu8wiblQJYLntnFi90CWRHSQBqycVLCwpV0a//v24lbZ5v
05q++VZ8hKNay9fhuXQBr3ZN2OvM9wG/Y6acxzo+rBquywH6omY/vrfjBSCEVOfaU1FW47Cyo4S4
NRjLsb8ATOJ+/N6tZTCw0A74uCuP0CcY8GdkUobEM3SnFvriLIL5ZJ157WjXDE94v0hdKSVLh66Q
eB5eM43NQ6x2y+bcIGeuQurTtcbWGggvz1IDxW81lRVyu7xkPjaA+nEEkRgete+YOPB+DXkqLx97
Hmq7u7Rqs9OXhSId6iN0f5MRkXZNJhQdx7lTeObEOyYFdpLj8sYqYawSI5N0uFnSLAgMV5rZwV43
PpNil0ycZGt8ipB+29j/aqlXGceHRGJ53EflBlWddEgybFRmdvQeN50R33bpXm3QtqUuM9bZ1ICs
YBwp31OOJKeb6vS6yWrMrsn+5XZDS/IqiSa9+h/hxLTCn9KdFGM3BLjSqh1oHLJtNjgt58zUHv3Y
gse9B3f50KAPZt0V80qaLTja0mrfCHnC9Ynid/b7CtENw+5nFzUZfjnIl/vsYqUxTEWmaB1aD7TR
knZvgyhVbbtqN4GDXUzrB125Im+iV7hJVrZN7mbKmpgT+qjFnGSA3AALtWC56rLsUoRZcEular5p
g2AkZwJqBlHnllohuKuk0CUP0oXJuaKUc69BqRK5SC1RUyDIo76EOQAFANgYJ+dDyEb/8RbD7ha2
0k8SOpMEQxXD24ouHjCQUXnMmW0fjrElAPHKtPb6zZGhUkXAzk7NMecFCGtn0qA1BLg7DeoiuZ4W
Ls9++tlHuae325msEAFxKzEIRJh+8EZUcYt+nH3GNnDTTaGNQBO0iwoKonDf5fM7k8YAo1aC8/x1
IRCD3N11IBRwCZTRmqeLhglFVBVWFOsMh3IFLwOM26b3qqUY0Rlg43IwyXP3tL8X7WZwj6855okY
lzutScbtS3PgeHJjuCpqqxPnwoDoyyao5vRtZdbC4UTtpBbne7CAqL1p6RqcACxwBvlzs2CyOwNN
ENxmgQZJ4i0EUtt8GSER6UGX53lwF3iwVkLgfbHzCXXPLeu8O8LC8je+HKvs8S+Ro9/LifP5g4zL
MzM/U1SgWOI7uP0jwwYSAN7eb6FJ3Pz1AXlHXnUw0mbYwVIHknSc6f0m3GR3gBw9mlyGk3JY3j7d
BYphRKw+bNzMPZGCmzR98mDyMWmw1LdhG6zMDGtSNVatOMyYJFe4cgwCNEXi5D7gI8TwCnP+D4DU
QYL0xWKUhAsIDr9DmreZInahPhM8L809qR5tvCfsmQBGUdtBvVOfAYI1OtW6lY0tLpXb63h4FfcB
Six0mhXvBxCiwZh3Qudh5di36NB28KK32jAuHhixZSS5c4fWlgIPHTatNatqp4brKZk/XhJrfvv3
L0Jv8ecgE38DUHqWdu24zB8n+Qh6Osm+1PoY8LGtKU+uIuHSIvPf0ZaJizXr6vk6pTQ8JSRa/fB3
GpUvCW6a6+8gNUtWnldOHEDwKIfgAiUuKBvhcL5oi3NjUPI3lmxn11WiFTNgDJuQDogwEhRM0bpf
UIvAVaF6DY81VcyA1iyV6HNmMcfJlsaXQRM0aFbGPDQ3DiyqJYzxu0Ey0Rs/Nj9nFft6EBkFe56w
/2rk3dFo45Ts3xABrpI+tCbcu/XuRFDd83RDKciub7JkuGwUqWFvvC/7hgoiOct9Muxsu8NmGWh+
PSKohu63tmIaYo5R4niaz4YWBlYoSQvdt5OuMgiwLhyQO72tFAL1WSe7ZkJZZzMVnixZ6CFx4fYr
PvxZPxZfSwZORToQbHU17Q1+clzyR0a+saxbsrMMREs0FQ0vA5JfkVNtfI7r1nOiev90EcU64s3G
VAfY5RwgC4S/Twzj5WJdJatL+LYpnT27nUql9R1M4h0Hp7FPOLxrJydsi/zgu5R0b/ftCtXug34X
unNMxsaPy3bAgkI/2Gs/pkTbXFPb+RSdpAYSBuBN0sekMGUDoiDYuhmiTSjh2Bmha/4slfXVmqkG
bPW7imbdccsFZyWaUeXqKuBIpPbN7YjVhj6iAwmPKkR1ip3+NxtRE46P+aBQXlpjnf64eVAd0W8q
qGcOjvksnJnoy70VDm8YnJNaPootpmTO5faMvfF38IGXPW8204HNVtYvaxW4DAdXSzFr4E7h4TQ4
0Xmm1N/8hNt1SujGWrEGZTTefLzxwpVkeHGVA6u9q7QmEqIbcNG2Lah5tXo73Aqfj+LCkCvJY9b0
nmNGvTEcbZkPfIl4h89uHz38XABRA3sTTQcpFjc7vm+wlokenP+orv4vMj6o9NqT04NN5LnkpZve
KrzC/W3clDmbVI80Q34yqEH9zNAIGoD9eaf4fC5sCLQECQw6SwRZSHbA3Z1Dy9Fhi2jcT5NsHdnp
uhR5+XJDhq1l1a6SjizN8hLutT7s9aLYIQYBzoMyXy1ElmuD5uSUyC+o4JZB/YqOz+ByQc/22BrR
vETR9RJCjWcDmx7+T57g1ipYsIqW8ZYrqbRUyJwK9A9ZpImoPaS1CkzcARGBXosP9anvrOiXnSqA
gb2uWl0/0UnwZlwEjIzqR0Plw4Fqyk1KewA6xqlaybHFgtWPcaTPLm0gMrcMy/ItuwkzB7+gSKL4
sfv1XCUgZ8lBfbvvSunQ2L6iSUTeyIoOPYLMP6s7mWpZSSlAW/6FcidI4fOj4qoGpbrYwaHIo3y0
a7Xp73Wbxmyt0h+s3KOWDbqreIWuAv/ODrZS3c/hitJfpXpxgQ6wVSMymjYj0yd+OPzhxnb5bL+n
YMkTqf2JbjT+daFxRXAbnf7RQW3bPOsk0t6XfIAszaQCryghCC833f6Ez+s/rMXN/iWJSLGQmYJi
K9O05CeBDwLJKWiyblS0Is8cacljut2GXPikN12drE0ar14MXQOrMFddGamz5TnI1C6RKBOhRKqM
7LXLHOxU7+fu/PwSBU9cZoUSBsU4cGfRWtJ1N5yfdkue/JScwf6LYHFI861vV+gQaJc2vNQ5DvYv
ycvg1WxQ0+6/QuFYjTw98z9Kviwy7GTrSAvElv0mUH7SLnTamxGtmcLiHxZoPHQSlt0nejQ98XfL
jjAvwvyhPcRBNObfHvS2KAQPJ+r2nOi+sYm20xQT/1MuwkMX0QfywYOI6AFg7tE6oZlMWVuP3Dgs
KU/1QvNkMd2fPJxvnPQ0x0XDWC7ujZDzQRVa2pGb4Tpyr0gZBJTmDOx/cG6CipmqjZpqaGqj1MDu
S326sCA+IbmjXetJfNOvm+A0O3zUEHgPVe0H/3gwJQdI515L1bQJGogGxUAfBLd63nM/20U32lJA
XtezIHgYUd8rgMl2Asb9vA6xkPpVVPDxYJZMvgZuXoZ1pKPAyIBk1mfOA1H8+jd+IVVsaoK2Txgp
Y/AIFegoHV5IU+QPvdUWkm3jnLo6C/tV0kW/++cG5FsjQiWs6x6OBWCRkPqN09PK1aOdDfBl/Hk0
EjKl9Kzudpwx88Xx8bwtQ53ouUUyIks0SzpBOpL3UuJ6VOPtt+Q9WsA4HEj/hHahc0vo/RIFJtdl
9rS1wJiCwDWeTX+rbZZDGBLkggg8DEdWciZ5Z+e8sPHu9Ep/OgxdKql2ImHjyXoR8zCo3cWwzCjQ
GujiLDX225WWYEzKNDO63u5jhIkOQd8iYqE9899UM1ok8+Fe5Eo6+hqel+rhfRtVMFLkiMy/npSg
KYE0fgW9+IMuoM/eEuv8EC8FGGw1UTVyLfYHvhbLlxlgvrP+6/DOicpIGta2139RpVC92SC3HIAz
PCZ7Hx7lkLnIkTwr5+naSuGoPmPsBmLtPXYHEfPEZUbdq6diHXmGDzcJMZA/1boMh6zrtHI96RKg
f/dB4reNAov/rehiH8cx+CmRjufK9lCeHhn4DUA7j2FmiCm3/bPQfqvqsoPC9fqJXk6WHQru8zvS
uIxKDNoEOIS7ugNjAPPy2elD8DCxwhk4pmrXc+nQfAuNx9kWMBeaerisUcFhwgPzMqFWQ0KYD9vi
cme7NPfs36AgFUVUvCCtf7A41hThrStWOKLLWszldPMS9xJGmthkYwwtG1yVotE8V4uvYyA0uxTQ
OWq8sUGtF7sF5SC9TTAH4QUm9XxhDucPxPxebZj4c7tRhrDAQP/beCXxEhSqDTaSy9ImdsOVgWGz
zgbLGbuQ0H6ajE1hDi3/+Y7qoQA3Mp27OLb1TCWQ8W0C7WdtA3yia+s/yPZroUxQMKWKCFbfPVmI
SwBbuUXQvAq4da00LezF08b6JNTrbpvt6vZieZPW/Ss9saWiJVXkIOaoEV71fHfwuSg3V5BEIhYG
63kak2Ot6k63bUH0znFLPpPyRF9FbJCxSYYA+92ZVBeXzT6wB4jqrPXV5+GJ2KZDFwxHdKV5GQlE
e0Apsx+PwlDgMjsXFUE/UzfLvUrKKJ6SGh8Q/Q7gtlZMsiQQhhuzWIIep1GFA8QYl41Un6QDi1YL
nFwIffegPLgVqOITulE8gzyhcsqqyiIPHoW2kMeFJ09UhJFVCKA9iNLWk588dGFyRMTs+FZMZAxZ
qm476pP+sxSwKd46Qt84/v/4XIQBpYkMZ/8Y1QpjUFu9TYA2nH2kkVcZZC8ah6vGitOjFVOU/0lR
wPYpA7CebxN/30ZdTrtrNOehFBPs5PXtxD0w4hiqU4OmDlOcHevTQHAPtBHUAZVvUVlk4quUbzYH
McN47zNyJE3IQi1f2g4Vu4LxVAHEB4khdxZwlcBe7rNiGL+r8rRXKFS7xGvKAZtPc7KSKewgL6JX
yey3vs5MZ2Ii4JCFN+h9Wt1m0A9Z+6uixNG6zo44Alma6qnCEsHGoi5qjjaMl9NmavLaOAkSqnUF
kmgtKGatXg9eJ91ZfbuCQLnGVpBHMnsi3R5IFq0b/mHanZY1jLC/kSauuZ9X0TTL6DdWJRP4Faxz
wBo0rQYTjhLfelOFFEHt7wstgpdRehCKTs/PYrAe1WDnu7JpbDrSkbPpQvwPVcXA/wZz31yaxOxc
h1PQRVsc5gLKXlBOSWSq7O6/bSNTPRqSn/xggGZvQOUpe1jUhrscsON9fiuQykkMQD1C0HBjwGgn
u4zkxTqBOeOWU89xYlsR5ti3qGy5Pm236s8VjXQ119/LT7kYuYcbPVz+OkWLzlYSllsVQHQPjedj
RQ2N2Ww+DXZKwoOK7aSlrfWbIbRbJq1/wq6KQaBKHBEILwWXYGWZOJ+cAPUMpC/TILOYkSUohu9o
EcDeBuJxyUuB86kchBpvRisW2hGVqNItMm5N/2OrrSh+8B1NcKP+f7sQ0nL0LgOVfGmInkESyyG3
YWEKe6FojeIvMYfFw9Y1Z3vKIJUgxrbiDq/96Q+dcbNoYRyNFqjRoPuznltvodyiI5BjxgLZpWnA
dVEGv40SGiXSDqrGBv037ZqVxZnSgGW8oftKWCIRTUM5T8gO38BIfEHzACbGuku5oXrNSFVTaRsY
tgZR6PE1TBs/Fb/PwxhYfqia9/VKr60fQs1Ie4EPY/I18K9g6Ahdj9wSdS60Tg4XGJt5gAm2cdLL
DhQQhzbsay28hhiWevvzAmQ+7JG+yrbCgTZMX+JTS2cTQmFjdNkYqGkYsffg4DoXNiZnJ4/KovPG
uaAKKhH4DNeTlWa2abO6J/vi8OxJKFE9ZSHW6vl3hoVyVkzY0rLKNs1qcvOnHKENU0mcZTlhGH0h
aEOPurY5s9Mk3j1JL44iDBx+IXHxqsVL9MgbPAGxELNO6gpK9PKlgMhKh01xT2h+i1Bn2aGSzQ4B
DBxhWdiMcwsjfmFM6bC5w5U3yckTaC/3enZvamqNUIB+ueuGIgVIfasAPs9RZ/I/qsW2iUwRElan
Vq1q5LBmm21v959OQeJZFKop3M83RGmyEZMjAU8srU3T1Scorl016rP//Bmfo5QVzxkJelpFZDRN
6bD1v/AsZ0sfLauCSWSA5gawf09Z1CJeclhTtVyGmdClcpz0ioV0IPGDLU9rJUMW1EVofXlo5Qlh
C3rQmgsdSDAvUA/inVI7BXC8Wdhp11a+qj9R/0gw4I7B3fETPu3ouU80kQ2fkTk6e1rhWET/RVXK
sFNlfeVqMeFMvG7HlOfgqNpPBUOyp+6RxuvD7vUIxOEOULb3owHOUp9G4EjsiHok+AVXrCVp0bep
xw5NsdWFDDcSqjeKDocq2DLiwFqSe74YVeBJ9WlaYjzUVu8BWP6b9ri73f3iETjmc6iKppzQQ0IX
TdeXD/DzKQPBj9fA+1T5tz17vw4P5baH41j7o+aYrk59yoZobgntY4KPe5ZVvkoRMguVbU7GOwTQ
P/SaVRFUwJ6gHR/U63GrTFh3PxMahfGrX/YQ+q0j+UQRekAeirDcMX5yE89P+lRpKoOdNJtPu0AN
srP6LrCTyTb9tQkgCVQF80eSC7TfCUYiBvqDrFg5m1Qr+/3UFp19dPL89O7RhOmbKs412AlIJe3W
qsOWpSwlXNVE7zsH9tbExU2f3SdZ6mQKACPxHjTJDWyPw//4fRk74lOYHYJiD77kRFutpW6LzWSB
FiNptC1ELyfdPzFibd/3a04+BE2BmhOyxN5JRa+E2iaPMv8RGep3DhLDpfkJr8jki1rm448gwatt
8WIJIXhtEUnT3eYnZpQIUZNDksHK1i+rWO3HNjpHCn0dbYIXsXyx/8JUjWHTG8lWlFuVegqelrEr
65QXQEaKQ9Z3TMzDBBGDhhBnV+IgDSGnWOc0NCZcgOdKMUzyDhzHjJ47QUm9y5NCC2W+IpEJ9x4Z
vxK8KhVUwcdgEXWpGW93QiDC/kEgNv8Cu78JryE+0B8DFPZVbi2knYLeEpt2zyf+4/DBmfAKKBF9
ebX3XQ+okXl+lQD3qBU2xzzudN0cX/+gXQVyYLAiY+1Rjv8RVmTZJFnXVXyt2Ho0Gky3DqLXCYEl
VPpqi7D5VvlFEL1YqPcfycx+85Kp1Jbb2ay28TE1ykIp2rsPJZw5SoMT6vfgjAGCialRLEMRT04o
rnC2MGM1BmD/lch1XobOCPdry4ocaV7Dh/XbT9Zujty33/s/gBFDCyr8AyEtKCXZ1tMJuJCaFeC2
8f8imBn8ZL3toZ17haQEf/Xd7pPlsVBPbqg4nEPOT5KGbRJupEliumNBneqlawOT5/a2KgEw8H7F
JysmH5z/7Dmu0KOfMqVIBD6jTuhhxqeaBfxNW+p2pWTfmSI6h4OGdfVSclJpqEcrZIfXvCfalvLx
51Bh2mKQ580hXdf45Ac6Nwg7U9M/3qvcGqrRsXqEVmMm7tAX8p2dHj61TEvvA3B++f8G6+xzNNEU
BZdcF8zxu7IZ1NTNdxQ/31Awswf98uMNxioVJih5WsRAkoiUIgfK4s4KSMCps57PyGjmhEyPyc4B
y5eiPFvSXe1W7bGidIfI+oHf66xON9oXbWY6P4BR7ZJLMZhYVJBlVOqniEqRs6fLXn2KTunhTapg
tQ8or+3uUKaTGFnSMLD1EddZyK/12UQm06UMSN7EQ4MBQOhzvXcYKKHKe000DvYMecM+fp7bh+cK
A4m565jqrClY7rbJSD2jyWOdO+x+4DZKhDXeG+tbC7zVWW4p9SscXwY25xyJX5B0sw/BHu0VgtRk
QxsgCLWBlxb8RMtoiK2qU1fQ/XB+Zj2PY5pMJPSWQ52fkeNg7Ybn8BsRtUEF48LfFRXAv8vWsZT3
6FRaX5LNHABRwhO8xeRMRQ3ntFGOjcj3z3DVKsFCEG/35K7wXYgzC5dc8+WG2s5gugdIb+6Bz++m
S5Isv2nj2m/BtVzfaTXHhrSbaGOnO0HAjAYneecRYW61uXpxRBqowid0kKirPiWprorYRoGc8n/W
NwJIWsE/wERnjsN4IeQnR6DFmsT4NCgrXbEoLUg8gGYO5ExIg+tg3jKXSPtFG8ehXKGzIKD5EE8l
R29EMsRdEIwsX2rMvIhV3Gq1FgIlZQEbzf3KwnWDv/X1ubk408fuS8CvCNlStzeoTDSjxDiQG20S
EBQ4RhF3shZey7YJgH616LaDLlRuHrYQH1fGQzZrvCDUR6jD4peh95L3ofj6/fpQhALwD2kNFZXu
NH5IfP424TrJ3UHzX3JdAeDu76wC7tZX2jyUGGfPO7/NFrrnPeUFMEHBdp530IUcyBg1+cDearh4
s2aOgoBXiI6LmdU8onDHaaEStLF9bZ667SJTSSnp7aV/f0OxmpRYAPd4b+OhwjlV5owsTYHPoBE1
9HzXJudEyeAis0sBjL7DD9u1h0IHBLEbbMcJjrTMc9lENFMWFB7pSXhNQ5WJL8NkKU4MrAvz38sP
4AT1S2orDGGP8o/Lyf5q0Mr+bIXXLMx+DPooH/klH1AQHcv/sOcF0vyjspHclUIdF+Yd7w1I6R4u
Ovep7VExGkdAUrN1pdzzEwTiFue5yAdQJBx+CthHazzpbIhvX4XNF0KjzNRkOMIWNAzSsaCBtGE7
aSMW10Ehb9hNakx+YVWXRRQVUjPK8X43/XbBgifAq37yJwD1VNL0xHdHXsXS7LOM7+xfTlP+cnyx
j7uA3+JjAXg3oaqbk/udRxzcIHEOyU9b/TsKu9bVK0yZJe0yKdjXCqO//h9Q6YHpTFK8PkNN//3c
21y+unPxEQZFMnAp5GLz6ZDyTsadvZ0BF3wy+uv3/9kIwc3ZwCFk2B9ipw+Z8eZnauTjqLbl9N/L
YH9Vuqej4ZE0MfRES8ch1iKfvCV0kLMrinZpbt3cU3zWobRvo5Z8db+9apUPn7DqINZB33948FHb
+dxdsyIS8FGQUZlyl9LKrRht9KhEst9izqBkgY+xI8A3XAvppQ26SBvwL1l/TJwk8fqVw8hQ9EPu
qSvEN+4OXquMptF4VqquhuaJ+yp1cyKYDJ1gbePEYvMEItRH85zSkK1Q97RUtbVbGwE8njJv2TcZ
ae5+ZkSLoCrCVLHYIRtbeHuiVHWidJRNbTDeUBpo1Se/1mPm80K4KdilIDVbdOwx1emhyC5q8X2p
RG35drIFv88pYz3tyWwVzdy16chNXDpdvg3UVDxtokTDryaV2bGOXoH8iljuUcC6sKxqeznXUSsb
n4o4gIXit7rTkSR+OGc7G+dL0jhi6j6lvLFXU6QyYpuN2QdZMbKd/BTEgzXEyuZVSGRndWMtxVsy
1jJLKl6F11HrEgCB12TxkdTqVLOQfNUpcyAeYtYa+xSec1ziJVsGC6l30g5H6iYGeROYjkg3dhHq
mG20uwEt7/8GmNGFqnwHkC22/XKJqxLB6f3Lun/5/RUSHrDR3sRuOMz1y5C707iXlnDIVw/e5/8j
Vxk4xONa295UxvbbZB2ZkN7ktinKO/fIswa7N9V+P5m5W8BiOboYVoYuWDHzVc54MYXDx+QFzSuS
HIwDdDmNp45QO/ebT7uUuIPJcmN5DJIQduyZWw/SSdVf1mm+Hqpx+vTWeJrCPKI86gIHmYHCLj+k
cZIvo3QsdGh8DG1xHCbp8YYak9xWtL/40Ka+2SPPNLgY/T4EWZncEKlCDX8hmbKL7H82jaMmlfhN
HQr/0jj1YMNBp74BfLu/VsTmTf2G6ap4bE8rxdk2Sj0NQOlLDpzh9XbsAwtTlu6FIzsJrVqxlWam
VQdMzPoLug47pVtFF1qSNfQae69VjSnQn7O3VT1TIAe+R+ZcNG+1LartbO1zKbMZaq0EAY16RCOq
Syly2CZ2InkagajTryAFJ8PQ2H0+8b5vrGlQ5T2Ujdwol/IM/G/u3O20WMqqlJoQT/BICtSV3hpx
zSckeuHa0ivJ3tT4oUUBwRSM8TbNMVfeL17A3SM1slfs17ny2QJLCxQVkDtsZWe6qMMM8ARHJWC0
unpff7UtI0IB9lKbE2MJ6Z7PgoaZ0J9VKrOQY5I9AJWUi6lYWDyV5WoLEC396qPc8fk3m0LsthPF
17ckNf6LghLYF/6qRGiWXgVU9G9V83m5nC47PnsZWVIoAYG7CIFq6V6EXPY/gUUgoBFICPVsf603
uEqNcBx604yesFVQvyAoUbvhwZt4q69T6LVyrM8SefgNxdneXrQG/ktJGqdpx2zPHcgsxt+dB/BX
2nYutDD8SRdb3Ji4hV7g/N+SnxvzKz7jKOr6Gve9Pwt53zZvGX46HXkXqx5SwukrbtcwfJND9rsZ
CqMD8CWtnlP+nQYY0CwtxFEeX5x3jqfhJsqvU6mZklad9mEKsdVDceDvC0trt9kBb3PMerIN1DyB
yHSNju1u8BeaV+eRalMgNXd+zqeUggb4t080FV0EcQk/5K79khZr0bJWh+sOkXNfNDk/blDP6QL2
cDFU3t9FyhxUEbyTs0HMJEkezByq+xgN8GFSgHAlvp9WLEk72kG2+Z9rDT0J+LptOlOqZbR1mr9R
YSwE7zMyuBeJkh5FqLtSuqyTKdq9zn5W6ad9pQpN8N6NM0sSkKdwjydqKYpc1Yib32SLWDU4/vIP
nLlf3ZCffetN+qVY94OxmuBPDk+M8dmpv7VOPzAaOvS4mCRmtLF/k70GOeK+HhVF3P3FPs1JbzAW
qpC0iZZpdaPf0HEy3Z+N5xJr4DzvsTRymUohAAvZMPEBDveqn7Hf0nfLLQ7HDTokurxtkQryfbA2
sdCyNrM4txncWLyr7PxCdtXjypAJv/KGbJUPoQehcY8b8zR1jhx8nAwXoWt5BRWk3Z8Dx+N9Rkhm
vMXvqcvzLZqBC5yqeJK7ZlQKrb0b/VqSjn1q0+Lp2jSGhnAsSijjezzEhhHOkw8ohsreV+tTSv8I
qAPsD8uYcCP+7lWlSxTKPyETleIPeti2pkmLQhNVa6Kz9yl2MZU6ysEPo36uUxGGjCQ4tJKJtwpQ
bBA19Jyu4lBGtLfG9wo6Jy1bCJx5YaIbveBlVg9yfGHMbMvKELmm/m5fPrF14dH6HhnfoarBhgwP
Uk+0dVj/LyzVIq911P4pzEbScCTsvnAmWFn+sXKBtEzMfQzjWzJMyUfvq8FrHHnij7MPtnQj5oOv
a1hKWD8ENSLk4kxgPUQusHJ9t2sBDwrIFRRSzQ/m32aGH5DcI2qkZs/oBS+EcN2sjooWy9OuTTGA
Gsysr8oke37a8Xeri0GvLj4YijXyjvjtbRJOw/QuhX4jtBTg+Zph0osX7/U4hslhlcebxBHoEG2E
UkPQrHNB+ne7Bfn7Ug0UsKiVlmoovY8qknv37iXs5sNceBcZaJNrTz0z5V+qFkA5MukfNVtyvHEX
9l7v0Jl8eFesR5Gj25oEdI3enFk2/Jg6/09WjpF0UtvT/9gr+qbh6Ih42HkDngp90o97aNYH2cFb
3p7TXb1uoVkq5jKs77DKDi2WFK1S0ll1WKHgt2JY/f3U4+L0DOthGK31c7mwGla3o2r+HYRooCt3
Uwh5eSkSXEmWONvKNH9h9viqScW6W8SYOq2Qii1JXgqslDI2eTD6k/1Qp5jq4rtu833Iqk/3d71P
WbYtv7UkLuyww5+Us8bfO1q4jOAgi/hugQvc+V8cHgIIiqXWir7nzy9K9LmI8vNEgb0NTLiesjkB
Np0oE1cVrdsokB69zXiY8jxJCeG7fnCGasDt/on9TtRB+n5Oqe9GmBc2d2bjBdMV5XInCQBpy4ng
7pWFPLwxbifgSvD35ughSR+T5BuBHK9Ibcck/y5rw2V6ZfSJeNuun5pQ4/2xXB62vxjvdN5NVizq
pYIYGNrRcedxKptenQnuOg93HruTjF70Ltw/StlV8W/19sM5TvdjWoSV/khMY2mEPjWAYZbwHzLq
JGxdBy7Jtj0+q9XxRjHFlVjTMFmSHiSQ+MMnxZdN/uE76ghLAFlIcussE2tTo3SF254d1gNIP7wo
PiGarkW8MciXPRP2t39QsZpdx7W5a79ygmqIdkey726/6vOlEcCHiT8FB1Qleg9S5+kyvSSez5ab
ZyirSWoGqqKUddD3vMDvFP3CTLoy5PQJuDi7jZm22vhTuw+lTGsE14GvheaudKqc4tmLIapp7bJw
F4zs5oGwUt0MpPpjtfB1cQNv0ucV2F2s2v2+89bJcDUk3GGU9674XxS/plHjED0rRrR1zVV5hdEy
Hj2gAvhxvA7TIxPPNInuTwyqisppsCQGeLr5JzUdEiVRE6VSuUo1/5NE+k2uo4of/3NealU7MSqR
qNPYmpSdW4cJI5Nll7gSN8IlcY88yHZeIME3l+9PLso07u/vwHqiih2UreD2y3QhT5RnbCvf2J+y
Gr2DwW/LcBtDkr89MBRkyHcm4G2lbpQrWt2fVyYSbiLFQAzph3qk8UzkHwx+ya/No7Bh63+zE/zt
nLfUz27EhgXW/ADP7cUk6OD4+iPV1crZtOozClUXOeDp9s+Ar42h2Hh+MngyrsX9X4L9WNnv562U
1Vp873wh/mkv7G5ulVeUiFXTyHvMVuEpieglt1RkN6hDq1v/ASUGTvTU5VLnJoLPFSFq7NS3qJ/r
4tflnvAAjkJENmXgbdvoHT0pqULsrYMljMldO8l5oN4DzgqA3wr/2Utf8Q4rPf960tNG0wo1nLJS
41vXhsGWlg+JYVS31H/eZv8gpVKzvbVyJYoEXa0f7ZsTVCouHEmQTNHe2gFL7gnzA2hANN+uuX/t
LgAmiFp7OCpOKtLst+N3XaC08Vds7/nqHC7ZyAAb5jaPNSDaPTHpnHJa9zQZKPYrrC/7rgdJI1ag
SlPj9lpr7xOeWAL6q/owiDsTT7owgoiNQ3aZd5Jqu3IT+are6LZD+jOv2pGr6apgzqPk9nhTm8SU
npusXLqievJh8ThEEPeWCDutzQBAIl+NquoJKnR+cxzBqTKwAK4UjNSJhxK2ZEyXSH230uUxeMqn
zi2GpCFT23G7uz5upbRXkwG07ID49zuFobMmu35L+pj/HDefjY+RM2Ifm7W0oVZjTXQpFSgt9w2i
5gXQ8Lj4g6bXQuXGg6TfP3meeldN41TC904Y9QADGVZ6zRBfuFBAeOekHhl3LCpxaxwxpaJH01GL
45zUXBoAXlOwWVGpMHbQ1vgGUEyOVUSGUo0nE/wZixBBUj2DKW+iz4PQyNgHEl8AKoy8iiMjwLTJ
6rQeRdLJSTg/euTCFMb3O125u85ybeWIkRP55cxw935/W0r2HFQ0P7HZbxTMV14W3s/qt8kcfo5J
jlD9j6j7GBtJExG1CRXlFIr6wOvJ+XDOfT+HzoCsmOlBPQCkoBukVLtBgWlShhFCqJkkrCNsM2jE
Jejd2iE8/oXDZyZ9KCojwVnrPRGh5bep1KCjcxWfJOCHU0eLqMMqTb84r7FvTpYbWDfZZjAv8udb
gzVE72GtyKiiYqzrx4T8w//wpxjimNjbJPe4X4k0u85CZmRFx6O3I+DiCA5qICtLCDpWQKV1ZRSX
G/mBWh2lnD7w4MIZvfK14OhnJLBzJiYm5/zh5VsITF9mWkJRKu6a4ZLhpaglvgm+iB/LjcV2IXdI
1v2FW7KBbZR1Tfoc8VaVRup9SyOnfrcNeUDFi8pKwNxj/stjomNIOv4jNaIig+WaNHgxe+GL+qKc
o6bbW8q3RNLcPTs1YMVpzojJXoMhgGJXh3Tip9lPEQQsySmjHCDC/luEt+Yln8ajFKMxhC1JEGMk
i2esq6FkCZAnB2VNmHag4R+yGTI5y1oClRw91JlZSFzI4AFTl9LI5DGLSnMjJOy2uF0j0gl9kN5D
O3kRdOX17MNQGD2pgbmpLDx8kd1VpVOcV3g4VTecI7rymLqMYKTQbNeBWyrcvSy7F36qGecWq8na
nljm06zLisAQ9FAkvxdqdmj3I9SgaFc7pDqJ/vzmehkuW1DytzwhNzbebEh5nxS6nV5GW8pgUf2m
bqXINzLI3sg6WjAA5Ixt3x2ir7YCpzpS+wIxQKEpO2w4jQNAdmWMcv2+euxZnyrUAK8n6biz4x+k
R8ZYk+/lZO/Q3lnrUWv2LCGe2n6iWoNkbIlPeY19umDNzqEGRqYcB07afCi7ttY1slEEV6L5knLs
199ajiczkP7CSd+1X/4CSJSFJkOmfuhzJb1pcWgoiDNCp19Ea2xSLSfvyfwpwL5Gx3ZaMQdLjgqI
7kf/E3mYaMR6ezNyoUwDAeNs5wEt7+QmXZuU519Nl4qr1UrNRGYI60vWtIzMzGa9Kj8Y4o7wR9xz
sqIpok9UH8cdY236Yyj7FliVQwGtCstU/5oSBI05FQgw/fQyh1yGU3IIRt01Fnh+AE0rqvKIZRMb
vyYLmVOb9WWVdWbFa13jyd5idk8NzS80zvUhG2+eVkVypsGNE0oS96JMii/TaQUEUHStBVz2e3M+
LjsbwD1dha1Kom38x/J0+RP8uXVnlW3UB30lBeKAFqRubDoxpL17H/uBZPUkCLp7CD5FCQPzN70O
5aiY5G7aPXl/VRNOLutKkLa2i+OMkR5L7SiE/OWbhHB0ybjoLeWRXGRlUYjZnwgVe2qPnCh250Fi
t8JvxzTWR1Q8io00JDuolMJhjxdBVrgQuAaFxHKryayKieY40P++Wi/8ZKtrFaIJMIbG8ii3Lpe3
eu0vM+F5e4iTyph1DRJT/7u2imAp08Nq2sCcV4G+yg5PZk9fXgwrnj+k7a/emaziEGlLZSqJ/cfp
Yy/Fz2z3a5pw1si3p23FBqfm41aga3cPpbfeji1T3Pb66bRDX6XApoWVX1imIXL4PR8gYuIRVWay
15wZ2bNWtlnVF3ZsdxUHM1P4jwRLLqbCVkJCsYNiMCZq0Nl7uR4fKmR3Su1vx227xqNFr63B9nf1
82EttCkB9Q9qp4JA0BijyAFLh4QXUI/zP8QBA665ii9dW5eO25WXRYGd8GybVumA7EtcK0+80LeU
8U5gaxDylVfAbam/6VZFTh46YqOeqCXe8PEkujTlr+48+A4lkDFmy0TIzvgjLDvVwV9x+s4eTPsg
mmplDQU61zH+U/mVkoPdcfFv9E4HSnroSWOveXqry74zTWR3Sl3XtkaXzmyX7uG4uwyNOG9Eoeg3
cmKsPItMMFp8zriJ068pz1odbW1t9Q2jEtgzarsodFEbp3HOJCrvoSa8BDFUueciVupBEDlZlDgc
EcBnjtfkR8r/OCh98NULG45kbTnPFQoNd+O3kh812yAdTCpWFycNfAHvcWoLJdwWOQEdpQNDUe4H
PCKC+qly4W4V0/1oYyARDqTyQIMcleqXcIgPa0iQLi/15c34/Resvbwf3NuXoLMyNfVeLK4VX3EJ
ejH5yUeQ91kynm0UEWOLrXBUt6ZUlqkMUz8Jml2V8m6Kntp6BR0EYXOWb9gx3hshFiwlEWOmI/VM
org7z5Cq27Mf8/h8V4vOBs4rNkUwZi7RB+93eRHh2TpWhlqbXlztaI0LXG1bHk175YiGARTtE6Sf
38Cl9t5RuR9fSXMxShYu57BWitgjn0PkETQiwjf7apDRv2a1wKb7YvFHqMNYrUz7D4QherqorP1Z
A/kgz05uRoIoM8vAsouD0g2+e8ecKv72mwNyodryxaeXVwSDB8vyxCjIqJhe5QFtp9ItWyUss2w4
TI3igSZc+csiWmM+5ccjcMSy27kki7XZ+mKqysEFMvXY7652PutONd0Nzkwr6en7/rFN4oxwFovr
8gm/18rlaTotwA26JU6/4+/VBYLMgse6nT1I72+en9H29FiRU1ysUaHwSdmktKbPt+kJGCdwTL4s
iQ1w1LMuVzjko25KKzkckZMcRf/MjmENINGNHQlnQ5Y/gqHdbmhmw9tjDZvTmS2GxigHuU6jzeLT
l3OsZ2Ufu/sPTXeaSBjudJo99iteEcxAyJGW1ycD/3RXeYy7MZt49RVGqb0OhAdTO3IV3+RrHKyk
ZunJ9B4ktQMzkXKBuAE9+LjeBSU7KlzrVOZZ5C4OJHuGqQgbHT1DMeZO27JhfwplOyp8cDk0QxR3
LKy4Sz90uwNw+DiDhiPoWMc0RcGCy5Ja8i8mO5K+XHWI2BZwg4EahP6vfPAIbhJNGyegUyyzo2VF
8Sd28yOmp2bsAGYaDPGq3lpM2g/W7xwZfXICKOuCsep+uWpeDFDFosO/96JMGqYr3rGDmby/wyQG
RqZ4zddSymO9g82c20ima3tHnMRzrHhm34NkpUEqn7rZ1GGr8PmoviO5QBA1Non6LM4BCZhuvXWY
JEjQD0cvvFjI2/UDdYsSp0v/bK9E1hroXbVdP0ORc+zomW2LXago4j8PXOOkbblCuQa+JisX3WVI
2YGqSMOsQFqKzrfFHou11G++yOPIXbQcv/Gnj77AumkE/K2mZefcqMAkVNYn0v5+NloSgM8x62a4
AHa1yCuzVu+FKzXluIOAmSVW281swjBD4eUgt8uLOD+ShupaxfVYR2itwWGyFalgAy+Los9++1lZ
APmhAofAYFKCqoGbPFSZdsh81Au0ImoJ+x7jwXvsEJ/BhBMXjxUh4R5bc9nJu4dABqK3BvxHRMiX
vGH8rAe1NUPnc9RnX0Gdv4a6PmGjks4ST5qpWIX9hNqqhq/MJ+JU+Ao8O8la4OlgoqK8p83/YqVp
V/c4g6RnPuX5BaYFuRsplscXpyUXIN9hudxORxuEnUXk2uROSGLUWlA1BWg2bZjCMVXKynVRF3lC
GrCZhN6dX0hmGAEsC92l8b3RHwWIZatOEwNeRimI34TwPAkkHaE3js2Q0cymbuYOnuDguGV3hbvX
OLVODksCRTFoaxCuQbng0OFWJwzR3PlUswAuEIBr0biIgooNTJEVQF9cb/h9hQSC4r838mETvY47
2dYyC+XLG35UCU8ySiDKRqrFsymdn2P2Xic/EXpKcx/PeeN2ATKAadBLNCzycEFxdIr2vUjjVwHD
1hoZbK4wTkLQkh5AfRxy2+k3gt/5weigVeGspzMAnugiHrGLeeclSFBg3QnCvabSw/+qGxtpVs23
+8xTDYVKJSRZZkaOqT9/b/bHuPDxlpNLHCIsokVq8mo6J4hKnv9AH+r7jyj834vqAxjGBB+ZGqN7
wd7Nj4JzMIefRRG9mlVJjESMgwpYkbxp8ki+RvV2pQWCbp6oZsOoXaDGrRVVJ7HD8ycH1vRmBevb
JONKLnH88Hgiih6MK8bJOzLp0cO4y3TVod6IyPWrVx9wrA4EHu0N0DLg0myqD9BgiNEk0oCdxl7c
AxL2d1qCd4hpaGsgDQPq93DVKBuDZrR7s8Nvb8Xh7wKVFgbuP5aHFyq2Zz4L6/WVEM6vGOKisMWQ
CsanQr1qHuL15ope2RsdpzUu+C+Y771mOXXvGSjbObkwQv9r2foeqMzNyYJZMgb4IAv1G55W9Iwb
nVyRq/rgvEkhJ+F3ldN9AReBrK3O+oe4XIjI9h3qg+vAjFD+1tB1akZzmRUihklGlQOnq4AQVPf0
C0gcQ4k5jS4mXBii+eE2N1dQipo/kHRtdjq9J1ZVe71o8eqFSF8bs1WVD2kl9my81y5GtxsGnYed
w6k1gnUI73ZCs1iZwkpK5CL9Ym+SzUiJPV6HoocZr3ien1z4w5Oh2bmDHqUHTeTvrezFJOad3hD2
Qq1/w+LkYST7lWhsjPV/1fyflETYhp+P6TcFbuk9cha1hWqN5u907RVTsIQdC+344+G7YaW9fBkR
Q2mB+wELBkpyZpoV58D3qlwJ2V1yFn9KutmjDEdFRS8fVszrmbxcy6JdctOfKpNxszRIra3I1R8O
bLKcRWPp8ICw7Do0zmQSqu15NfgQ+dFkDwHjRfz+U/IqLseX+AKYm4rKBrn3Za7pQm78vst2x9+B
9Bt8B0i7QCs24vT5pyaeZssZxyf0DgZYmw7eldrnJmc0ssZD7IdAPHs105tg1fRzOehingy3aBBM
oApaO+Jxs5r0C7bwSQpUoTGEv09Pts4iUqjduZ/pknQLYWa40oS6PYcFlSnDzuvm60Nd8uRHUIAf
toen16SeRgN7JBZ6zF5y01X5V65R0jV0WnyjCbKLvftksEkn2vsmUpzPzvfwRthOai8hubEFKI+t
UqudSRWBO5m1QQ7hAoAV3lyuqP6xuhGhNtyHZSgES9bHK4zmKvAODZao2XPfg6SM/JoLz6fMG09j
tvInKoVqttyg0rw6sp68/hPWYk4nkpxX3fa8VP/HuN97y42qaKmRYya+jMZAwP5bY0TYlezzR4fA
Oj9owyDAcwe1X3dbH72bTFZL40N+T5cQL+SEYrlLBG27Xkeqyslg2JBuDXqDSQfK2ECQ8OQb7C7a
Jkmpx0aDZkRfpDNUzJAdZ9pEPHlsfEwiBsIqRnc9H5ox3cYserFUBtym+AqffSh/v8nZID71J4Bm
sFCwk2fEU2UdwA31C9hPp55JNFep+wdg/2NEABqxJtnETNPHDvztBcfGJFENnMq0ZVki3nWPkwZc
tqueOs09NbiAa1KqpGNuTJv9HefqytPabDsO6LUtWjc2KP8c6/rY4ov7grPqo67lR1YF1hK+FAy4
T3GH0jEw/dATsWxJ+mtsM218FrQI4BmKzjY9CPLaZpesjNamCl0xyaC+x4dVl2fYjeu5X+RBM4L6
J5AYrKwjTtaMGktx8BCyjpNDCN+GDpmpQU4REbvtfavBGksTW1n2kXipAdBfuA58/8elHo+uvaDM
LteyMeH9kkcPnbt5nm6gsLUqTMjgT4P4uSnS8l4uwzj7uPhELKeNQ1RzDRe1X9TKYlrCitkIZ3P2
fAZceUgjo8VioSXq4zpMtL0osYyPu4aXYsheMSUtNUN23N8MJUBv0u+b8MwWSd8/6LAPizBPOqc7
xGz3u9VlfZP6ngZaZpdKozEF7EbZufcX6+Gk8/yQeRMBMw7TTk/1tp+BeE2UWB+ylX7IweCvRKQg
3EosLnAwjT4r0mj4JxIlCIBJ6EroyyNsxZ7pV5yQNTNrNKsrwtXLiMwGJ4DTqbIxmujO+SKOtDNe
bjJycZTRDZHiXDKFGMlNxGZofkCsBcECfApOx5Na7w8zvATKNxbkKXEFaliLU/eudWNrumGXdEpg
XQMtod0NkJnPYf+wrYl0jIyXrm3AYW0xEfg8imyI+obuJZCPFe4mqp1NtvtaeSzct2YroEjbQt09
8m5Dw0WdyVc1e1d0IWL9tv8jYzwZsCwmqV262tEKWL9bQDL6oWdHPtAE+QLMyIuXTEBMV2Pvw/lb
vc+rW3ogFs3GSAN+prtpSefI2ZhfANz5K13sd8l5D3RkCoJ6NPN+r7SKdYqkXkM0X6h19fixWkht
xbIX4dwbTPOP+3iiXfHRRHtDaLebzf7UoG9VT31MyNjxb3fiPQxnHVpPGpHQR+dZtnMR33abfCSl
QMx7hmkunnWrf9Pft5awEfYZ+c42qc6llV2ndbsZBUV9BSeSb9X33z9HLl31okgqZTcC1/awwAU7
NNHwMKVV8R5aNHMGm0DoZewLaZDEuo+YnanY7hWDbVJ21O/KuqKnToP8TvoUdi3TWbOiI2x+BLkS
XT5yd/kqRKDyDYW5dbmiuizCRG6blF3Ih7aRmlARdCyaXhQGNgQQyfvt7/dpzD37JM9XfE4HkrKc
GM2JwGM/hJ7q0qj9kVFnQnaEGXneh2VYnSimWS0TWf9QyBzzcrhKsHUYjSp6oD80LsVBlQMlBA1b
Fe3i5VH+wi2WwosFaRxpKfoECrRJEDE7kng5/IQSwXh4sdp/NM6pLGS+TvpX5AB/ocAhJ4IUvvgs
+UI2ZfAJ/z3QQY/hf47z1OiViXZ0hkMVPk4v1Uz/fKI7ZFDYY5zDcNF3WczGFLSP122/9y9e6BqY
19xjgrTN/OXY9pBYbZBhh3eR9orxRWW6KHxwxp/BIkfVpdeN2X8vPEooAGRlsaLh+r5lY9Y9QGPu
wqxx8Dcqe5LcPu77rjB1V3WJVi/uio4gS1uv17UtVUkaT+48uFYnD04Ood0ZoUMp3+VKG9RFdzQl
Qlgy10XMeCbrpH73bbAd0nFMS9RyKC6GMszcqwOrfudLdRPFRYHkyhuR9lXE7a3zqgT+WZZjNa7z
G+GZKMVa3XEoCDq/2FSqWFBY6M7goBLvRJHwA54Qb2XvjW59xPWkks+zSa4YsaCPvm2IzAWWNpa2
GaQiFbEqGQ+hfxqbgb6GXsY+j21qWg7EnTzHJ1D9DeF2tCmXdjskWmoaFNaKhxK1aMo0xm6osT8/
NTrNozoe2gFNBUpp7+ELWUTunJl0Ku7qWDJGFwF2VlzvSfaYLprsiuq+795xJLznTNRrn3z0Id8x
9OEbHTsJrKaDNDYpvUSaOlDtqPHmyuKT4xlf1ze9yLbFiEYC9gMHHGfhjCOK2CW+jA4rZKStyuJu
65kllKd7CZrMHLfeVVStu4YkYUAVnMn+tXrecdmc60s5uL+ZgZY1dQ1aonH0ug4tonySkcrLx/bq
+T5h4ZZyvQOL1/LCSFwZmxJ8GGVVKPrSm7Du2t7KwsxhZP5VrDmx6iW3H5FoN8NyS89qE8XQPnDL
d5mWnp9YNQ1dUOxcTcV0UsRHeIA2tSaWb9WH7o8b5+eJVlZX3KEVv9vZjj/xd3+oNdSID+SCIfvU
qxDRtlPFXV0N9my6Dofc2PizC2UoDlRMrq0LYnZVFsw3/BoZkhsQKwQZifzAa6Rfpv58Xt7rPB53
SJj/FCyyujzYgYvUUpgJLbHqurdBYBsOj5Ghng80CQuBpNTfJp7aL0BeGrrE2RLcZPbSaHfw40CR
7Ia/jfIWrlf2Da6wbENbp/GMlvMwZINTsJHoOYvwhyBgRcwuexQk4SxF7k7KmFSSP2V3AnrSZ05q
w8pvPwo4C4eameCSC/VnNmkkc2ee/0W7sZUYWmwF4pCkMBKXuqQbEkF0gSyfLhDbEIUHqqyEm6gd
MUZ489pi93i65wuAV87cpniY1A2wRaY4ywYtd3a5kK73uQa4eOQ3QbC1/5jg9rsWwCZepjC8qix3
yu4wz+iC+8CZnjfAx9H6O3qpsmfV44Adp6Xev3wH9Xgaav6pnK1fu5dgeu9bF2mRbfCRN2tFNj63
A52mFYPXEtBOQSq9VqLSlIk8aIxQpZF9dp5aPPJ88ntiAqTIeE5HnLKSSahdAWfMrCg3enGQL3Md
F2HmFAvPlGXlYaKbkHA96Wej5w0uiMqDlE0/vyZCrUTy1vgRWEk8a8cGKv6PfFW8FluvRJkIwhAQ
jaKew/B8USkLdjWO+A3S6e9fdD6sk6DIepylW+BLWMySYCg8VIVLOoW9qQLQNaxjBuUulD04ECdI
eQw3EybEzu7TpEjtcc0JxWgUq/N3i9b5ovALkAsbLqP6xtKxttoUvuam33z3pqKLse/Js2jwiBQu
ay5KprAEl2uQEXclkM0vP7Y/XD/tKfTzI/IV7AQAurYJpYoEhogH9US+FYASQPa6dUYxZP1KG6t0
YNV/X6XaHWvahmhhiNVmUTp6EmIMgGAecaxjJp1jwU00ui8mfyjjhQly/+7SK54O7cqCfGw/vcfX
SEHmBH5WDE9PJo8TsciNKEGMV0TCZxnfizaa3/IQijhndPuVPWyQSOgKkzRQ4N3ALM+x/1v1U3/j
QLhyKq9nwV6+9gVz4qhTQiuyOABxcFJESyxkL/qAneqINXgNCbX6fH526/x6TY7Z4iTQiHuDgApr
b7T777gPYJswRgfgGB0m1pfoDhpLXJPUj2hk1rz/81UeCdb3CIRv+Efx5U0YOKUG1/FZOirOwVN6
inJPZUhRW8dMMN+hAso0m1ZZ+ZRE0C5Kh9HaV6HHFwcdgb3dGHsEagbA3JDOvuFPc4dTjmJ7eU2i
R3fCz2Sx6fI1BneyHFvJGabdf6a7hX0JvkAK0so686Rn1VLLlWlcR+QswEdUPnwal+1mLwMJUuMC
I3zJtbeugLFw+K+F/dzGgSiCaJpUevIpSmnXOrnu6JfKhZvrrEMGA5zbpbyzebR9LiJNPNm3/Y26
OJJcGNGf6roXjJ28qm/Ye93k5XQX+cjMv1fPTpujwZxkNm59FCtpoxPeVhAubhFtqYYdCzMi+3kb
TLVr9L3QJAfVAuKPebgOyNc9jVk1LsDLMBYSYeKoPMpE9uEcdZ5yjLORx08s3S07B5Cjh4Xa0RfG
AjBT3oJNAwWug8H9SLHJa4DH6PgbUvOnUVqUw+m8mIvmv6BfEcXAe6oGzbqJO7QHhhjNj6pdOqkl
X3ng07jQpx5Y+4oAxIVslE11rRyJcP8khz51EsT+Oq3vREp+27Z+ykbKTXNrrve/dPUZM5MXHouY
1lJmmBuoEo5tgJV1CclpLlLbyQ3REpW5hKGOCOn4VrLjVBt+ntxI9vq0RNcUT86MkjdYW3Eyq2XR
ale8lNpJyOseyFzKtlxpzvnBWDkhFWXNgza2Cv0YXvdhAfCfnFgdhNyz0l4MF8Pa7dNNRGEwjcQM
JemBntHZFxq1GlAQZ+LKAyWkVHOovqBtpjT01Iat5suMS5OPNNfSgO5e5lCY+F7zuGSaGTqExVH+
27aP611Krly6AD7awYvbMUR39kLmzhafFBli5VZbKCaLbAvNsCQY6upTle5RPNNIQtoaGkDiUVSi
cjW8604TuWg9yPenZP+pHyVEc0zTVdH9/AcoYPPGBVTr3H/Jg/mVZ2ChwORBtBw8r1wCbMenaOxO
X1Hf6pWeZU6CFLS+Me8rqv3XvUR10l/MmO4VfImcTnGSO7Z0PEkHWqgQd5CvDvqFIXJ/mZgpjD88
cwRDWb++Pw8rCd1G59bcbHsPcxb+HxiYZCINyP3kESNPWEcGHHhePV4mGwtYT+N8P6hCEIr1uypJ
Zqw/QLLHXFbbj8r2ty5JY6XhVQBN8+lKr/mnap4MIna74L5Zv68DKpfT1iMjyfTYXwdG3K3s93yi
vu3P8IJJwwgA+QxKBajaRQkrmjowuhJwvN6rTrR20nFCZJndIhKHMZO51Sik8IEOTWkpyKPxPtUN
PiUlp8sg1ixrIFEypcjQtaNATTZqR8Hg88mbOjVImVToWSl/v7DvM2kQFvhBgULrRfzNTHPBde5G
0rwgDwrRlHH8qjgD1RN5R9s8FLbYUf2ZFX6X4pZCkLwudoemZbnaA8ykz5eXwLeUFdbnnO+8YOZp
Swc2M7AeND+5zAbBuYF4KPgjPCnofS4MVcihkwPdXOBlfLxImcGw0aOw7dWlKF7DCwaBWE8IRpY6
zO92hPv1bA/8KKBzUorTXvki2MWeG0LAJGnBmeNePDaBdfXkLUbWsNlCf7FxSe3PrwFvjbtkcENL
ZmFUiDWS343dMJvmCC/1T5Chx0a3JFtkNLuRO7GilXL/9xOGedaJU/ZoGsLvaF1kVMNS+R6aZVec
scl+CjwMVcNxwmqNsvTn3nt7QiGeIJiwuBymrKdijyfzNWen1Cz3bZamZZCAQiQufwgcSSU6YWVv
qjP7a7mnFZ/QDflipjoDgjD9N3IqBPv1CfEFdls2Ridt3VgbwTpRuNqQRzkRPPSRdXUDK+v/mNa4
/rPGqWF/oGaKBdyEDUYpZIKeOwg04ofMrWHXK0H7hlprxNCVEZa4/HXPtkdx1LEI5qu4gY8eEEKV
WrfUV7ORsDGxqmkg8wSo14CAHauwweVXN17y5AkOxlsJwoFX2TGwLwsawpT6L4yN6YP8OebBwJCU
VtvxQHBM+mpVa4h/qlAmOiDMnnBT9Ly0Z1eOOfFS7dPuoXNyut245iwbyd35TAIjcn0zUe5j3Ppj
SOxJkPL+l0mvicmKBluha6JJcw5jKrcukIe9Kyg9317I/ayWjrFTa6FO8qaJ0JxTVQ+8OZcCYEzk
GbxEHYggNGvq98Vmre5j+X42JMJRFVUt5RqlXTotWi5YmEC8y0v5Ln48MEfusFDgy8u213JoWGQh
fhQCTU+5tlN8YpZf7bQS3FMi44ATD5xfQW5aKb87DILBU7lj5whA3A2eosWFqE2J+f+Pouy61XaJ
Nb6K8xklMsjxIPTvo0nFy+ZoSV34c6us4uA/9Wny1gpSWL1inOHo6LEVC4nxQHl2CP3K6ae3Ull3
0F8jQCmC8FzBmM5SfPvuEL201FZBpwIbn7uzQUpPBb0CtI4tM/MyF0ZW7+oeI+VVkUmyZxUaZacq
7dX6JbUBXn8IEcj0MxTEUZEyyX362g3RzMayYI/m5nXv7HPTdjqpodllDaWTTgXtmtUEGjdOkveG
hs+1YhpfmaQKnY6kB1Mi1Bt3XLv1rJcO2h7HO3AJRpUafCe0q4r/IHYY5AFyUBjNmsLR4jyQ6pt8
cNgenG6czL7oTmkme+nE3ewp7BH9yA4ywlQ1cvAdgkaCInF6udFqVnJyNsQoPQIW2I/47H3swL/z
+zyEDgKa2oMA73esLuDoWu4teVt/dG9Qn49zC0hTOh0fWAHWKNFRNgmZCJzfgVrc/7n2GDiSIE7u
bRpHQmqsH9svJG/XbQMHt5NjLbgMwKBALjA2FegrdJu45gSWvPnWLcK67MdKcgs/uRYpX8B5qBu5
9Bd0hfFMO1LFZIvF2n5sIv8LhKWQ2FY+qlCr+MK3m9/iPFGDIu/lgxeUHuqlqSOslwRIkM7E1wEV
X3q4Uw1Elklj0yFy0u/TJbuV/FSBfPUa8oAy/VJ8nfQuP2E7EZRzelQRA4W+4nG9J6DzvObvhpGB
ZXS6NtQum6btZIX/WLFb8gOFZtZko4kto9AH/OXBgsfOTLoT5T6sULKag0Ob4OgCs5yYjQry2Svt
wXE7ksvmy9u8r69Xl5EG+I7WP+6StGHUuXjV+6ZxcyT+374rlZQR7wFRX119nY37/Pkp+xAUrcrc
i7RkU7yLNoIirYjGKAOqBuE6hjg+fHwTe+wg4fnhYvRH+o8hirW3haEx9Hs8u4BELrEJ4WcaAAJk
C65SjcndfIc+r0smIL3pK9k0xNB85QtXm8JHX4P1VELVucwyvVOar4McsJ33rEyH04ORMSmelZw2
5UIw62fUB4LDX9jdBuhARqlVUUFoywJ9Ia5nFSMOqM4puaWS8ZB1ZgdXW4eUyb5KurbX4MYhigK9
r0GzyLJ7GWQUeBESCbj5l1yZ+v/4ja8jZKjNikIjos0cLCivKA3bngfhpZwY2qWdwinjWQgFLKRq
kaHtsJg6XTG0HNpDtQ42kZ/0Ik3JlZ1HnV46SwBjMJyrgujH7aWrckSIK59ZEOdT03h7BX1B6o26
orOLn1tKbq81eE0u24m2UuZxlgOOgczTyswqcwuQlmCjUSIofOrVHz9DcmHMVOSn6+L64EqdVz8x
hxLuw0RRXBZf5gsKznoDgnkYJI5ZJC/M8Z1wFeopxxL3peLJwYA037u7WUYchdigSqUEPlmmHR4r
Ld64ODZXZjmxa2zV0UlbgT2i+a62j3A3GYXDCHto1IZIOp532CnFRDmCjfBSHX/YgHKGKHihMppd
khcYNeCuwWOLCFPmecEMcO0EPqswZRILBK7g4MxLtxGgKHztzDP50D4Jzx+ZwluWKakdjRU/8yrQ
KfPMcnVBOqhLsh8PwCGAgB9iZ8A1lqRfnB/uXTd0F5c+ojzFTbvmTxCZzF1ghUP3dnBZV8p0hQf5
gU57s0SFDZkAznto7wgoljS/RjkZ6x/gmHpI+e4YDSl9P3U4IGdUi4598lmDrNN2jKHdpCGGNLuW
a5G8qzheq3Xj1/eaW8HWil4gdWRJxeDfvd5/9oTNQHH66cadfVeea56PZ9g4r7dus+fJ5Brohe77
XMj5Moidx3gBEivzEFA1SCM2Sc+yc5eNTJvaRkQQwDpjJSLHs69u3V0iSv2rHhFRZpGZNWxadS6i
p/tGj5AB+ZYCrTjnNioHuNNMdyjUgLDkTPU06NRqXNRPQKRSJ3RGtJo+mltcC4LxeyiPff9HtE7y
q1oTxCpJAGoszykxgx3w9b21mlo5NMSFlrw76a3Rq5wC0h57j4zUalTdT2FZmAeFh27ftJDjoHZX
+QwHBC2kwnHkRETQBgn4eaDr0mdYR2XWa8jgf+CNzL1mzEfyKlZqNYSHzJztseQYSxvPJoPIE1wD
s0QLPNr1eNXA9mic3LU12DE8nwm36E1HZz+BFhHs1ecMxSgrF/o6baZD8XO2/ksjemdj6+xqk///
fg0G05v13uNebkuNBy2p+0l/19ebheyPtOWeuFfpY5DoNgYaov9Naha/djGDmrpOTp6ni7Z4b4Tm
lFNdmsDWgOeRIoDsjngpMh/+aDlg4Tkp5OyQ/7s7+wpPdAAyToco7b/of6OwxWhrQsqz/TJNOdEp
8eSk8i0vrUQLPUIrwCSd9EMxL2xuPWBamriHpZzikelsDItTKdGurtFrT4FW1RDyMVclGNEkUXe5
wdZ1U0NtYpD07nITtUUhADnybGU5BqNG63v7wswk8jgQKjXeP1kmF+CI+q1V9pF2ybPlaDRVyzSv
wQMQXUEdUYGVMudix8Cpxc5dvfiFeL4+I25Nm15uSe06+sAg6QZca2m3PBrdU4NO8+q/dErHtoJI
1loOXERi1XegDTHw916snro93EUonAbeAlAfpQ8YPovxue+raqWCKXXreZApK+4lkMBKtUuTY6aS
5HGKDr6ed2CuXjjNYZQYtdYPbq5yIfLFcXaTYTfTOsxWat9Uq4gqlcUBKGJTvLFf0p+CYVF6gv/C
PMiH+NeOlC1xbzKWZIVB+6KQeWzgHWsADnCZMXOntNdRGIBH1Y9NlfsQik/IKdUlFGUVNJ17bHXo
i1FnVhay0SmPp26uL6b7Pet+DFg40XMTpy2MAV+p1LhP3hGoMoDF93c2ybgn3/n8OOyMeAgydJC0
qHMr1hW9g/LAtAO7+GSLsvUbKI6txNg8xwcpskny9tgxy2mJpzWeReZrdGeJHRGGK8POupt/eR+E
ShTK7cYAl7hoYe/3HSiXBLSpTMwUayyUnNuBzYX+Gc0c9K0vXJElEbh5cK545ox0kODvf8ytWpkO
L2cs6iEcfIVVTcscReU33ItCoBMzIYmmJjk7LgPtgX5C28c8Yx9fJeFRbdVYHD852/Rn2GpDplom
e4JmDZ5yT/BprbLpeMfS9GtYqL8PaAYBxpJ/J2Ti1rYUyTSXnoZjoEtUjocK4gznOUBxgHCLlPaI
DdvTXQggWxOANR1+ipIYLTLsdwnBEcrJ4edElMeA7e09hkV4tiN5KfAXbXL2sfQWJLkOhD30GJtV
W4+1DDntpHWua8+wzQIPgml7Mhfh6anyYJqohaqdzGBZ4AtilFY1AKHkmvT+xTF+qjfYYcrKl7ae
7bmFRtHvlbH+QkOPJVOc53a1urlnAyJ4LJZk2KEKmPV0mqbMaFAmbLThaK8uG1BpBPVdUXj7+HsA
OE178Cvwkm6khUBOSQDmyMmFKwj7X6BPDGOAPyLl4pQSI9JdtCKUR1TXPjJ83E2/yeBBbUVl5uPX
PnCm6RRtexySCuL6Au0gG7TErLKpLexBfP+Ox+UQobqBb5OSBFnSKSLxGJKLayCn9X1muA+/CoxN
vURMhKtNbdeC/oUoAc5tXb32GPf6xdTXeMwrO1TAestyj4nj6tBGMLqLn6WNJwEGLaMhHhDW2us/
PPhVJSP2uN127dxpMXBoINpYVDEfFB/migfqBU1fG3Vc2Q9YTLdZf8d1xjvAoYkqkxpjhClRfWnd
4fuMKQJeHdPVYmkkAyFqU0raR1/DvFXz+svudScpc9HZGqCZ1n3X2l+H1mWQRnTnI0uygbzv8NEj
zsRXRKU7ph+0vRYRbBheIi9NcHiwmKT4nfABtOdUS+NyhiFxg0pTREjyO2q+L3oYjik6Ef6fsE3y
RS1ZThwkhD9T5U6Y0siNw9nQs/bUNpjRYZ32m36MvP0gi3PMpBEDkFR6UHERROdQzCstAQcS6Lyt
x4bi5FhXqdaNvCDARekv86OvjCjfwqFOZmQOWeUQLgn+YpKYxFV7+sTZDV4/YvAdmqJ6EeEuLNqy
9OBj1vT4q1XQAVY8+8Mp87/iHUb54djqBqhdTUBdGNuKIxbKuv9xiYs3+K3pDuuzUsRwkZ7T+BHx
v1t2ZOo2+oVyFmaBiPU2OFnh7XUggGw0wT5NbKdCJJxvaUCyeHzoteCsZkC1xNICFzH7e2JlvSZY
/DCom1rdQAuauE44WHGDI0LEBT9f4cyEdkI+F/wGNyYz63K1O/Z6t2ShBabsRaX3ypJVTFAJKzRu
pORk8tPs6AODL+vm0hL/CcFICOjRwUrPOtA0S7XQZS9wTKzmL8UL9aXykzsR6+f014b41Kl7iGFb
AZetHSH47CQ/wZwEZ4P4xo/3IMZ4sCFm/1rE6PrYiT6HvSGx26iAvTX0BLadJLAJEV9BEwQUlRhw
imuWZ0eBWyT9BjdjRIO/B8PcNK8loGsTovkBGE64nBBnqqHjNCCNmUSYwzNYZsqRXPVeokGBMSIR
eOmHvJPCTqTjQ2tscs6bzZbPv26Bh4NcW6pAqy6nigR9qoVHy1gObXtX8hgkm9FIpaVQ7EF6qzyU
blCSWANQqIp8ghQY6OnTvivoNVqBHfwoGSPQCvLT3aagyGa32fS00bP/U/9ejCT9ULsdybgBHEbZ
+OHT2Xxy5Xuiaix6W3U1XvEfLN3iH9ySXg9wDz87ZLXt7r5LKtZPWEYUwtRIGiEG/1zZRL8r1fM2
zG73jtzwbHkoBIOFeiAFJ9QewPl84/q4ouhH4XGg35PH7WmIbNlz5s1JaDrBa8jmSVhvjIfxrBoK
V2xlBJ9fJIcuOtO6sUDft1hNIXbSsxjnlZVYNLqzXCRVAtJ5Z30AQOk3TjWvhWzJpX163USAWEyK
pPPD38xDNdz+GHB5xIDkCRbtgjGUzOMlJQAltyVU2VtP6Q8RZujqrbtuBIBR6PIWkn0ZUXTplSeR
59m+wT52i7+0ceBnt82kRc3rVuvt3nya0/4RoRf/ut8nMtwwrRVlgQYZyCKh/0iZ8sxo+jTG/Rur
V8RJQPo0dGFKjMYkJn2PtT47y5HFPdaznLTBaJXam5f7m0B+xJWFXZnqjItluxWnO7zx6D0xtKUb
3Egpgx3ccq7ZCpar8ehE4VBX0lHXr7ZJOqAwKVv72gWNk0m2aE5qyNbDmoV8hymrzFPvlP322TCN
YKir7rXOqhodRXxcX0+PCLArvFx1o2BV5qAMnPSO8+nsTHvZJ923f6DoU+cVJxXp/nB/7kai3Lst
p9QyqRUZS35AzidS7qnpv3M42fQmmmkFLmW/k7jevc6mU2hP0dsyy8rtzDPppjH4a1V3rZkQL149
IuOsTXejrt3+4N1zbRKxkdc4qQCQURLTU6PRw73AwitA8RS4dVdGYcr65Uv2fd7QwrHibvDMz+ok
1iA3i22rcxhNkgi5cGCyHAh+yGzpj4i10gJbNCxZ66nFFEBw66Ed8NrlXRPkrOxg0QqCJDgxsy9q
qDoqezY6MT8w++zfc0Lb7bvMndYGIxOec0W83Jf/GabPY6l+roTRUSO4iAoadEiIHl8U/62cximu
VapCaCB88k30S93NAV8znP7Bnu07TpbCYjJNWdFT51BGjd0qlxNQjhV/QJiMNsMmdxL/Z0PklSpD
uy8iVHKO1lgK5OWcU0woO1J3WU54iaOXqWasffslBpNSO46SMEpXs3tN0snVnk3pH6XvQMChIGn7
lEvuZ5g7WZaZg7DXkDdZ3qrNlQoB96GKhdmqHRcm/2fmgaA6gJ/Yu9WCN/cY8O4Bwcasxt5iMnak
8Ai5wGu378ZBfX6IJ1J4MZrQ3Q1veHsULksy0uYnHAdUOiUXPZAJf0UZ38ocF4/pY1tr5AuB3CO8
Gw8xReu/9iZsrQ35Yz/AglTBcKyRoWbwK0FAmx37KfdZVnzk/CvoC9Qwl3O5VF3gppd+Bz0sfmgJ
Tod9InBzu1/suVvVmP+3bAJ8kNuUSDSL57J/fwEUqyAT6y/YldiBe0rNx02co2Q292xzunbCMPYk
Eblx8KhhXQ/hWJD1ZYsNsjH9UGAybzDJ68jW3fAA6RKTAppWGQC2uNgBFyVIbuPnXR1jLcy/L/hq
DofDKFQAa1LaXzCZSTwwlWR9DPjChgczZEUpV7ecISneRSqmPGJ0US0aCHBLnazxGPdhoTSNhU/k
XJd60SQMMlH6nS7lSa2eCLpD869ELle0IQMb6rzVCNMU8orSw/KO9s5mitRFTVWxMNDL2j7G7fnT
wazg/LdlnfQ+qOlciRO4/do6sMU6pPxkA2Nip6lmgKnrFEjFdFFbh1mVUAfzSx6NK9CSBOFUT7kQ
3TDhl3K14wWWTYPNoDI62rliBWCrLzjyLsfYaoS2W9cVGbAOghPfPsGbgvoB7OnE1Ce5erLuBBk2
3OBX8fnjSWJ1/i+m5l1LQg92y8JAXt5MEqV8KPOUs7P7bDYZxwPWTa5E4yWps8r7A4IR+lX+T/gC
5x1f+5x2Kc8ep5i5tREsstYwRmf107Zt3THI4t6Y2Px3XtWuYHF4nlFZaffaPoocl/p0f8DSB7rv
ygMJz5h7eCijwjhIm7laMqiehrm5+ssf/IUh7CzGcdN0SPsDUQHUhmxzVUVmzBx3HufZfORwIZVh
4Q3WPrd3N88V35s8ergYul6syCqnMGxNV4HH3t7cIn2okkiQ+yofmFd1+EL3ZjH/GJ9dSLelMr4O
SIdvoaif5uvzaZP0ozhE/X5FxVXLNFszeSgRWcE5KfIp7uSkSrtyQyPGp2IQkV/jmg2ujm56e4CU
spUdv40D2lJaCHnVl9XZcejQw5E1jS0pSe8tPhmHI1y7ICw5c3OKHoAVL/KKsVoEzqmlTk87VZ/0
A6T8TtNeefKiqV5vPZFOoUGFrazuhV1pdm2R39Amcq/7usWTd0Bxa62rY8+/qhBpETmbfXdBnzFf
uW72OqsRTEbXPxD+3mdOxr4VLLuVmC+jaQtpE5dBmcmKKnqh/d1qnJkdBaxTngzzENy+UjplVcsI
aKJmYM6ISs6qHlg4Wv9s7Cv8DygvALO3L/6lNQYJtDG6SPCxUIuitnOG8q2potNNJj+nrgl1FYPe
d2SLH4lRZXk7AE0b5BHyVTfTy/iokWaJfL7JacqDSYx4v84gCsqzB7khA5XFiSOYUXJNnijQzf9V
0Eqop7tkUgUfvVs5ZcU+pMUwFyxDZ2UbU8RjbD84GZa5MMMm/8ByrviYieLmsxfCa7Clwki624sp
xfwdXt8qKInUpfuDhl1G1q+kQghjtuCWaQglJ5huf0KnNyODcmq+tCZINM7DJWQd1NRfi85JLqTv
UzPZH1vlbYmgUq/yuWtcnOdwemM5ZJe7tbzY601WMvT2TVMvet2FxH2pC25LRVEfZcfHaEyMFM5s
SSibF/fkLfm2FrHgB+SvIQPO6y9Aoj+/wWX5OkPXdneD3kEdJzIZd8nAcO90Ob/BrisgBVrA2ms5
KarW74YNF5Zs4O+l0tKk7g8RHwSHBQZdCog3kuGh5fHPkfnB0ADM9vyOaGKc+8loPcdXVuJ3Hj4b
hpAgfLr35aHoy/0YmPJQoneah622xrRgBKL4ansrdq2EppBA5ox7l8oM/OvOKU6yxQEsPqv0Xywc
iVD8kNS2UOk+rhfmfsmTrDjKMVaXfEFu4bcf5zzYoNqdq+aeFgZ4hI21sEPRezIIY9y2RbsIns6x
MpNz3DU4HUIp/lV4GUQ7Q+Wb8oYTM662XKdSupgZ64P2AVZg2Kz36DOJx5swLB8uvYuc3JhiU9AS
qu77wgFUObJZ9eR2PZAQFQLZ+Xv5o0odLgQmWWJLEF+0xXaYzXoDIVStbRLT+iw5fACMK897r6xi
n3YN2e5RnD/KVsuCn3iN9t/wpd5Y/uEaCo2F/C3sxqU9t3HAXGACllh5kG7ZfKs2r78jTbJSXBgU
2PiSabIJAy9wSuLmvpdkaXV5HpKR/tnHYjMSHwEDtvHP62sPQNLd8lsSDz1nOQJv57Dak2VLknhl
dk5GHzu98S3a2ub6/LyYrPxlFl0RrpLQxUVxF6Tz8D7SIF6zSB1L9yGYDRr255tSXErRP7nk0FVU
ReFd0LfQH2gWgmJOKV6ejKa3WbNDRdr4zuIX36zdzxK03HjHw6ty+zCDG0crV7y+hiGqPYBlRiLU
bKO9fhjhDk0nlzhVbO4ZDqLGDb1PURL7FpgmPekV4/LlP3oal5iXbQpghsWjimQWv4EGTVRW2bHL
uFcCcGbCkw8QT5vbT8WHWcfjRAT1XVAKkQP2JfiUYA5JmtAsFX6Sr4ji3tzwI9OFH5xE7CuvPTXf
oJdf2+BXp9wVhjiONk2vNFHpnXtB+ES4Sytx96y12aPXn364m3LuvsVgSYCDBHO2yoKA8NeBdKU7
RymEeit2i1+415oMYfRHn7AQFN2y9rw2tZR9M6QuDADQhZnaeMfCeBmYdGpjmiRohanIlKCq/8jQ
rGchlCEyR9OrVhnGGD5HgcaZjNkAi7GJ0lVb5NRLrzU8IsHsmottIkjD8eJY2yo68uf90Fm6UyI6
taHStPpPXDDP3Q2+uU1ntwwUTOr6ZOck1WN86Ql7QnaJOO75wMjlzWFYqDpbQ8Ep3vexf5BvZVum
TrrYfW25Wk5VDLQfvQLxyGHxVR87vXC1snUMs+/Hb88yUq/LSvK5DiJJlDXeGScmvwCodVc1KRj8
Lynm3JlczLn7pzLJuJM2rQVqAQdUcG4e2h+gF02NKKCOixMy07QsTYOMaeUVZNhGiYH7vEXKNbSZ
XqvvPkR7BaxqH5pjjLDutfoknf2maTvolq+99PDtgWyyFKys2Xq0D1dql7Uumz6udptHg/aI+Pv0
BhM1Ck9B3G5ZYGypZxeKOGP5B/nFAsHs/MJFcHrUY9k0ZpYIq/ONCaoPdJDApqHHqSQNE3Cp0i1J
LOfgTQCUQmGyLbR07dhYcwc5kHkkGGq17hKXEzhPIZCqgV8oR4HMh9plOy6f7E5GReOy2hy/c8bF
12+AFkmcPmiK6yqWNZl1r/UI1VzCJ9u+R8rlZPN8+/FWHMODQ+CD5rWpmK/XtUgnOPdFg5MEKpOk
nX++b4tBDDeFwEd2r5mjiJy6MOws80HQgsRIMEzkhQPq1ztB3SkGTLyBOoqN8xCFxbCrN4A5ZENd
GsRNkfJNzjOybMJUpUrUyXLx0YPEgwP6/7asp9cF6QI4dddqYjRo67cZCkD+sZMGLlTdOydEEfaC
ivPfNwlenKMzfgnxXKn/fBB9uvfBcY1+TpxiyCui9t/nzpombtBpoJasA1zE0ypDFln3yEkY8Rvm
nC3HjwwjTB7B0/t3G/K2W9U6dfCrntuQerRNyjL7LS7mhEIuhGWpIVD7mpXKHpf11lvJSqdh812i
/FhMQW/B/4Y7ZLxEiY/ypQ2+/J+gsqIjw7+RG6Ax9oLbJsDfFqqDjZqDhVEXP+2wso0jN5UHp4Xv
ZgCII5f1yA44/e5YngvRkEepXtSMmE/ymOgtcjpqY330YJsJkWj4/rF/gLLoELNx1ogaCfv2aNhE
MLdg6cPhjWPhIEh13aY49sNm4SkAvgEJxYr3g17UTJAgRtGcP9d4yGoRfP/t8gUcg9XAFgXTwOI/
4dXUaIt0PFxFiYn6FP/HOQVPVQi9mWixjZBTsvOe3r6LKDtJKAKrO6X09Q7FtYIRfO/K2+ZmeZL8
ujON2giSFiZIRGBOeakFAWZWKUnclsM623d1n4JD+3/bo2Ke1/4eHUorxoIpIBofIakOdjscLb1S
sT7qj4uhPZ5QeYY62sxyLbndRvh4NmXUBqPa4BubQ3CkxPYyIx3uA+BpcfzPIqaJQiXQPxmc0l/N
6jyuGKQzeFDpoblhiLAqMsLwBFlfK+2nk7zRKcCCMtm2NpXlDzOcPrJNr3q7y5hRkpimK6A0mY8U
Bv2bxMc3P3hFkn1eha1dwlW+E6OZz0jN8dg2eyqYPMUXSR9ixc+2wdlgJ9a1V3em04D4EJ5ZGS7w
CRmYKYuvDf7Ylk2jiDlvtIpyy5sc6WUPcJafHiVPt3f4ldAvNncYIp/y6IdqpUPeQY6/9O3gJSmv
WgQqy93HxpPEPYLAO2BWJGHX+e1TI6AXrrUVtBFhqG951eCnFk5TSm7pDRY4rD7OjZBHTYmTZ4WS
kQyBKk+n/gGmEAoESCmZi97QItHOP/jQ7eC1ZKaFEvJFKsWtiq80ZSRU5vJ4ZKOI2+FzzWt7oGni
7Xq3YB9mO6okJhv3qzfudHAL7ARrD+Bw8MtVWpfWwSTi7MaTBcLDH7sRIHNITrJx0UEd/KNA1y8t
cI6Xc/2w8FU2A48kMd5zjFM4FsbPjI4ePmtmgMId2yO0egU6A6eU+u4vPq8upM3zyL8pIalvoOcZ
h+wMbiBSaXLfL9DS2sZfG81btFHYFl5YU9P0+D1lY5G1B+BzJ3LI98YiWWtcz2R7hIq7whRgP3XU
R/sWYpAy6DntwH6tQTkVLmm22LcyP15oEmiHhsZXf0xeEWH/smMGE/w7UZckAqraJgVaaQryRrKu
U1RvtkcDbpRWE/ZQo+LUC4cSpmI+rk5yLowIXwOqB00r8ANwW7kZ9cDU+Z8l7m7TyVHK8FTKp8aH
9Gnhq0cazLxEEKrm9ptwmO3Kvu6B8nsRTGl70MxHNcCbyQ17/Q4C4tjj0PpT+NKg9EaPvzK7Kc63
w8pOLdgSRFyDlXYAQybiUOo9NPFGIbPi5Pj8ayJAsDcPjFaaYFJoy1WbxTW+0FyXtiDsTZdcUoz0
RRotM679FoI/z766/Cf263rPAlTxRUrAK++TDSovYuHPdJaA+I6h8f5GRIZ7La39eTEGDGtowKSx
Vk0OKKC3qvlcHzjJPdegrDZLl/ZDYISsTWJuobUfEfc27AxxxTmw6iVM09mYOYRVkGDbFBFvoz/D
mR0kyoIvhmKYeGw68R6EVwzDyGwI1uw/4Z9u9Nh6p9r0Bm29DOE0fzUsno1zTBGY2PAUVN9M1BjE
CQR6Xw0MOGmrUk1sMCDsCP2sJaPOomcEEHq9FYBmaF8SvaCRV+sQjDLBiNruBn8ROu2uW5UL2P4Z
u2xs+/2DVFR1T6qzcAcKbbR8Aaf0kDRkDuXSpRoGSNIdBRPyMCoUAYBXMb1vql7qnOSrxBmM8IGd
JOlD+rXAFu47+ydRAaMis7CoEC2miuhIO64/yo4AkwrQ58Zv4xZhzzn6cvWqJvCwfo/5LbGJH7jo
0Wf9/GHBZeg/Vf2cRWfSaRiVsbKRQpzcLpe8jedB5dKHSF8sWEouy2rCwNpixtjuTNMdtDow+itK
nuTpxAVhPWSLz2/CQket9C8NMMquaAcKBC585Q5vLi+x7B5QVa79zNVLdWYelqUq8CjS/G8CBTrG
BCU+lUDMh46jTdy6f0s4eywQJigIN/DA8r+AuOnq55bMfB+nD/AhWAcOK/sy/74jc66D4/SMWvuT
mo2eP4Tjj5dG+eXlYtL9G+t1uAKkXSaeqVCpUjHTJ+l5RMFOVYCPAA2x/bznXHQzkQYy2CSm6bUA
FLYbGVIEDcyLDMFmw+2Lsxc/hS29GZbg4VcZHjh/EkLyxVn7o+fBtjT/X6+9Bby6VupeSnFHxots
Wj+Q3+3bVroLAtfOd9bxXlP/j5S9y64jT/x0kcH1NOuCilhEpBiDs01a3JVscC93Otz8QcrMpRfp
+N6dPfCx1fVuk1JY8oUsmx+PT+DC0gyhmeF68tb9LhLaFEW62L0QuVkWwOQxbAIstMO4ulYpcBxC
YLnug9E3ZCVzEbeTEndjo4+0DwSkZy13OLCZPgH7cXyKhjZOjJc4LDu8sZlzQfFry3b4NXUIA1gB
PH+luaWtEq6rJezHR8BcFKpeBGX5FWiVLU9jhmCOB5nYh7WB26WrZIFqDsX2QknbT05Jo46dhcas
cVE94uIiLZEjm7u8Ybem2f+PZwQFX2yb6/4bD3FyAgjfnpT4S8iKhPM/hICvzzXpPMjLaqHrNgWx
LdVlSWEJNLo2ab2rD/55tad2lvkKKeVH6bTcxuSWqJEg00OuynKpgpLKCsNGe8/XJ8F3oePty/tD
W3az8Pwj5IA+gC0Xtdtyp2Zu/u91d9K5JTMt3Gq2FLZ9oFEWDZfkc3C8mLdC1Kd2UZ+XOq35TR5S
z6yYboryYNjH4CjLcIU3mRKpLQiAAJlXXx4R84A/UMVVKFlG2eoIpSPAJQNu8eNPSAmP+BkV1fhG
I+z7kc2pmSYvizTlj93yxRBNfFQzbyL+Pp5kDdFPVr3mA0v2KDfE5yJdEwbIQJLXDvXJPKeWQCEB
emHuJCpSNy76F9IhOcru5QUaruyox2V95ahnIgP19CEnkugkkx21yCMGS6XTAA8v50RrEEfjOQ2k
e4GbOI2LpB1HkcIHzBXAjdtShf7xtq3KRP8yVREJWLnY5MMOK1XkdtmLwV6Ukim9m1X/5GK89Vv6
qT9D9oSJO6S9FTPLsaLwa9lvXs1blTU7UmCRf7/HYWAs9KnsFQT4bd3wSA8V2GquhxM9R1g6p4Dd
eYBc/6RK7xNNh5HN4E1myHCi6U5GDLlPKxKtlBey9GTZPvZPfVViwlFlqRyIJmS3bhBxaSFq6LjP
6kCJa9CzScyqKpoIGjnEpigPqZMrOUbsWNA5hw6XUJryBLdZz2VqZd9PifrBuoevL8QFAMf9UC7R
pX8KSlJgyuIKwoAOUBlwMRBsx6wE4N67lNogifhU4nAo1XSiLXroh0H5C8b9qxu1hMtZumawP9D4
hbvvZeZ44yemS8HfZ3shPRlRZQIQafHF2HEBk91EYrjU9jlPDh1jIcma9IdFQVWaVrbhppVsKzri
GP2QjUJZYq+SXc55FFqJFaa6SiF9JJIW5E7Zx4aLJnWHf2cciX0GhhAO3FwGumYcwsljC2I7m6lS
MhCLi9m/JaZTzY2zlNgh+amYSawN5w12VPpfW2eWEdWT+RnwNlTXvJ0e/Mm5OIgd7xcKk8Fcrmed
EUhPxicELQRHj1B66mKtb2DSyiS/+qcAHCciiVJ7gySlCDpSetsxFhsv5jcOn0asH2r2UEma4cqA
t97D5hy5gB707WADX4ImnIBUwwipRAuBIRVCDqpeijRgx6p5O2bHfiV9fni6PuIsXx3HU7t8dkFA
jzfaCunKa9EwmZb1vZkzEbBhfwZ50GCRaOIAl4j30lUmT/H14+w0TH1e46zutJxWGkRG0vncpdD+
HJfPgdQ6McxT9EKufvo1WVh1cRDyaMqlnHNBrK2WRYBeGrdunJi8EmXEv8WcfVatReMFHIrwAv8s
HVPn296Zdm0jRB+55keq5h0DiUP+loiiASylMGoy5QaNHu5z7DUXAhdtA6wuvxYEZLYE1wvZcKvF
Y4vECgmkHJz+UX/7Q89viaAwFwX5bxKGksFv357rcG4QyAbG6Y1xTDHSfKqiumy379OYpeT/SUrP
fXeM0xY4mZBcsz2+lm1Y3+86dEhC46ZnCNUlhGxeJEQrYNvMk6viHj+l1ESsyP0o2f6bBT6G/Q/2
oAvD/GtFBQ9mkhuKHp6h685zfz87h3ScPXfcQv1eqQn8sTYqW7RnYt2m5aLsE3BgonB8GwGcDUNt
6Fl6rB68oUbWxz+7Z8HGuh8cxHDHhsVP48ACHj9y6ie0nfFHkl0XZ5+KKC2FekNTMZzkdZL2k5KT
IeguPtsC/PnzcZCptU8PHTCxZPLAtQe97Na7oRzmbsi2WXGqecoSgGtZF+yqaouy2c9JiPJG4Qp9
RqxdRlici72cZ/Uxx2nqHHlylEJ/FXsN1W3m/4GNBuaYGpTqAhTlZcUTbcUXL77PSKnxbGPcuM3T
XIIPO3+dV6o28eD2EJhl9H+zzGkXI1MpS/o24hEwe6cbacqWfk7U3H0QY++ocwwPh2kP6CCeStAc
xBoj/bwBcXe6wGrPZvTT7JCFJexZB1vNv61RvPIB96sZYsNZhaJktLSy1RdckiBO7Iq87JuE1f8c
vzUSb+kWQ/ZvDY/zTJs9JXmUzGZ5pkme3YnAuvbUSBKGyD8QBqg5VVtL8zAPbjf2/sGSTt+r4cXJ
S98ZtOp452Dxrpkgw6BrPrH3vHzQIlq7g2V42cK4m+g0Hl11Q+tXHerMr0d+y7a6Ku+43AsQGqCp
br4UMJEnzNfBhNasGokjg0LpLk0QqOB9Oto9Ifn/EP4UK7u9G+tAglK+C6BayotJjhLcZIcQsIn9
2sqeUQbuxaVBPOQbYpwQMxhl6aFKrHAzWGfPKS9OH7GcP8bmR7LcSQHaMBtRaBmCCIgrQu3hXemZ
/u+5ILKTDjaCs1nwDf4ol4S3NAvs2Vpcguwms2zE6bB62ZNYRuDOOogMIBMEL4wrTtqK7i22HrJ4
kagkY0WPZVZigbUCx2/nAUWw8RBdG+KUc1z2xuWyWLKEa0YuXGc+qrq7Re3SKYPOHMC9s4/KtvZm
Zu1JKED7GtTl/m2aRzcuFCWK+ZOL8bK1RWBNv4O0SpMwHxow1vQkaGyyeIRE7KnzbsiktBGUW0Ex
C0xodFwKYRS05vMm6/hoZMgrz/VfxG+jdzQdkqK9IOUkRmNABcHoxi2Ch5ePLJoq2GhIr9O6hQTt
/ZsO5YPLmoGGHP7D1piq9vFBRSUxi/wbOE0Sl/AB5T7K1gZ849+gESf1yDPcohBsl87U4Q6ru/CM
R2bIpgDhZvfMhwDDyccCw/r3Vy5pcEBlSwqo7BBLi249KARcDNSVdAZXunmnaRocLKc1eHkac8WU
Rkso0gTkB9+Tmk69+Z+bSpVAZswvR4fbVHpWSe9M5NOIS+s/WqEVmdpCE5+4JeNyyQDI+M5/Nmxe
ds09XNhdr0ACZ4XykGsNPRWnsgvpN+yxoGtV0VZ160PPKPHSGZAt8RLaeQEL00W5LU1DuqVXclRq
lP0jwN7Ci5Q5Vz+kFEDo9ZthPhURNG36VDJGC4dNtPP63sGRv3cFFfSjRe1i6ka+1VZmxss/G9Q8
sMD4nh2BJbb+MnhxhdI7RsC8/jOd2oRO7xqjT2DGE22Ju5zPwxKGaJsUJVTeaH5n28JCk+orEjvP
GCOJP5lu3VKaQ8LYDzX6dQioXSfdiIcpHloQ3IKIqo4QBd7QrdoGyxvlEFRRmQgrbMUGncvfx6PS
skNKFgKGttSZ4BoZHWlFZtGw91iuxv300MCvGMnSP5uIHWNoi4R9UCRZe3yHLR81GVN70YIgJS7F
kL1cdDQEfJbQ7JfCy33hOzLdO6Qo+g9ujtHZvRP9LMzameEQ2ueXPL+kRzpiEUd5kt4QwouqDpNh
5LOcTW2xV0c3LV5mv8HpTy7gCEeVqBvVYs5wqyMqeoEmBw2Y2Q1mv6fll/GuVL6Uf6KDhQ4i4Kos
gkvmlj4I6JYTWiITqXeCTI8HKOrSfJXrI5Ag+PdcyB/rXZF6o6IBdOw1Mmtbk+YXWofnaQxYn9IN
x9WmGx3/60TMAqSkiOo1RFLfkROEH1herKW5Kr5/ncnme0GIxnDBwCqObKz0rbfPywPB5FhsdOt9
qMlyb6srKPiyx/x4PJO1oeIYk5/wvWiQBwAn5USCFwg+Ebnfrai27bWn3HhmyH5Tt8ocdpG3pAkQ
W6ttkRfN696ovo5mlQXsdIevqOX/pZY3E7pe6iHG/pRieFmDld+ntHdjf1m/sXiVGD6xgCbYjl5F
25vmN907O1JDZls19Ziq+WEEjR02GsOasFHoVEFsjK5ExoGW5QbW/nzhVT+cCSKynB9GQV8SCxsV
pJZtNomsCg7wus+uvUKgCbCV8kovzYgDqNdoJz8k5ClVm5/GLHOUJFa0fHmbkKCSjrO5ImXoe6bQ
Ro8KwqOe4pG5FlLU2iu+L7L/R7Xdfv0weUrETBkeqThwky3MKTcdnMholBAqo9kvJdfxC330Dt7J
c2/9eoO7IY7Mke+yR0TCH5GNwt61vMi60oPuNwk8/lkl7tHOLaN0GZQX3ZTDPGRWGJ+J0OWC50I1
h9kugQT+GoKJfuB+PkxIKKYppf8TagnS5OLk6dUqp7DGi/fN9n3AO4v7RVrlLZnchhyMbgiFy3Kg
SQfpQ/UqTYgdFmqKagm9wGXEPm3WM7tBPGU2Tt2KkvC4WaecfgPbZtnxZuDsNuiXiKxfvqgl7blW
NYOZ0IdR9e59rKEpO94ANEglqYMJmrEppO/qc6gXbYhoyNLBXoLnNSgUODJwKl8n0oy8itWLXC3f
z4ZBF+x6HWDefBCMriCKg0SqQX/tB9RUB2yQTPhU+QauZcil9vHghuJmcU7dOcc4Gz+iREI4y11b
cS1D0Zdsm/whiMuNaGfCg0/vO3cKmmlkSVWCaRyfa1PDLLtU4V98/EJHXb92TyoEYcENS703voKB
Hy2Xbof9o5k8nefZh2sbUk/iQ7wQi7d4ndu9AXrsmV/TqF2K1fT3Fr5mtxmUhD6orM91NeNArXKM
wmbOuC65e3fWisjaZpk8vdyP8aPkChY6S85np+cV4iSgytvaJpfXeGLXVEOH6mAx0dU1iqrbdTYV
t5ZlgBja0pdAEaMh9wAJ9HbIh219PqMbf7E5DXLmfbGUbiTKndCH0o7C5yM+VB83f7waOCXHHc+e
IgvR0NVb8KJjI+5AfWVusL9G7DAeNUiKy1s+dv97VjAOTtYFXz34EBkqHEeEYOS+sAiF7UoZb6U7
iMk0D3J+524Efrv2J5v32qeAqSb/mYS2yMr2ETzweabUogFEC78V5/YBx6J5Z1sFl+FpauaQfywI
B1NSb3JmbKQOarH0ejFWFJkxhS9WkXhkbRc/RXUfLVm83dyDVFl4x0zpHkWEZkljovX7dKLal+vb
Fg1LcLhR0EqJwbkIp/uWFdiF2X0wMGEDmfyv2wzZKUrBX8VLKITz4kS8ub1ZYorAnRD4yYYXX+ca
pxWYNQ+/I/3vHE4GfeFrR04zU14KZklahXJMSiFilRHz8fLadv7S6zbojwPwFifac8ns9IYdibwB
JLWaQW8/9bad7hF+2dOfMVXgynrZQZMcjdH91evDrXWm9LV6u21LRKg/gPnCmzZckfnT3iQ/hx7C
ww6zds1XyVYgBUVoitKM7Be/LFVnCAR+RCkBepm+OoNsCZqTj0QSLPjrpA7U8hpiG0pBIvUiewxF
biSivrDrbfdTHkAd+NGE2cXDoJc8jazw6jfbF7blR5eMO2E97UTpOAvXgMGULWTcXEzrm1p3JXG5
qVVO1Mg6vO+BbbR30mi02JH5F3+5MJNNOJhNhuSEDNlDIl8jqbhcWPeo7hMce98xx0uLnJ/9z3Hp
6fh1gX2+eXtcY3sxZDi/vg77Ncl7wl/sXdwuNSa27yjZKbXiQFQlDpBoSJkBBveL0yiD8SOXTrKG
kcA98qBlnRbcV1vTVT6GpA5qvQOkepkClH2y4zKVjOONi3lmU+1eIcxcJKqKpqNEQOXFqYFlGVHL
XD6szeCF2zrckfkEq8V7Sy7kZ4ctRVJOeFfksvDihRPAtYqO2xKBp0HndswKEmjL8WFQQYHNTPVT
eSM9syHXjGcTEg9evbOiJ6aP3SmmfBK5cxfWXDYyXRicZBi/WIehEwSFKlvNUX+vDwojgn553Raa
6XHSu5FAyJb61PCatXMvpdrpOWiayKd+N9TRNSnB/TqKY4K9aV1H2tbPb8KHLRh+fFriogllbg56
m5Q753IQQ13dANRaWBEr6jzmhTsihOU4zUxSzmh7oM62NnETcdsEvEoDcOUfGYCXyoHSraAEKr3B
geWm5KeDcHI4Gm6sJaZEKC3E72lDksBm9VsvwUGL3STgVio5OHlenF60eocLadlGCwJomRenz9ed
+z/zF9wYt6aM+jdIAa248s5JwqJ5LZAi7fE2LjEhMG5Y02k5DbtCJ/njnEZJYKBWTBIUVOgz78fg
3B3YuijRR1Msex8qk3hT6xOIm4oE+GcG3e9YoGIoaALv0JNfmaJ9Gl4lPjfqd+LO+NfKFDRGCeG4
f7lcg6As3w/RBWR0stdWlBSd3cmBE02PgqhNpa8KyYpic/oQ5yUeCm3RFan8L8BzXhdKy35QjgKI
wNCfoYXLR/XBut++Xy0J3zd64KRBNjz68c96gFowwXNKXAGw1LEIJW9gqRsntpy3sKp09yxc4o9s
K1Pz4pxdtj7tFE0SpMM7vHGrbHsEK7QvJsiTw26MZfF9LYvhZpWBrQUCNkkM9XiFKaLk0rCKZMY4
HmRZLHaAnLtbyrGGdpsg6ZZWoQnl/0CLg3+L3GhtPu7aGXwL27ul6xIBKJm/HjQMqFQt50DvKA7y
zBhovSidNPwNJlDDO7e1iOZIwSyMKYwq+LihV6z5AKwpmgrhmlWCwWzAaFuJblOy9w+XXz0Nk7hz
X6ryP7i5YaAjabVW819yj+I+SbcAB219SBDbee6svqdoCICAEhIMkhltBw8YC4sPLA1SPoI4O9Ur
+IDtXo8Sa56AeAU2f2kNHBlBSZ+o1aCNPNf6uKkwTc2/6HyntntduIa3UZOiNYZmI9yOJUUUyg/7
gFMEDpGBYMrDhU0lfjaEHFT7IEwqGUpkGPM4oe71Yl8jDTJK+PGjmZAb54O8JQfHuxR1bTShGYAX
+VqO+3jI9+ZTSraTkUa5+N4VmFtcMMoDp0JtxNtV5eV3XmurLj1FOTnL1h57GPCSybcfzIPKM+rN
YB80AM01ltwWuGqJwWi7JzF+ESxx70dq8Xyfh6PR2h1lSrXlOMAcvwCbNY5QkVXiq814lHvcvgY6
90e9PDAcjDjoNK7YYnwFgQDbDBujdNER++Bw/I1zvszyxck6O9Vktkjt1QGMnrjgEQtLLlQ8ZwpI
Ziy4RCChBON/JMARAChTpo9bqN1L1a96kN/HUVsvaLZ7Y9gHHCqHsKNOLpRmR1HE0SVfZzWMg8gT
sAmO+9CLcV49VfZGx/TeVcxH8rY9n0xfE2eIpXzbEApXtb95QdvzDYLp/ndiMxk7R/fmBZ1c3HjJ
SviuMJFACWNFhEo2P1KSRj5wS0FFy3LIWWHbM86NytIBEwuaLVctgF4dcBCbgim9pwVhncqvd5sl
afNURjTa/io44aLTcvgZHNUq7qHT8pBTJPVvIP6wGfWbcEMNqjMSXOLCO5fnh3RS8GAk0h53ieFo
Oo+Vei58Yt3X8n/G+R1ExSPLOFUlaAgi3laRR7pFLMiDOKnnatxr2YwerhqaZOSsouxe20NcCUGf
xJhW5zw0EhG+04+eZcigEppY6d6DswwYKZD1lrIloOzacOhBdYhYtxhv6gkQR3IZRdQTpSpEgUni
VXNWJWyH7JTHkPwiftp/kSA6yDspMA2mqBRm5hPYpj9nVUCDjhImCis5b5cyy7oSHxk56LTDMdRS
qTKa160mFbnX3Quudp2yLZVHSEBFCDF1ck3fDBuJkZv9BUMX7ZV5djmny2B+Csi0ywoXWmR2nGCW
m6RTObu912r+1AwcQurdGyQiSbVj/7J3/Qa6uRb6xWlD4bSROJG9NZ6Itw6yHL3v90nyk2iSrIgE
5ksf/k5CB6q4uWLrm1+icVoOh9YDdJcOASnwtjfFfNH6U95ZfpgJHpAm02itZaEK+Y6TkTw+MlHD
hUw7rVCoqUSEbW9JX6GA7OrhHwKj9QY7hzPF0FgvaSCVvGgiO5sC2pEaz5x1a9iu4CQTsWKhXWTy
12m5nrMCdEO80kHnYdulr+1CUhuq1Ptsbtv1Q9pApDokBiktU03FTyajZ6bHoF4+55SAfjs2j+Ps
yev1qg4o0/iTd7FTMD3INljTjHnOzvVcpUUqbbjSmyQvm07YmQtumvX5s4e0iputvUihod2mEuci
82YHqB+oUDtKJh/tulpq3lCLjVKIEWcsK6xt98khFe8bjY1sNvJaSoqWmALa37o+WApRVdCXGiG5
Bvvl0snDS8Nit3UKLOdbWM2MkgjAnGhfiFIIbiCWjeLzsntWtHTo0OLIT72rBxlKck/Hu6RD0RQU
sTdx1HFTPwjP5O2XmDwD/JHDVMPg9prPA17lxV6TLZ5GvlH76ePr6djzflwYLnEmLaqjnfsqC/Z5
kO5L5TjhlsCUPgMQ/FRNouxQl9Ez768b2g4Doi4la8iZ/7Bk/5oOVX6EyLzDJ38k1FawwdLj3gma
w8xiLQoioJjiQKGES2Zra5bxCLkHjsw8kiLCQ2fzw0NeBKmHcD19ynDCoQ7yMlzHgc6XB1M9s1it
oYLzaTISaYbUOqF3WiVPD1KPiUyupN/bZDE2wOSK4cM9+TDgHsGEVtvJ+JG3rfUjwr3VWoWQZxFE
x6WFd4Bjrzv0PLSUi98s8pomA7MnzkSI4OOqixCAQmiS7SZtxxRISbqWSVHhR97dajtYpg67ZuEM
7Z1CfJXxxBHiatLAdN3EZvfDkRjavqYO2n+E8mwhQf6ZG7bYN6xuodQs5a37+snNDIOnfUhZ4QEn
RV7j729Dq5AdQHhiBPR6SSbv8Ghl8mCRdi70SOTkfkoTXpOgsMbKAXoO3g9XYBd3cEf8/48L2zS+
msL7iFPHkiJtu5H51pvB1sIP0lyGItA0yrtQ2FW4DprB/osgQwhx8bxfLG9PAARgAITzTzI6et5N
yfK1Q3dHJN2N2DF991Q1CdZwY07LkmOJnqnJIOUTkVJ0PYUCWXn9L9cri2sCmTPlT2aDGvlWWXK2
tPSzY0xZhCY2JQfHMalxY6DhrndwM1TAbnmtX+6UvHx3uh4IKEgbjTjaNOjMxubg0YiBstPCkpyG
k5rc9J1Yo9C1AyCOrvhYp/RgFCZjQHT9TJGMJog1GVklFDwc8DktBW+Soi+02zuaZS1ZpoiGuN4B
55X7iqWCMKx3hcCPoaVDqR2e+tlsbyM+RCh+lQFDSxRg1ELRmwp+/NiuuCkN41d8ACQIXykQXlnK
Pqq87ae1m1Q//o8KJOd77Qu3JfDrOeP+Psqst2T0RwrsLSgInduakKvsDYsQNna24A6rCfZHLAUg
2BxZ/DYMR3n16f/5WveWWGx0ddBMLSQZhbEVZvTw7QzH9ByFvPRIKd2juu2ro7XggnSvjbjngWxv
rgnsWKiHch1rAk/ZlI3u5xilHByKvIkzc78VDBUjNZICgmu80oVy78+OYJ5HTQVHbEqndsV97oXv
4GUf7BgOwDzNxFWnXWJztBRD0MDCEfF/m5SgG5B7a0haUSxrGFR0N3JqfK1MrlUOCG0mv3x6ZwqQ
Qvd0nQwwb78oL4zdCkELOGkCX4GoSydmIc4RFOOnghSFYsnVr6ZRIsbUn1IS0n5jufwsvReURh7E
uoO5jDFgIkQobfierygg52ZEjvuv3LKtLvNghUEM+BvhbLoPbKtsqZ4Y5dQa9PSyuktwvYbeh1B8
qyBtcJADUDbIi40NTtCDWjGmrVA+Fp9BDbMCh+Xm1xAZClUK1HqUyGUs1OLN3GeXXW2beQXaQi9G
M73joXZCuh+vDMH+OtUymU8PQbr0pnNHbBDB5/OVQcMxi3UKON6kpvz5Ym8XfreDfBW78r2wJzaJ
NWMN/nmB0ElU/uuRUSExD1u3XxsIlhXz+OaepnUoaMjbw09MiyUuCxk3KC2Gfm2cPBXTzabrnSDL
Mb1bgFwXY2jErAFJXIt9Ee7hZHuShG551e8U125CuTZEtogDTRMviM27kLTVQ2TI8rEEEaogNsXl
UDyJb4w6LQf0LU9I6Fb3JY572TZGrsTvFwQLWDkvhMhME1kb2ae8+7cgS4cqAy3GaXdFmRb+Cadt
D0UqzlHepgVvsaHGitEVo59t4PK1sJEVxT6te0/c2HRbe1Nba60+I8NBBYOJU+o+Ft3Sd7LMa1lc
u35v/A3ZusOuDMiTKCnkunzBeKZsZUpF/aBtkiKhO0o/gip0ZCtuMZ8EHh1jtpIqcvcdGnvvelrc
Lo4DF0u41fBlmsNS7Y9a90lbztNzLjPf2RRpj15bDUy2JXG9d39Selh/pZawST7XTXw1v0MmPHjq
tRdEarGsZ0zFwmhcneyAabkgtXe4HvX8Nbbv75XPgTTe5blY8P1L2GMnjZsvBlzEUkMhryTYxnmi
ABiettdZQdQTUD/VkQC4GKQ/3OVGvaOXr1jKkBI6K/LCTvcpLJa1j06ibioVnGrF/GtF/ugby+0v
W/+5ceEkdrpXZyWhLcpbCk66oU2ri5+D7IvWpyMgE/yP7V1qhiw6cs1hLrkjmFdfuxsMFGVEc9kc
y1dqV/Cx2AwC1vyT6/C9ykJAKi2z16DPtmM7HpXOfT6ai8pA0TcIOC/xNNaAOahRMoKMZ7Mw0q4E
1kmS3y4Z/KfEpGgqA1zCftZgo8oQgR0VUkRHvQcIy0Uh8EDvYiDo6oCaSkGvMHB0F5hOD4oHVBWH
a/ZIlUeGApTxL8ts8rg0Fn2VXc0nWBaX8wRciIbwoutYI0zesPndEr4DrkSY0ZxMIF+x4Bhte/Ug
KqgOkSak+dKAE/X0fBjh0nSeaFwVqCPFtmxMf3c+DYCMuwaoh1hyVQTp5THizEMPDLLR61kUQFUu
/zk9E5L3jMx5qMl9SHuED3MCT0B+AYlIscy+xcVpYwbdbGjBFzVw6Ea4Rl+vPHtnf73dMrXgHTBi
xGHHoW5WovzoVFdwgBsiVpM8kWcQ2xc20yrd4dhAab880Xvy0rY+Z0bBCgea60hYdqQdx7h2HuTk
rTVl2+vikbOWQxlfwjy08fBjwN/8nh4BloWiEHp02Ea8K2YJreWCyPqN54FijD5go9BpiuwtAmhk
29wUDxqAoH6HV9vnyH9qrt79kKewvH114sTLtAjp2+YplroK5y4mySPBQ711mVCo6HnLPcAuGSxd
NM8HKj44AjIudze919ZNG2D5omsOi/oNeg8KEA+Sq44ZBLUQkxGON7vkayHfgPFLPbNfepr+Bfzr
cNdhsYRDd2+1ToW167pQRDbFB2ZHfFTcI1wiSz50u0ZQeAJpwHm5s0/eKAOlWVUKANTt+E7x/MiJ
av44JMYh9+R7zIQwLa4ilZXMJzdCrwXbKoyzg7/hnTn4qS1NO+go+GBSPe4XWqyVSwWnQ+IkShr9
7ynRlpCGBePMZix26jQL/B6K/KXPUadsI2rzcvuB6bVlJS5aRCVp57FgjEI9/g8K4FSpHW94p/Np
iKSvCCJuiSie/sCoLK+e7AoqAF8QTGwtPWhAo5xyDK9w7ujdpcTybArth4bkIQRNkyH1KI52j36D
eqFBqvjwqV7NyHiQu2v1IN3bPawiYugkI98RcUUlXl+ywHKOxKnURS5IG96jN8/deiT+aXrG7ZyC
6vWBik9h9kNniPsuUL40mpLxhZ3O1xo/QUcqtszkoQOGjG7M459maMezqt4tvkJKUdca/Iz0i7bg
QgvsJbwd/g3WOu41+DcTBwQwrF6KPFESpLEBNF8Qer9NmWpgDL0eUB06widsTC2IuVHlwPdhIN8V
5QU17m3s/bRP5ud2vxXYYgqUB31UhIs95T0dDkZBPw1fD0LB6K/Nd/942ja533/ZfmM/dbJ3S2eX
AdKzDKfApLvnqimoTe9r8VzJnC4DWxy1EgX/mlLHeV+OwvdRFPWNQ+iI+BcwkBClb24s80dcdRAC
ayrQBbIrQiNfWJirQhdHGRDvtjC5tcfeE+6mw39utCagfhCHPtciSKeof46TTrJRHDa7smNIWNPe
0yDXhf35AjfMVi2BCCMC+zcPOT9RynLH8WVwQE9gte7vlpXSg0bNvKRZ/mBOEox0ae0KiQSFWYlE
vBGqmMpGEXfONXgGmTU8HlJIMkBCc3UZhJCfuUG6Ez4BeGEnVcLq3zZ63yKo5IwdgkEoOvkq4Qrd
5pOFiH1AH3njJ+Yxjx/w6+2STk/vr2z4tiFcR1dGROKUNQJvTwuuH6hWxkuJawx0gss89LPLJeAp
+3/wwJk9y1VSIKupWYFucO+ytLaBfJ6bOy4Sx6Krafy5ZdXRDcJTG3d3qZRuIR5J93fX0UwD/lco
C+rJVOTTYDU1nYY//EsW9oyFwqrOpA6Ow6ruSowPU21oPjKthPkBikltH2H4Nba0k8DKrNTIIt3L
AGWxMSOqxC/JNnYuMH+8NJqgx9inEo9aDErfc09mKon35TdoJL8C00pQotAL3LyGy9WSY/xs/BjK
TS3eKvWsLj3MUPbaBBJyAT9N5LTbXvQs9XfPm8zfOgTEL1WmZ33I7PJSc0jnybO2qToFMxtCuQ4C
4iqHdqq/2ryQFNJv3ELOv9H/BwsuJcw+iP+uij/pKTX82OPH3FXZvfLqu5h6q7ZR/KTkdU6CcLAe
gjvcoArIKrE2+zDF1pSxMRq5RRXXt3Uczacs8+VBAlmm+sL4cLer2WQ1BF/WE1/K/X5MuAWUTL4E
ynIAD672yiB941CoI3ch2Ayqi9ZkClSH6B5v1X8XdG6noWuRvZ1KuXDeF4x3RuWG8MPvB5Yl5aSH
hv4oVgxgjPN3ht+VYel3gdopmpqsXw1YqBuZ7kDUx6Ve/W6APaBPOix05hlUW7WmHzifNm6yCNFX
1JoRHcmMy1HWZiXIurUCwkOV4K/OtOCtRXlGmEFdgBcc61mD0ozel1vNGCC1YeaL5nNcic/XXL1e
R7KjFAFnxJSGydv0gAxA08wEdTa41yMAjCMnVI5pawM8YpFB1BkGlRJmwaz+VUdy1FVceDm7NbiB
x+f2/YB/0uAB2UpikfYdZh4WGlL+nxn9+s3bzcZqPWkzYdEvlFY2gZzehHWJ+aoOJdN2oHS6MuY+
PzUf2V4gddujOjQNB1rEpGHgB1I+mkmfc5GhzUyuGBAl1yXK0N4zivLUlpVBz7y58lLJ9qs5L3yP
BpWmRSIfRw0AsL1SWBEkoYqDzJwS86J/JraolRbKfkQS3BqWqSOQRFZcSRbwVemjCJ75pmbyobfv
yeD6JpEUKRFPCCgC4N4rfTr1suAMbGdVskIMGPZSPvvoz/Ogzw3ZFutzAW8W8plxZ9LPCZ3NHum/
jmPm8p7c2vYamwmk+BFBaZJHAHIOEPt4ZQ4vR8F1rY6J5jG5VnZY6TitNyER0PhCi+TuOaGGE8YO
bS+kLDoSmLiy7+8WI+8glj/bb80IGhVrn2CLTEDx4uoFa7BbP8j8FmtJ+I5g1YGS7pTa0OoZ68Dd
qXqNuN6qwPZM96uIbaI9GGrQLJyWdWDF2a8GZ0zMwqh1CVgeszcErz7oyWl8+1m1Pc7TTaHwisv2
V/9HbnpxcXMLhViqBxGYB0L0P5DFB87kAsb4bfVIXrwc5LZw7hiAdJ/HSf5f5Q9NQi5cDWGFHHgT
oCms/TdgYRovpXhcfAo3puw/PSN7PNOVwJ/WYjntMUQZvLwm2vg5K0HqpLt8cK55bhloPCe8CxZP
K5+UfbsgkoBGPGqig+gdCUKWN6nZNvesEmMfzoiUgbGxDS9MQQm023L6WaruZqPzerYhZOsBLGgb
w5ppRXNPg274MIlmd5gy0S69BtiqM681C8BA6qvEh6YzE7/eOv8aEW/RYZ3k4go5jwEHrPQBhvBz
uyQBcjsLjKjvYtMoPy6GF0nLG/Px70EtrW1M34W6QKK3CXBaiXdl7bZSZrchHf0kntcMqimA4Bsj
DekVRco90a75zHpSglXS8z9LBftRvt0S7YFjGFrh1KA4ailv0HGV0L0onscxjmW6p56c1cQK3K9x
Z5hA44RA0kJnQeFrxbtc65J0Tw0HHviDop97QN+w2qPwpZx4Mf4LITmaddS0FhyIIEuNsOXnSrgn
XGkvQA7Ipru4Qg/8jW+ZvfAIZCrqRO3mlsq+s9EUYd+E/2YICX2YlZuzNZQ7DqwGZdFxkKwJglfm
t/iP8RArjP2rruW7rtJi9MxCBZ4ZgOMORcqGLvo4Lu7G2eh2uy1LNqQ9duh2P1dju+38TGl2cWJJ
RkohtH8ga6Mz5wJCK6vsshbe8F9NUxaIeye5ztVaZAvf1Yp25vfuRj1uKusfjkQkeL6OFyOWx3Ba
XSokD/5xcGWsV63hpHh0vKaib8+R22MjRRx1moBuB51wSnZmzomG+OTckgB5XaQOLjdSEpshtQOA
SeAXxpKlWDjmvi0tDAofYPivdYHf/Tp9hPGoXWLawnnfYpdwgMBucJ624V2ZMJbZVyEZG5XjcpfS
WC/xjRx2dlu2PnIfGwC/P4U6yi1chdYET7hOEXQhbPcyXWTfr1sR6WVXLjdbeDpvFo4DoPFVelzq
QnGQ9uy8ruNiYMVM6VTCy5G9GmroL4vDbeeTqCqo1JpfItAdxA8smd8He0s473AGs3ECz0BRlR4b
Xsd3vJ9uOYmw2uFewa4/L4nECpKjWtfXt5eLiQj0ry0gHDPULysu66mouW/9G6+plXk1YTmQ+uUX
FMXd8KW9R0UVF3wDTU3INDjL36x/0cWPbaw0DPxvKwzAA1cA4DlYGjF9hNKVpZGDl+ZhAhtusGqZ
ZSTUfM/oIuck9yEAXtFL3xdA7KeY+r7HDoPGjtW8XSKg0lpOvE+W50RhUlC0M4bQMPwdnAwtb4vR
85FcmqLPAHSSbGQcmqRNofdOykH1rMn3dSUQxrhkmHaOwGpOlQLsiA5ByyAsns3hpH6ebPmG4szk
5JVjT9n7u4v+SJyJKvHSX1xEkC5EmatacOUUEWxqCIjyjAr0HP2dba3yHd4u3jn583yb54Wr/+pJ
wKJ6+JhgfvkpIrL6zUx7nubhJPA0Bu9syorOKSmEEtlKVRNAyIa49E6ppxbyUQPIw9Wk0FyJsyup
MykB79ET7EbiKrM5Wvf8YeQyK/wAd5MsbYEqN5IqLY2F6suAwleqvQosEIG/TXiugyVlAAj288zn
234efv/WMqw5VNlNwD/I5T74OghxSS1qB1k7v7GQ8B8xubTuUCfzt4JSevloMAJACzu+YntkCIIU
XShTrqKUt134HJE3H9lxDGb+NDYvAjhBdJ5PCtSUTocV+IKS96TmdePVYqmEy26hD3d/OkILYUdP
RAaUvEOuRIblmjEg1zWvUOdVSVtkEPuTD9+7Fvfk+Dm1HzJN2agOCyEz5LCORzt0BKs7OEdWPxZy
prE9ytoItypQxDuR0i2+ADeTisZjs98eiHG0kwiS/Xsbh7Erm53X2EhUTwF3j2wIx96+4Fp+eu7H
/duklT1257rFiOUubp7Kr0YToRqbQYmFhtsGTqYHGFVPAb0DDVahBZllga62kP8/rhcA5anaX9Fg
VFTpJOK1H11EGxFJiJacELqyyDsP5NxGdzvMZ9YstZdFTQjwwDDWMXb9Y+zpWhRy8gLLsURX5vsW
YURNDga3SfRki4XgwERFCHzCs41jRt90C2kWRuP/tcIBFvPH9R3rdtcXPbf/9ZTJdzFFBc2/e0cS
Qkv5zOU7Oj4g8NIpKPrDuHHLMdimAozGIbET9kDut+QWlDk0jTZbXdCjQoxL9vU01srtVBRlSnNj
Wo+fQoLMxPEylkrUHKcGCAz4oPNaLz6xIUg9ooPvnaT0waxhii05cocvnA1a+mkA7zJEuU0tI5Kg
HgURfDAP81yVdmjxs+7bMFhthHpS87X+bHyRA0Dx3l5heDvuvALMEZ3t70GOexpCBUUFT/Pz0jF0
6Xt+Hji+fIXuSY+HQItxLfEnBhoaLJeF0Aw0zlgQqrF4GBVbSCsjS1jg6hMRz+JVzK64Apt5wSW/
KSFcZXLxrFXxEGAFGPGVDBbfKZnXnjpIMgYdB4HuVDxFI/tTV9GSE+jo+/mgmllGIL0Kfwy9c8ez
fDxivS/3eKdt0cLuH8zLXz7GxCnJtPHfu249FWSBPhznGgIPlTk9vWsv9MywxOA0YITv2Crn8+UP
CSnZIpu0zRkbKB3kOqxMxgsI0z+YRMUeJWeSKrl2wJrrZU2Uz2zAnZBDO8wdpPafbxhXAlYvVKlr
2JsOsKaHiILlBsiBQ/RrVqRK+SoFPMHiPihezImHU8WRa1Hz/Uf2I678EbXNz0n0aCymrlvu938g
o+OTMxVyEhqqgY/b220rX+DZ5c4nDjMa4znFEIG0DC+uRwTq3e8BjH1hfzk7bhXiT/nBwHZH46Cy
qdpyg6rLZg5DYefMEjZI4hjvrx63LkmfhOioSZ2adbwaTkRDvN1f6zgJisEcCfcRApZetA/eftHv
Bi6UHtqeTwThRKDU8pOX/XmNBL5lhG4NZpGVV8eQBZestd6Y/fOyy4YNIsxtXkIQQFLMNRlkVq4N
r6hIzNkmyGRw0/PzTB3r4KZByeOxy3E9eXjxi3yKyHEg0sB3l1W+9aWm2GpfySatZe5aPUKT2K9H
YHblupYNi/Wj3Tgx6deky+V48iwqT2JKXJM4Q4IU/SKIwvrwkh+crtGRqE15oyyctMZtE/l86PC7
yPBuNWUCA5t2zkoVSpA4AbZdpV7F81/U88QsRiRfFaEY1gAzzAtyd8RxwZkTzKqk5eU5sBduvF43
nl18DcvF+uhC/GZ5wS0IdDOBpq4X04jnMpN4KHow5hz/OXjaiFRc+cnvTY8N94zmmq/jzDkk1GRY
9om0wLRHcDTkbYhGGTi7PeW6qfo5L+4dhxXEyIVIZqR37K0Uyq2p5hd/BPOpHdJbtzKhskRbVGhk
rEqcUU+zbihZ7x077eUssJg7qhNSHf0tUMQ1RmVwnr1HVmLlT0HEDEQHQPjAK0E6vPF4G+vwXeys
BGis5UhiB1/IyFggzHcRJrOkU8eIJMckGoxkYripo48oSKEp7DohnAshAv+SpBcUd/+PEbxGh9vx
v61uy6zAUrSyN+or9S0SCmELuFzcJyBpaT2UIW9TPJvHu+H8ccf8v/Vw3v/qjgSTlLZ11m9QH9eg
xAGGcB+QRvIBMnwHYCovvL/1xw0OdgX4cTJl9cSDgcMRCyOFm7xjtnoIpFd3jfzNzWvMvGuRn2Cf
+w4M5I+I4Eu6t8GcqwyXDkdJ/aJvHNQa+fZeJPEdJL7SUtbyyByRKDZNfNtRMS8Xnpg0qckv5OWs
+M4bDFY+A21PeVTs5nvdJFlHCESwBCC6hSB89kKy6FsdthDQ0KlFya+7DdRNQbpZ0rKgy4rQBQVj
iH1eQYD8cPjB1Um4ah3ZPI6My9eXRuY3m3BFBcKBMM5LeIMV1hyJk1epkmWQ7dsRILdelRU4+2Tg
esvLVAebL2vDLgFMX14rZaiWN1D2vd/QPlQDXTxMoQmhglMbmKmhuxnjwQ5vH0VSBqR/Xe4D9wSX
/U+mTvYR+9in9M9mZ4coaVacaNkOE0kPwi/OPHPLZz8fRoWeLz2bchScDuTKDrIQcBxNWI3FVgua
H6N/9DCg8mw8nROdvPD7hIovXucKdRly5hkq0SQBjsC44Muy+qDqndpRToVrGyXHoCQGu7DxD9O8
Rnihzd1Bf32nJX/sH76Rfq34QZ6F1+wDwkyo9TVbpqbyJRIgUPd2+0xVHsSZIeYhzF8eRyI1LG81
ZyCAk6GIxh29rNlw6e6qAiNAeK7lXliIZ6qFb9cNjXCx4sa3vMcMK8OiCtfXjVAzjcV90V6P5Msr
WN+xGzCVIx0huMAJpt4e09tRMic9MXbv5aE8F03d3L5XayLcfXqUOtclm2fnp8i2CuJcolnBAyD+
uB51uSxae3RP5uI8KLawooEhAJUFrUeVrcHh6Cg2h4a22OnRm80iugDwiHraXglfgjllByZmDlPW
nyjuRIEzpapTXMQ5wB0psnzPzyeIc/x83ce6P8IvvZNiNAoqwlbClVy74XuAtOLW3P5L4QSPgbVr
eq6eKZmOblnj1rFhahGU56iTErLdfmrBUQP2xLpv7XQSBFfFkGfBrn98GnzO4pbfYOHFjZYMsQFa
U1YvJ8AqmCZc5VvmUTPDVIHWsjW81mTrM2DmzrP8uGAj3R/CZ99ZQYO1Zbb1oLrB99smfLGaVBpa
jWh9ROH6OnjRo/VWGpvESGHcSXAzg/xcZNNTgx3LCb5coM1KG6XqA5s8dnZn1Cxeu62xAXt0iaUl
z7I/Rl6p8xGuU+mPBSwFdl4+j7smAMEYXaw2mitN4LQuu91XUbVX7mvn7ntWXIg8iIep8wBVu1nl
hirraP0HENktzRY1qUUKctOXeAqatGu3x3NzHhRlQrxPojaGWIjcRqSHyWLbANAIlLT4ch4NwurX
H7DNWPHvgCTdAKHmyI+EfGPEU+gSuvQ6pTeigIT+HGmYXKojRaAZkiVcH9KWtedC7SU/90rxq4S/
hZ0AW8fR8eDHvWIeka/EFCSjYmDqkA+H/Tvq++Q6IMut4RQUJg0KX/sBmiuWRp5IXwGA8qE+RqcA
YRk/FGW0a5k6RXAdw7hW4LIbJhoVX+2If8wOud07uBWkeoQsNJD1kD7/X5oPLVVMv5uvmLFN+jG5
TBGmelHJjcHDgln+2AFoFJR0WU7itUGsfQbKFETbGVUmYa/QHNjA1k4pPJIU8Lf87+nA9jOMVrjQ
YenhmOdEFUSzagEu7F7lC3Ow/yetL5c72TNODxRyr3OLlDN864+ASDhvCvVP/yC9izgM6yRPmGTK
mDSRaLJwgmjOnppEL6BMzYlFYh5iI7M21y9Fp/KbTCJwCLrPmZTBLF7JQjrhyJcrXM5exMrjEieD
eqHdSWh14MqgmVEcOx/IY/wEXKOWoHu3lg4bELVQuv3jmjsXvWuBcY+Ej4vhvAwNmk4mLIeClRRl
+0noH/W6TaIKbSR31/ktVP0WzWYuiMU9QdVXHO3EU3bq+eE7I/i6GxHoM92mbOaEOk+l1Pq0L44y
NSBJommoX0cO+S+gBGgemsPBqHP2cMLjmR+OxpDkdlVNqXyVUGXYRikfa7sBtyLG34hMcDs9PTOj
sBJlgLoIB8y7z/o+ZVwszBoo+QCJT9YLnszAX9Scii9L4+b2s08fYuqy+hIZeR/JNY4KOJUdm3wV
aOJMJNx/nzAN3su64AvPrBDPle4zQ+OfaHGQ8snM5KLchCz9MiqxbAvTu4kgdE+bHl1efwf40m8g
wYIlUJwS3pj2in8JwFGk6vUBoWFPTRYO0dRAqsRvN5TzdGgdpdVw9a57TA3aDuM7NBhhAqVCLDI7
zucqr7TdsuF8LXid4R9H3kYU7xV2qQUk2gt5uaZnLRn5DL/Xpgd2wSXAtGqYTzQuWiqAtuGWVan6
zXII+y+CIv0H5lkeCTBxprorCPa9lHgeNJukJLKLGiO8U6qR5qB75/I/WJx/T8ZP4mTXsaYx9I/Q
w73ynTe7ClMcKOKwUsVwzdHWN8l6Yoppi3IignPEo+TXxwOIK2AvJkzQ/KZjQsIhBY/yeQq+vumU
xvj2KJTrRZnki2gT24cKGn+TkdnFQNAOVxcaQq2s1OVX37E/TOzm0cCE7xiljcFhUEBt7+8aGsq3
yZuKFJYxGtUo2lJanRqB/VlsYxcLS50HT/r9Qn7291ZgYaYxML4hmyYbgkVn8OGkmK5/Hkbskil0
OpCD0C578vNfCRLT+p5hGmwrn1DN5X1hEQfpoeSd7NbEfyHGBrY0/8K9eiDAmgeQ/mdOich/eLPV
IcoczNUch9NmiByhkZDbwztMjjk34RlUXBwQcFkrO/a/j0nfQZO/TeThf2qKhdJGCPistxMPCzWi
+/TwSF2r693hW7PyiqTtIHqsUamHlWp48WvWfca6+OViTDUicNAkvPom3EFRU/ZmrmLPK9/bpu4C
+vh7oV/xVqItnlmmSrsHaw2QHZqs6v7twFrQrzUnrK8FK8n+c0fkdGLkCg/+cxiITxjYB9nXm2xb
DyJDCfXKc/HW05tF4aDRBmbFtQuEqq6G/+hNT3u1PQQtHrltpn+t6BnaPYdVvBVq7ptTdYf5+DFh
r+3t0EAT9ICSbAGNZi9OyvUYqr9OdyUDc2TPt3PCgQATJaB1U/cMgEzPXalWSncFZEMI60XlW6ge
//rpJD5DgPDgSFCKVyTQUls+xK1rCUM9/oD99cb+meKcAtx8ugV8IOQjqG0x3xJqawcijgyvCNZC
9glknCxz4RCUXI631dIQvx4FejFe6zYiwPvxCM4LLz2qrSHtQ6Bo9kYnZiHJAyjnMSI9KrK04yHt
laNZCKBYLbUcWfrMjkoT5VzbBmTpZ9WF0werCW6CeoyzerTzUX9k7nNGC3mpARKpc3rGdUs3FXKg
qf8r1TdYlB66oVsGRqcLxG1mJGUsYNaRVfzwhqxzLqzXcNWYtZSsgVtp9IHPOR0kLspnHSjczdcU
gJXUl0JHIPhHwFCrt/iRXfhPU5vLoUAMlxTbg2bxbQYDO+6y4VRphppaogLnkD7iw60jhrmzdRQf
AKDpXycSG1ac6Au1SmL271fmRvUCDBW4YCN3O2ib08gCSwbO5NavroHcjrTybkZ0eNbV5trvLz3p
js74cYaGRLiY4j2jkyxZ7ktP5tTPGdIgLxnfBzxl2Pq0RCD8OinjhK/DisXgpBFAYANPmP8HXbmA
oTQGW0K2+UWqDmOtr6G1SjNW7hCF5hjqxOPhW9aFveyCNVNSEvoObCDjuQhpa+5Ks1pCpSfXDubw
8y+/Bq+u+cZSMHN2gjSlNFth0lMLUP5CneReKi16CM9PTIsQ6CeKvUjDoP5uXRj1pE4ItCT6As3X
ui7fFQ5Ab1OaVP2qR3PAlPKwz6ZShYQdEKqMb4hUCwUNA30GWYXppu5oG6v+bXmfkGnnaMxn9hCc
R3DTar+EfJGtnl8RcisWOsPeu1i40GSw1MIUqjISUqSVebkWxnbCRNKJjyff2yXl7OQWA9OS8W/w
vqVWnBl3tVcWg5BckLrn7IY0rwY0KzkaK99exDbg2Zj+altG8yBHabIgwVq8GTz1ua1QFc8jeXq8
GQ8vgOZjP78n/M0gddgi0uG+yyyHvrva0YS5aXbeXjWgjuPqhHi66xLoYgkegXC6EHhXHHWNfij4
zgUdlvgn0vU75Hx360eDg4saCP6nqKfipJJ32OvwE4aSXmTJz8utflxboZ/e22GkNxH2ton6sFk+
DRPsdYR3EIivDomSJjtUc33mLy5+cu13vI5IkYaBWc4W/9ubta093P6kGglHrrgKZcFQ2rOkO6pr
871AH6jXvhIOHTvjnuD2lgt+zjsqVkh5ERvqLj5nXFKWQAaz3yxTSiut5ZObCrkrXjGjkcw+bqfm
nUM1mppLY/YRReW155NP9JFQZU5lDhYz0mMmwPdT1toMNNYAN4BqA9REVI93c8r8FrmAOeb+g6/L
p4rOLKx1NgCVumZZVKMERvpvQKVcWgnsEaFHd8YeYUha46vc9gg5e8qa+cG5F7Yr1ajRybKwSDrr
Gh3jSs1AfNrtoR77OBQkbBAhoPKkXwnIHCe2xreBDKUxa49N1ByfAVzqqGMy0rQ652Pm8c/Z27GQ
4iALizbzHDJZSWlDqqfDU3pff5ja7XmmmwIVWHq0DGFsId1nU8eAgx5QLl+QAt2yWZuoE3YxlVl0
XdApOrWdtuOpPtHUa1Sv9TxWD7sFrQevaKklOY9DGJp/6ZKj6XrbJ0MhREU3JLjj+/5TnUrr4Ww6
xghkyE8oy1zXtVTvwGxA1+zeN/kaETJCAHRlln4ezjiNMFRd3LhkwhbR167PhJRNOtGVN2bcOYjL
NT0uvvXhSkQxm+/5zyeTfauImiiMxkV9jGLNT3KYWGN7YYiMszMBLYEtFuRVJazbICA50fRTUDQ4
67NkBvOe/CSSn+bzYl5ux0eAFppuv/sYr5FLjad6Oy+MX2e3jUcVVTvJgeM0bI7MfI3jwKSvngM2
bg5K6niI4F+WkroM54v+aFH0LAACMjqolO7lbkdzW/57yZxuay5nzwpTuf52OVmPboAaDRlsHHJv
Xa2L+uJzqwvBvrB+6VXc5q/lFHFBJYBPGAHwJOC7k0XIW2h8P3T+LAQYyhcazq4K58RNvMVGIVDh
t8BpTs5g6ING6IUAS3hG0wQw+HMlco2RveUy6gPFlP4d/Bdt5E5WO3kj1sVCU8PH0WQXbqNYv7g6
dbFGR8R4HqWe5GyH6goQAsFTrie8N1Cm8QJGwK64Jq/WdR78Kjbr3LsRfBHBXBXUYorv9IUb+dXA
V9NmZzTjBf0DBXVCPahnGGNeTxPIuRF//yRg6kgZB7vsBv7EimAGnV/1EG+6rEhvmB8239lgt2jE
p5Q4qLVde5c4oqdY1wOKNlSYJBQYemVNxGSRP2yxwMVy9/h35cWFWpnTtK4B5P+WPuIaNMZTgQCI
Lc0IBHHxKe+hGoKhQU5Ysbx7h/U9v32w7OfUaF/82FXpqbCw/ZMQ2fy/J8IuutBWGuVIH3OeCID4
nitkxzchDVwzzXIMaJbGtMFm+l/EOnL0lr//hnLkzF91bs8veW3c8r4CfMhoKFayXjIbPZ4JVEPb
xWXJJg8m+WhygqYAxtJKm692XPK4h/+7zcfDTo1c017l8XRWE8lcf26wlBThp6vTfZBduT6RY07O
gU+U2/AIuBkzuPIN1eipyMhgMfxqLduiVArouRvtHbfv34iWbU8hRbRTuIE5rgoWK6GKBl9LHWx5
7yr74AraW1tGKwnnRYJ37Iuc6AxhypDfZXjD8oydDSMeTYyUsD/D8O91+xoQWsF+V3MPI3p4XtGB
fr4wzm56lDf55N9ES8/cqJHSLlFz+Qt+0qDht1A2BMTUlF1kUNWKZCtghOj2n99751JFl/XcWU0E
cLxhesUD29Hfn8kTs2ghiHCsTvh7zoEBw1GnWa9wEEpm5z1FMK88b8jJoD9FCqqqbIJuRan5apHE
Pr2bMYvp74tCLbWhOMLWJxytFUl8xSIJCgA+6Hye54zrGU5l41YnTw/3TqT/7Sk6xh9iE1S3TQEL
/ED2pDTmM/O80wXtcaeU8ESAUAoxcLgrdmlsjHB/2+MJM7yRGbeXVoIynZ5ubMb0c+LdO+uq5T8d
BfkSBk8bhnuxZMw8VAePb8A6tpBua+yzL3sKUJm/qsiZBmA7JmN7bBVszSpqp0thl16c9GRFyAvb
u6VJDRLiCXTMTADS1NAXWL4YSC6IbTn5r7RnUQH7hF94oMzlShzu9AISFUJRz5CyijQpfwyT2uTG
Jyj3ROwzI0zO3Yh3DZpI3BEgy2ZihjHQsMVqBMr6hqByem3zULRAGF/6Oxb9a20tExyoIkzV5A2A
lMPiv+o0TsAidt1iNu0CsNVOrLDKqLAu0CC0Jav2RJKlW4GasRD83/pZkqOfdpy6uAEtHXJbBB8a
3+vOQfQ0GZT09HDmkAKr87OvQ8pVf+aLnMhpZffcO3IvdpsoBGAuHWNzRpLAtBooUJ2btYOEg3Yw
5Y58LqU+8Z80JhZjhxi+zZ6LWZgCnk+eNIRy1WSztrh6zvBgyugCWLaYhZCf9Ty1QqxSo92m5WPM
XwOpiaiJclsIkbpM5y7bMo65CNp6oxKoBMbvEkcyIM/96bdgMEbiUg7ONfrR1om9fq2UYZHC7QbN
YJk4FFguA+X2vN4tBsaz6KMAXwczJ0l0YRDnfAMbjqxzggNjMkuFYoa6bNnLgWbgg9BKW4TJCaZW
Osm197dKbNVHNsd6Uo5/f2YKu74uuyG7l1OZiFkLuUBaE6N+Fy9ucju4ipRH68DiCzx3EqCnL/Yq
+frUdyV+C8LIzKfD8xXjiPf84E9wkx4DPumAyqQcxjnYegu+XrJcnO8xBiCvdAXT73oi6mqaFYMp
sRcAyl79puRVp4BmV3Ni725ELS+gfXobywxpMVWVOfmP+l92gycGYRgtUyPdb/eITBKgdMsF+WmR
DiPut4evDcUiPtDvIA+BB40BYBVyFrGVwoLL0labnNuzcN7jQGlyBnoQ97w4XJJ2CL2/hQCv3gsM
hcO9/es+8ZKC3eoozXNs7GEqUAN429sICMdy9+yW4jwgTsZJfpTMJCiVc2z3fyVu5f8G25kkMjFg
Tn7BY/40nzTFmqrv2Gck3c2vphU6P4VSD7fHbk2WZ3pP7rTzuHrjWHR0RPGHDFmPqPDdochFUiZI
pjmufa3N3QqriqZo0ecXvDtRIXwkUeo2BzFvo6j5sMxMpo75XVVPkHJTsXlaOgLtl6fknfAIFA79
tS0Mm8gVw9rLC4WEuP6lL5w/0CCIOvZxBk3iAS2tOSmc+166+lQddT9PcB5i1t9TI81m8sNRpAG7
dLlTgW9ZzLGSyhXmBZF63QdXw+Bf4EFdsttHPCE70uteje0P9PMFS6MwqKcJbUOSokPD7NX8uqXU
lXCJ0EPfjbPPNGq9eFeCTxCvyBjkD6oC7Se19Y8YTCWBnqb3DQ5yOH99OtB29qmLozKEg/Kwz91d
nqQuJs1ioqnn4cUCuY0R5YIa1x1JaiqrQXhGmqwrDbBlSJe9qB4aaCwG3AhKbJqB9tGJDNGSNmuA
U+96tPg/Ah7BxaaYJHUdWMNRLASGa5sRH5JmlwxSq9gmAyrKEJWJOZjl6FrxlHBTVouzxSIy5uD2
w1PqeEsdKdGevTGLzl8laXrlkvM5Wj3k6CpGib/L6ngPw3E/nfF0rAm/ehDPqhZrLDpB5H1wr8y3
cb1+EU0Ym5ICd3Pj2nlgHaZ1/IRddkG1eii27yK7UbDqRgoRmjpUk/kh6NHlKZndXJMRXCPkB19G
g4K1FsFZGEtwU99cno7zPfKxLpLKFlBl/s6Ha3rUCDwqyy2jaoOioaXzEoh/dWGWfQJukQWmPHkZ
oIBA2gOxmMrz3Zks9xqFbtI15lLSinizSRpFk3ii+89sth7oVkZIWfjGNQGmBt+o1gGW72u71KLE
zb0+ExAZJvB9NY36tGuITZn2WgwS/yWuJCMU23ggYxSI6cjMtoufXzSxHGW4Vetjr9izVUZnk318
0RCxlpLOQc7478zFW0Wcy2TizOUoTuvH5p06UK7U874rGEEsx8X1csOF+Vo3bTo/Jaz5tLcN47rB
IYeMtfG1x6F7VJDdfxZOmMPQvyvaAXegFOz0nE9lGefp3+ePq+o05/AY/IV9yetj2kjIzvFzeJAk
8XSP55OQuud8rdnQ4rWiQLz+CeeITvv4trrp4G8akq/PW/IO6625KAVSalOoY9EO3p7Zdrk9vMB+
G5l3UE6wUvS3Bn4ZlqMJno5CTax2JuQqeyjKNeR5TEermXhIimZukGN8oFu+tSVPtdVutiOSYzB3
WMNNcZajXBJNloB+6qLTue2g/fjukw2VHuHVwKKMyZ3XcBVVwO/fA/j99HCiF/ZZ78fTZpfB9C14
IHWX1Bt7vTFv3g2eU46xwFoEchm2ijpvKhW36pmXGHBUB+MjcX3zi+J0vYuTd7A1SIWvSdPv2jpS
rJp+lXfd6nIP+bberwsMSkcPNtgjNGujfgSNL9nqDVU58FgerqvIs45GHZG97vlZ+gQS6rF4rDvn
P5pRzhHyzGHpLfSt5UOtDnRWmCyDLRd4vmoz7A/KdYJCTGJdicAqV0v/tPH7w06djAz/yKBz2FGw
+4oKJ9mCp7/IMJHvvZT4lz3wl0fR7NNfOUaqVwYh8dx59iNA8kGAKrBuaJmSLnysZcE4V3NrHrLr
PA09mvTFeMzr1Z7dafRyt3NsrsilFtaMJzDnzFP63knh6Xc+6yRkoKc+YJJMYq3lWVL6B4y7M7a7
o9cjVOFBeum3CvMrMnKn4BhEFhXOEz0jOPHuPzIf102ns9gAwf3SnSx5y9uoA98b7MZslAYy8TtK
TFnk8F2qPVxERZ4QycLywnEMOOoIjhvq2zOHnCMYYqXlkRB0/Nx23E/pN3PBPvuF3+8NzMjQdUik
i2esdAXG/ssLiDQWySGidVRhaHdJNn/ATCETZaYscdQlbObND3j6+o329wBM3E7JvbpZGKLqTtMh
UORZixmNRLZZSjjmf7pGkt1oVr9CvMCrc9VvmeX+eaM1oVuM8gp/sHUwf9X4vzemtXvz8cd4JCRA
frM7wVnBB+LEfqeYb3hKRsWkXTupBRx8ytytKQL/XTwxiba8cJBIOlSwDnnhL42P90NI2L2gnIyc
QPrjxxU7FZJ/cGCYlUJcvTP9Vtf3rOp5imSSsQO7OH4nHxdBiHAaqVFV+ZQhpQhfBsH4iG1iRMuL
2fXIV0BAdzgJ//ntbgLrsSKJ5CxM0tJ431kqWIKD1+AwNIoFdElPUlsKPqffo5ZtGu8WIB6c+77y
B1FEazxKqDs3i8frQGp954c+wiO4HZoUDFNaUITPYyC/73HvK2siqcp15ltJBj+fqV9uP8NDDk88
jPgv0t9PffvPUh8aLiCuDNv6kqyoj6x+fzsOtc8TdK33G7MyLiFpYoLaqp1pllK/+dk3KOVfUBBB
1V1npaDAUgZrjIT9lvDNyUJWYJ92j9MZqJMJnkZDUWykfKqNYLyW1MCG0AKm6N4AMllPKKhoHw5m
KZFteUJw6CTBwOpeZHfA1qcrU+rJbPbtliGO0xVGmbc72XjcinVN+IJMmtKD7/WNS19K7TxlZ/1M
S6D/drFVAXzqGC/ytE4MKk1cbg7y+IA12mG1cVRUd1czKlZ1LiGTnvCZhHyl/dm8nDKNedT29x6m
cJu/wXwPOlhM+5/BtFhvoqTlEP/r3qFjPqBaIxknSkLq7RPQTw/J2uh+ShTEfSupNADSTJXIt2sp
nOPV/H6fj5kU/Ir4eoAB0wQFYf9zbDLiGN84ePAXZTNpnJpcMnTERl7adjzQOvwn3YPPvWe4h6I7
RAE+AOBcSkbpIHXQanmRMc2LaLereTp7TX9npFHNhHuOJ1qWl2tWTwTT1H/de6JzlVgCrlIu4DdV
M2wBi0Ob9yJE2xk0VGAUjanxLRqGSSswg0JZhPOswoY4WHsXH+nnUPOmrjdWISbJxOifsVyWIyu1
pIfB/Y3eolq27Qp+UYzKX1rLBTqVeumRfN6n1IlNtuQSJVBg6hTNJQChmXgPRL/bKA75vhx0imP5
+M/nBlhikXKPL1C85+sua981PLfdhI2lOXaLaNe5Y6RsSkdRUw8YMlYEw1mKpidwhFcTt9pvsFHV
t6Y3z58CKPjUnWc+Bvi8bnlpgpezgz0hJWrznoeF2QTqPN/HjoM01bYRMB36b+e2EKa2s57H07Xp
m/nXLwZcLPomD9Qhm9iQjS24gTa8PZlvdv9TBibLk9TT1xd2j6tZBMxFbBGJtrAEVT5EIEGPF4W2
gxpNTDpxQtlGic7kg3gHnfiXIV3cgfQm6fQmSt4z2kyCsK0VzjJ2hxOr7399MLKPWZw4G1AZzYEd
JGu1w+FIZ8mRBhGIcUc1gGzWx30C4bBM7kKNZzo9CyqkHed0Kzk5zZL6i4YimNERq1f3EkjAsp9M
dW4w93l/z9RJJoHuD1RS9xceq+ymtJA8252SPygHG6WtPEyRspM3Z0+B8WJEN+FCroiO3yhIo02m
mVQZNL78MRSqcRHHx8ZPqPoUVr5yMSlyCjz2VCIJPk5hNFqTTPTOcooZhI0AQUO8DsnjPK+imSpe
RZgJRaC3ZICVp4BJQWwsndllfyXY/e5RU7V0ZYSIuT3uZUN0Zl8/FoMmsfAkKOHn7eqYx5rMHhQB
ozKP/b0cATW0pS7UGO7wklWThd56UkCyfIT+BL2rwGP8Zuv5HA/HLU+zntuZlOXnHt2N0pM/FH9N
CZolGa2umu3JdqOkh0f/EqrtlHS+yRgpxcX9uBVjhMG1JmdA/SfIK7fUZu5JztAuB1jE4HjGH5wr
1iL4G5u1NWis7FZabfF1LsoObz4+3MwlbntebDPp9QGE1AyrJ5hZnd0ClUsCHWU3eEFaJieTaR3r
RR7fkYhOpUiBDLA6FQNZYl/CMy5TAr/shVBqVvC8KVEEmhcCp7nUX6LIoE4hysXaQ45Kt2ynpgRu
rGMCiNTzxtInZKiyxl0y82rOfvFCXuksvpeFosehRIzrK73j7YHbCoIlsWF42xd2tfseg/PS/d/L
xCZLj37W5G/WbFqMgpn2VVNftndJ5xRC9Rogb36zA/lOtYoE5OfRzowUYVYxIE61sBCCIkAv6r4o
4jx1ykHArqnrvsvE+tdgjiviweoi6VVjSuCe7KDI11bRZ0soTnYJjfJUS9AmmCNu2FviyJ8UOlgb
FTJ27TTK5xAjmW8d8KbhJ53TcwwPxbS7Nx4CVouuOmKP/Y7/LGbZLSZVtvVPiooqr4AUiRXLJFsQ
X5FmD+j4QTazf9XJ62oa+bd6SBRC2HjkYgZlOcRITIeaH+byRP3uOtMJDbrhI/A65tNtdohe2TUL
Q5urvJ6ORuUKCHA63kXSj77Cwb92gfD/TfQDa/sY+lHxkcmcYBcdTKQFMqv4iGDZE5pJ8RtJdZkU
tgS0jiHBI4ybXx1dFY0wpXbHJg51OJb2RYB3geV0+hIubJs9SJfADM26bPYRYw0ClREHm3r3D19Y
7ittkeZs5LTrcgG/8HgKHHjSdmPM4qpAnpzah59bI5ZUPejhbyrFitPR15EALciipOmCJPSmokoF
xJbUYLR9xdcyZFErAdAcVWNNWdO5zCnQ1XQMX+V7wA3G0CXPU1m2kltDUI4RHf0MF4TXPHOFDWMi
r5NpngGIQE9RtxBBWjqUMMzDE3AAHiCkQYsFbLoedap9jHgRlxjnR+8OCwlYy2FMGu6+SUMZd6JJ
TJiGiA/42v+xF/yTBrF1XHVknxS7gReqt0Sz2Jo/3kdqp6kogU3Gd6dah9vVwPmP0dxZXH6Jq0O3
vQl7TwUE9dM5Kx6Y5Q2LNhoMH2AJI7rgEODLD+WRPAIXs/zjcIqXC6rUykTpapwdONceoupH1+u5
d4rlcCqbguNLsr3jXoJ5FHofpSMwjezN+66BSgTd7hlsNj/sbs9RT0u1CW4VlG2ciOkeUKRKJ5th
u3pFe+JByEi9gn9LR8f/NOfQqblv5rQK7bv3nWkykVto1sbRsn0ySYEgL6vw4EzWp2h8UbrSPJWE
V/LonDFft0oDUz0J/si/XLwZ3bmSIYgS384TZ5/oTJsapvf7f3slsB7TipO7nKPapt8RYFXLtB62
dTOErg0WVC7xK4jHwsuEx8Zq2eZH5OCQwVC6+D5B89XNZVs/f3JDfHBCWOl+EeiKN/jazn2ZTLNU
7pdM2vwuuH7Uqqc/FBBAZoIryVY3qLj/dxCn1q/Ao+MZGYTjr5BW+Fnh8E+qNvpXmvT/F9C/YwEr
XWY+pDTrIZ8OexifMxWT9hiqq/UPLm3Jug0aixs/oIPFAaUU6MLvelFzhgy/VU4tefLfXD1FziDq
vtDHCqIvxOuGQZk7VrZgKlTAz2i+B60zAkk+36u03QHl9RFgFg6h7JL1GdKm3mZuL8KWyfsj0OTM
JeMT6Kjm5hneS8yZQDrj2WE8UPJu57vBni48uhBkT9o8zo0edwzTTa4ANu0saq4St3gLWrcA9OW3
Y6chgbqZyrS1VvokGBm9i0evK5uzigway7k3sXQhP8TKRjDc4Xq+tgQm3EL1POftFKNNAFe1duQh
/PbaVtbGXBcP6Fl0AuDMBucbN9V4eHvy5g2o76ZPN93KfIfdk7xSnCQ9xeWruVzMvMuKPlZTrJx1
dlHCYgWK9aO1MFVvd3PQls7OKcDgfYzjoKY7arGE3h5qbpujAJgTY3DpRQBcHWXzQrZbmZK2I972
sa5tsiSkdwRN9275WJsjIHlz7WkTzH8z1KkGMhzd/lZx7WhO6KygZsPM7QOh0XVTg3qZmmLyO0fj
h0iA7sH91QEikSRDv+71/AiZTYHOBX5P4TBL74bNVthd5HAXXpGv6C5jBHVRBPQzgAAj4UlrzKs4
WOz6TNJDnPzfKLt7YuPRYPBns2PAImYPheiKq0RtYPwwJv+s8bkPyug54KE6P2xqbLP0Jl0MOWSe
0dAyua6rZVp9VKpCIlbys0AYBuXG2tdhYhMr5Kch7UHs4m9URgCKtVvRfMihr0mGDWt9XAQHWrNL
6KJLcedhnkoV9xvGeYREZqPImdwxTZcwOOT8roXz5xadWgPAgWRkBBd4kdcSn+rD5AiVtAdnXZOv
wPQyExLH1OzH0NyqwjcJK3+6XD8BS2IHW9C3WglBLXMkP/D3w1BOOAxN4BRwi4o+fvnpRbq8f/D4
Yaj9/rtirk2jEqqBonokLWVbP2jjEx+5NwhNlz41Kq2jfm+hScF26EagIbOCbKezjFZ8ndKFoe7a
bLdO2nRa3MfZsl6HwTNpVrhfMnaRraJNep8gfD/Vco/lfSqqwxEJ/R87WfD5GtZfr+3h5FNRLVI3
9yPtUk3dFYlMsITI1omP5NFBI197Qyy5PAGT+QZWztKlYus5gfBfPDzpTVU/5JcKVdWSXz4Dsi2O
dZk3GZBQ165l0qU3LgijzCKRf8PljO9u61Oo5c5Mr2j891Oj+ttvXERnJ2D1XQ3W3SgTo2DCLMCI
yokgyrztIXA5XuEjuMP6Kx8EozfRjW7UznJNB106TlmwhtoMOd+40e8USSTYJ7KUv3ibxGPAPPVh
461c/qk0iM+rNeikl2yTwte9MGSO9Jqoi7NtUw60NIMko8tA+FYrC43is+yDykDCvEpB6aWcPVbI
omuelseIKqiFdZluNFzr74QgpfV5X8LXX7fGZ3CDTkktqb5m4OoANuEa46CO2YVGBH0/ObEwB14u
OU5+tCS0ty8K2DTcBaoB1+/5oDY6hhJynKcncofYipJo9lXDIeiXbsqmp3EOOiu0VFZ5KuGInfC/
Re7OWVAqQ6yMe+Km2p7HRAtxO1x/t/W6eLUBYQ1H4XNF2Oxn75+IxZOjdLgJw63YCZXw6d8txaOV
Sfsrvp+xPshI51MYdbtq8d2YfRtvDOi53UUa2+FjyTn+6fq8kWA7fHliJapmrHdbPAq+MxRvhQW3
li/QdLLy4p/6z/pkOhg25GmRtLDumT9LO3ASxANQycYtA9FbsHN7dMSFnzsovGe8xh9ApIvBUYb5
//v+LsfEN3gMHn9xb4zIzC7XDO6eKIrWEMI57Fo7VCRbZ1sYcjgGjLXlwW2age3xZqFtH1d4jnuK
Hbcw5F6KkWktcSU4+2LKWmSIcquGEmz9NjlsYyugLmCcUchXGvnVfLRCugNpneZsP6j5cTiLAJs4
hRtCwL6JW+HtCj5fH6vERnIMYskHhOhDcjmOMBEsDHJzMs216Cy/Yn6OethmbFnu1+mytyD9qawx
EP792QdREPyGsTZqnqYaL4Yd63hmNvcGbYLcmuCuPRxUnSp8o3on9VORnvepyXb5kGw7mZPBNDf8
N0rmUL8c/dCQMrIz54ctkkTMkLKNid01YMHKkzzgo6Jbhb9tPmDaDSW8YaDfIOiy0UeyfXBnwLTi
XFyXTEKAQYlZxt6fB6KDrQsrW6/4e8Q8eRRAf81am6zDj1sgFmmKVJDvqP3Zb3uOs4+l/YuzwJ9U
EyqPVbO4WADfZLV7ybMujEa1Wq66sMXPYFgvQBReBdnBr0/gKLVRFMALLnp9DsyPsV8q8uqyR5ju
+joleg3qn7B7R2OmbBwR5ufUEVfAv37bnDr3t0k2tQKHaQS/eOm7NPvPgvztorzsBfjVYeb9cgwb
G1Az1V6+x8/ZvSyluuPVr1HHgvP9bsuF6JxOciLaZtYJfnkXfuy7lLfkcSZJRbDt4Nvw65gnBrRu
yeZ63w1pU5Tj3z9H/hmKvWuZcI7a+UMmjsWF3K9Ee/VZWyxyVLUpElEFfUxCeZYaRdPv24qlyT2/
UKOBSAcsce+8Z2Y+gaKSbKXwIDy712xG4A2KCpdpbBgBnx22QQnUdJbSAkkEoaa6ubswH0qPCbBW
4C2tp9aM4KkKEAtny++c8OuAdO2/E220Tf80w6p1y4ZsENYQE/xKuiubSOzxVPVGg3TFr1WY371r
lCzsN80NMmdtnxvSiwxyHzwd8efpI1ORKRP8z3Olm2paUVE9GNUYRZSIZ5dQGMvhBTeCtMwnslrg
frpJyIVlaAisxLFGATRBiYlsg1KVbHogjtNKET2kWlypBUgweKtkyrEeKQ9zWZCc0qVyFbuGn7jx
YeJPFtpP4xGdgQxS4HgM3JlZ6lWf+PSJDu5JbfN/QXU14nyeHq6dtdzJBCInKLsIZLLf+8kn82OI
x4oQtDWhtdQV1yuAYsqQ/6SliLm96G8U6R5mJKb5J4qBfdMWoR3VWtn5X2zo3yq7ezk2LaBjO9kp
O4SmIAT/BS1BIIXMZbwN5QDNuC8kbTDW0US3LZ2iX335QVNtOq8Kr8cGgrpDXfAISUD6NffuVRSN
rQbk8Mck6VxSdyVtXpGhPOOzRnhtXuTVyqpV/gU2yeJVm9Mpgq30/NnAwfKWtrRBk+CRL52j97qj
PA7ING5hI2Woy4wiUgZ6wDf6UAdT26Rgto9jHE5c/2oWT98L2IpR2exG5s7rF5Wc7hxuzU8+G9et
yDPq3C5gSb2/ivdVMRCqwAHZH9LCRr0juMHLWiLYu1Drz8JKBWG2sdzGfTL2OMOYrJfnXQxsaxif
0k1m/IGDdwFrCkuxD6l+rdW9O+0quYo49t3uJzpt9WBo/8IwCcv00BPCd5V/hgGVoecwylWp3YqL
LLjfudOLfL7Tpu3Ijg0D80cpzbuZFo6poMxUNgbkZRGJSZCNqUpKhROjtjItYu/70hqMni3QBv9m
bHFE8tk0fV4qooCEkEf4bbFz5kxVavWk7Y3Dbnc6mATjTTpN8y461r3IIj6glAHmagZEdgWYVTTp
4aq+pppJVRMLaHF2+daF7D7fzFZqREjH7yqRodx9gcywwpQFO29vHUk5h/TV1xGCzaEfHQi9UuRX
K4qqAYFud/eEjtBXtXaDw3RorfIDl/8dLGdJMKtsz7mOewn6tgabpNFOl/NGEB9d1AsbPlhQ0LiB
6B06OJuIquccHr1iJErCKGRQxe88xFGEcZYaqGKe0CGndn0Zqhg0HFXEIlQY8Z3EsUlHeauNTgH/
VlOOf9JUYkewsHhQApAcc9a5+8ZC4KuFo0npYJswoGQuvylvLloo+k0Vys/MFMgAnc3qqpGuA8wu
dTNFBdIYaNeokrP54HCXLBQY1bzEbmeIhYEWtHh9YvNGjsUYaqbWyGQ6s4NoueN4vNhO/D5QwVkt
FLMbytMuJyEU9QrmfHqKkyri11b7FuxM4mNNIm8KHiMVaD4DORlxxIh03/widj1VOaUkpUc1t8gd
0oA2/2RomGocnveP95n42OA5wu3BSI9l9i4jmHhAYbWlEuK4SVwErdvVWq1LuFTO0Ron5X36JNxJ
yZDYQhhnQOhvLEOFtpfpKmYWllRIFXysapHNEdWbquRNgfwE0zq0EQ9cxzinzIOH4ku9IxE5PiC0
orzr8/beK82EfjqUz8jYl9foAd25V1XZMc4CUAjB6MuBZPng/17YeaC5T7cXC0pn5qkDe0zem0rm
7Ge0SiXGM3E2CGTYm8NoO8e5c5ae3XHdrxN74TCCse+GlJJmbVYlh9Uvv784qRgDer9yweM+yECw
ejfNKWz4GyjFc+Z8ZT/c6laERFSaOq5hpxYfluYMY6UlikNu16mNB/lcUlfBUZ9vTEhOWP1h83a0
2PWqd+Ub1IKb85XTvXQIigBbQGhPFoVD585bdsEU1C0Pv+6KDXVn0VHJVQOIfl24ZQbbrSlnmvRO
NGHCHOvSiCYZVpauoSyXufeO/TaD1EyRrACNKnJTNmIsBI+nXbywNoxDbnU5/elO9FwcSPoXLVGx
TvocY4WyH0F0hweknmT5mTYKmqwM8xFwrUTIpaPc3MrWE195MVnDOCSB//1O3Eo/ZaE7ceSBaNTI
Qk6z5kvWPEMH19TP0KY/QGPLE7ZMIZNrKHxpk2GTCIcRY1XYdF7nTz5GcLkxV/s5SUAM8g2qz8Bb
NH+RHle9lyl3Hyq6cSEtP+2nPPLEiemM98CzFr+f94MAL4shh75Ef8n8HAx46NGXL7chzgH8c4il
bo5sgKZuxXpGKR9vtnYCEkxa3NzndxBhHa9cTlZW1khAZ+L25NZL9PlJJle4G/e6Hko9O6VIq541
6jGbA6XXPJ7uGbBeSWeEownsYKh82eA3c4XcB8YS5Bi1TrHl0DXHYa/yUmRP9vCgro9VnWVqyTO7
QaQIdWHpkcIHXGWVm8tlx/37FLKtiG7z35olvHqbCR7UHSghnlwOuASKcfHOXztmGxLEFoIfOY+d
CU+HvqxV/hMivdRrke4YWGE9oA4RVrEEYcSrkbOBs8n1tzMXzdJQXA8dG2+d2m7KrWsFXmg4Y3pl
Fmy2v9E9C5cKAX/vAM6onMRq52Z2nlX/pUKFuRQW/V9mBWsTFmx5PGgfTtNTLqmt/Gt2LSurg3EM
NyFmyumrMIfGvHFgB4joJu8E+VDunS4R7AjQiU/eoHx90Mha1KWDjLv2ymnzMF7jMMQBvqWNjpD3
B40fHNUcu/HkOK+IDslJn9jaGIEiAzDwtCUNhdZcCtGl7bXEtTpUzZHFlpRsxQz+T5SWcIPAmMii
nYiZ+9ff26I4/mzxLDGEnRkbAdT5lMUKnFL40Ob0mK5tgaoDO3DLJ5/ng+jWu1zMOAikqpDANsDc
jPDaXQawcuHQwep4id4d56Hxr4ObHzavosPSNuEzllq8lgEH1TdV2nDAt+2O++WkCyLkjzXegkm3
icnX7VRxHJpbOf23cHVnhezYgcSAEkOv1W5SfehOKwMKgIVohlgzLMMSvbUNbFPuY7cIw1Mliig5
XMFRWH0zvu4D9+RoMHdQ5k39eA79I2A3uoaGFb2DTNUzzoyH978tO8gof7mqnMIUglpQUnzkwAR3
Aw6x3Mw2ZPNgo2Gm4Ee1QZ2iZZvd2ftPhYHNHa8e+HIMvuKbwk9N3ksLug7tSljXVyhBAP7+R0hB
XesPSjd0NRT7/cXkf4IgjmRq9KI0IDqSJLfjEkRGZsHt30OSYTa6GNyRAsbuDfIvUl76tsu0Wbhg
Et2EE+0qWmRIwLolytfoNzvGT6137s5Q/pYd7VHXKhadkf0tK1dEsDU+Q1l7hcNTj+ctv5VA2x6O
bWKuWX1MAyC7c23bI7fJiP9qTYsEeAlcs8JMafyhjLmOSMEOreH2Ojusx4W0mVhvL45oo9BJ8L55
EvmRI5HxPxHltQ4AMKomVElDTZbE8JDWYBTdzscrY4eBJv8s8/uhugZmGQDqNl2Nqpib0vZvlZ+o
gjrRLsquuUlS64n/gBRlx4CBmKFFdGMHAA8TLPp8+QtpUATLsBkhBTxnn3aI/f7n8b7n3C42dPvA
xsi+cyorIvsJOWarSsJLyUD5v+rxULs7kg43tkf0GSIyvKh/4aZMKSRvKQr5AVoQlgMmr9YCdi7e
rSeIOlwmRDoujXGvs/mgLYD4xPLSLPodTTKJ/ddkdHpKp9oHLoisNuDQiVHXmiriPrcVL/tPAwa7
X3lKSf+cR+XoXaXVge1+bRAEuZFhguyYZ3FJtG6E8gUs0oN9PapGL2oaaAMvz4kJFPYF6AMhTDCr
kLDdCONVH+nQ4rm/6jq5dGX+mQymd4wGI33XGzaUSAoRQlLDtWfZuBf1Zz8vkG9Pn7IDV08Ur29C
H7N8gchFJrKxF9Fg3qwnUw4O2ur8KKOmu9p9AfdplaSi7q7zmmq4+vGWzOry/uJkGBNl/KI8IIRL
IGwtnD0JpGbsS4OpoajfcQShzhycHnaslVCZxEgiuYMY10H1SfFSv4unKyyVwUd5ahzipHX3A46s
bcQCzjkNeBDKZ3/7LIpVGmuJCfXpmJ/6sBXGbE+CMOtTQttNI8TllCMjAeWnjUdq4p7nZckU5iRB
Z2oidqUxKhPy9djjbSceg/jRV7I6Iak4ExS1vU3k6iO9mCz+4mzm2rRY+vxSrQNBWS+IGetIXSD7
IOcwlNotMWmBDa0t3Hd8+oiSYxCg4Yuwn8WwZ9K4gcg7PKwPNjdhyAbwZzVX/63PU75igybpwH04
zIc4CinWNLnyWGf81XcrH/X58UlYCG+4md0KIb+aMdy+wMYoIaDwexfzGpqaQRU4jZtgSe87kDzc
s/sgLrQZZIAFBBCqt2nln5Kj1TB4wzfZJ+jJoQCWeo5SSvB3NHOcIck+fo/T8ODewn15Jhx7fX1s
KxvYUOk++11ywwvYUjj5D5pqNYtUc1NESXMSbV7JZWd5thfp6shQjUdDeQDnhRhTtGs9a2wqvUtV
DSSjX6YIj5sVkmHX+RRrIMTIDQpMHrdaA200fC1YoEXdUZqUw/Y+R96SJFhVtcqa4t4mRBuZlb8U
0Chi87YK8lVs72F3rXGrRH2Zx6JiXhIril0BijPlhAd5LGwv26Tjk6xFcluurm32IcKR+591I8QB
IRis3Yrp8EJnbm85QZeNMR/GlZcjhwujkXNG0tnFDl5tN1sLyH7nE1T8Y2+MFnR35dJlxOsAfwEz
L2QNKDkPe8FFNqcGQ3thIcOJvIVANNAVjfpWkLao4C3w9E8b9gS3Wve886rPBJ1kdZ4Vo/D52FAd
8IiVYmbbnUNXJ1CLx49l3GMAitgKWuTuANhI8NzEm7nKspwxk7+BeuJTBUvqlFEgG6t5J96+N7fx
eV+ulEpXTm6NQqhlPhyQERBkoC43m3d1uk/9z9nToB6xAGUc+jWisbKLbu0Uttdh4f4mWLHl2yTq
V0RfeceiB0r/ajmZhnlc2qj5n9U7/KTh4ormzBhQDDrBRztE/sKuQH38J+A/5V041KaN3enhaMFA
aEVztIY69sEz83FCMBeKvUpIlvQlIHuJfUM+u42LRDX926eVFvynU/EsyOogk4VI6VBLAiL4PemM
0+iOpTKHwXH8QLQC8cFWOUq2OpnqKPK58san+wdz5R3csizmq9/yfWQ2Itpcg8zl5gmITHOwNMMH
QCzJ94qQsjXMAYkpOH4G0gkgkv4nBiDRSYpdKnxk8d7sNYWaOnt4FMfcbo1kIMEQ9O/JbCABrp4P
v10+IAKQFoCChmFpcY+vW3sVkq52fnANheO3YSoCfj/qHy0H6V9ElACjeDUhsTyGjg1lhc5ujp/D
3W8S84METZXK224aiYFT7Cp4+7reic6CCgb+9y66yjWJGBoL12bpHrH6CdCvgSEh/NW0DoF+6I1B
2XwUvDhWA5PmwEUwXNvzRAZJeHX99WKz+MyiADqCnH/DYX59oL1hGCQNfTdsRTUzz8zMTFuRiAXF
PT+ajOCRoN/OTKXhy0tLoO6/PPVjagbeo3TiXbLHq3jC9rC+NbivpPyC0UDyzJ8mzuyXf7EpchFG
AX4BtOi2nu7jwwHxgFI95fn/vV2jLelyGBpXdw/4TQpmXNVR3h3V8aOSWGcbSRDiBAyQl5IWUDYK
tKyUcZ1Nt8N1Oi4kqHPyg1Jtt08gsNk8M3xYazoLqay4N7FEEvP2t8xajfL2YlK4grrO0ws9KsIk
/Cfa0zYDqGE0p13v3pIdkzunGeIdFkvq74qYF5z8S0IFYGQB/ZY8fju4uqxG8ZTffSG5Bg73pzxk
xj2zCHbT1HrQiMPADbgsUBVqfehaCuoDO6f2fTsBe1PZZa2s+pUekPE+s54tR+GxI11yNCMktmHD
cdcZfytI1Cvrj7AX0ulDVEWHhUlVXwgTR1xyV1wCkJZywE3KMTu03YJznXh4hzeTwBmKKfvCg83Z
4JFVOGoLBztxA+WrssfKDa6brqD46+mPTsDBu91BmcxmtWlRM5YAWxlIZaRiCwQNoln0SCfIhmyg
IPyHTDpI0epDespDzSUYf7ShuBkAMHZlbXWRLgHMRZKEzyCZpxrcUIeeGQIact59Ih3k+JfI001m
tb+OJUIAKwceH4HcdnJvAK5It7Thn5ZQnSHSezFhRIwNZVrPD9uJ/4DvzePivRyUm+a2jEF0Hj6F
QgwbIFHUBdYKC6dy4aRYlq1fOsn5vY4NP3KBwPM6TWLjMUh/qR7V9gXod0CdxO0+++qySkHUeYjd
t7B1S54DDKyFb7fvzJ2BM2yZGXqTP5/ME9PGCr8xZrbvFTcAXGavO3Wy4lEfqAoAk5kETSKT5HsZ
eNZiT+rFzJN2+YKRC2k3xfFL+Gh8JJxGXo6CaXGSZSj257B/2KK+jKBKrg0aNOWjoiif/nZ4hoZl
ttykTxxVR9smC3vOywOsNt4w3Q1ey4hj6eAMBLFC4YoK7mBFQS5+IOsGz4bvrZQ3lbgYdpF4Qjc5
vAvkbqMoUKHdvxEzUsqKLJupOmlmvkU67Qt3zINs3z7byUkXSvGgVw2lW1onhjkVsC6ZMIJIGvAa
ZjbyE7fkEGEwkOyc/ExI9x5VxQugWGLXSxUsdaRWFDHxEPaS1auXr8og0OSwSKPKX5UUo3Xl4//f
E5dSq+8uY/Dk6XgpnqKASIYjUc3UXb0HozE+GgzQiURCP3NQsurWg6iS25GixxVVPggyig1NUHE2
R4o+9RGm2jHQKPh66lQR1Vp+N7jMgV8ZhSbc+U8op+y1ynfGoZHJVSPSWZ0Lfgum5LYfNErzd5Yl
Mmj1SnNIB3JZf/OTauo/qbDWfFoRmmyBjCI7j6p+wvgicMIM9X0aQv/Nl5DT8j4IrFdQcAvZbpSt
SnJU73LCxQ9/JyJUswoWvzzTysQO93ZfQXL5Ups1zYEgRo9oH6n7fjmB+s5Y+j1RUl+W+VwQwpXj
CeV5mExJ615SEZRajTu7Q5j4ck2ONdylJ2LILnClE35eQBjWwJXcmSuh+8bI2BoLRUjEIHql7aPn
wXRrmnrAXNSN65ZaXyWwl/DdVeDITRweq4ws9ZqXr9IzdsHJXwjthgLY5F+PmtOUH9SZkI2711ic
n2R9on7IPsNgJO0SrMhtqavrya7NdJnptqSx/oO31F/lf0wIXvA41WwVyZ2q7Oyal7z53JiTI6fs
aGAH76OLDcS9mXm/H2VeJfBzgr7m7OVgml+7YCRbXWEWmTzN+gsGiReXwiLpECEeO45vgm1P2h48
hgbjylQyQvEuJvXVdpR3Ac+4DWh6acuIsobGnxu3096tSD77wYp3leDjNikLM2VnIiYLXDwiGIqa
S7pgS8aTgMWOm6nOKqBTYlQ4DUmuJiu55O933UqwNBkVH26BdJetRcDuJ7LP5oMlX+fKlHltBnDC
v0VvuycTmPxgel5FSLMZ73oJLqAkJ1DFyVp+SgskKbPRezt56bATnjyu9+iriz+NpzrF6lIfpuWU
hZmkDqEo7CtCtEPGXuiLTOQa4VOYiAN32ywyaFX2K7GVtUy0fZNpgWGZ5PBNTS+qpuJpvzGV2u1p
HeTEU2BTd5rZvujECO02/nM5SY5HUBrtk9L/CqgG7IcE5hPslOzbcXCu9IBvYkhpa+Mo5V81Ipm1
JhDwvb44p633qsrTGNO0ivgDpMcsxpBCx5BpeMv4pKDzN0fOK95ZUJRYGoEJHJzKPev48cAYMX1x
xljg0aAVaI9oBuaD/nTtJK/nmaN4kUF1WnwOXRGOfb4Pcrg3og9noKAg6k5W59DSOx1RKLH3a5GB
qUaTZbOitK+0HLKEJ+wzZbweJJG05HFaSS8/gJxmJaVtoCO7+UOMeojCBvUst8sHhJZXB4hlv1vr
UuvSV8Na+5I93NOFWZgZAgwI/PzSLQVPcaK1RMkfQQJ0hjDwCmhH0P/akCQ4GlJKEoSu5dx/ahWG
NwBq92qacNMcHwJ+rB3piCDo77JqU2bP/WwyYL4gRAJMQb1VbuIZrONo7MgNCpkHlA+lXXwwAG/1
9SOXhcLLKMTiBf70HSxp+Z3GDVDHuzmkPt4601mNEt21q5NzmpoG9BN90wdw4yeW7iBs1SXWNrul
/vwhgyOqrIw0H/n6tl/aUAeYoAAv8fcPWjWXWF9JtmY1mZ+maOD6kPMHm6VM9htbNa8q3Qms+F3y
zI8rPtMAgY7Xx35/RkGztp1heJD9nN9yuhHr7LDFfdpAFYY0rICpE0l5P0xYGpOi1V0QuVVwRLRE
5RZmY/KbWIePiI74HhxztdOp6ub8khyA3Jrt0ctYCJtRWLc/ngh3O16/051PRm/MQwewtgn99wT9
6W9xd7fYKzrawS2s9LYCcrz/sL0KpnITnKLlPhqmeRsOnYK6bpdTYC6bYs6WwD1FbVXwCl0oHCaP
MbjxN23ow/Qz/uPJ7mfZX3FnaebYJ5EQt0yqyh3HGSOhF2AWljfmw0Z0I14Y59Nv5xOSZbc69aO9
bZMh2bZk8MQ2f9tPnDPg07JulgHhCKGXmkeT+0lrNqW6lRR/5MvUVxrVoxAmRlbCm7OleG4U87Bu
dZMjHfxMidvTq226oaBIdUFVqA2UOeCqSON5FFGE0hwRI11rD/6vFxDPC17jIu8djd012ozPPKwE
Dk1zMKf6+9SQJ6SSm5CMD47muxEoo5I//wUIRfkxgOcx1HDhjb+WI7cW8lJM35dLXMEm98AGiAGp
LDiFAylTrQ8yZx0InBhQwpe0+L7n+US1YnhoJWv9gav1w3hIU9DS/9SEg00Pd66kPo5BqJOQTvhk
6P1XmteHRmjEVZmyDoebOjQJHCOOA1UmduUi6CvWQaoUvJnS0UGDFzVpKtWR4NJ7orXK6Ivxzm9G
KeaW/LPU/K9VQzkox3YnkfNGlfWBeEkcq9sRX0JRq0+6gHE+wDnXa4+iFBkqpyihFM/yOUMH7SQr
zW7zt5EdHhKPZ9JB8NR6kp2k3NE7Z61EakJPNR8u8wDfWMXd7K5UGLv1a3NtDRxw9QPIfV3bTrwb
/BeKAqOVVJeLNSucYV08nMl3hbG+zb4ianu4oI4TrBjAKDl7gQpzeqz6lAGfarRsonz3ahvdJaw3
HHDZVSQjpzbqdrunwcTF3cViMlm4GFI6m+a181lpVSY2mmqGIGreuvGkUmBBo1mAFy8wOpgUXl61
PvXyJwi/dL0bE/9m2e46pP5h4j5GjIMblbXp8po5ETUqvVPBezJo+zpir5l8ZbXLVm9H0QTYR1Gy
QNSPh6KuRlC094DlVXpgo/ifEc+eGaYbpJfw4/SdF4Fp1yG4e20mOBqwQvkoXmWjcGS0h5/pZkRa
PFrFaJKTq++YK7pqhk9rWx5OPr5pfnB/VKG3rTXWzHJLjhH8nW+1lhBZgt68VkLwPhDU2T4vP1Pl
oCG8fTkE1j1br4dVnsgB9+qrXE+f46QTL8kaEL5bp0zsKa5KNKPlOn+WzKbtsHRjJGRCxhZLeUOD
+c/paUzXkD53pheHnpxZNGRiZpzgp8fFR9pJGpC7T5rh13waQ9TBEiHlg/1LuCCaW+0EvEpmBiZv
+zpdioBwyaSA6LTIE4IuZryjmqczsQwPaZaWxZp1ZL8zeL5h+egRFr1I5DNW3MKJvTrD2M5B5fa1
NAed5xM9PCWXCFUogC8MuX+Hc18HJemhF80bXJH7YwF4wLc8PReZQoHzfIsevqP58w09VATwPI7d
ter0EupH06UdPGpBIGM4ToFWOxjFZXOD/1b5iwryIoWdBrUgjH1YQ4aqsWvEsFivZt4Tf59SV7aa
PksS9IMwxrJnOmBfKFpOOFMz/vCqVvTrQGIZVvhmKVrCiMoprmMolE4oBgE0Srrh6zmEsTMck/zX
/9TXnl1xuQZjKV+8H3srOkiYbdw670Z1/wusjKSVlOsTsca4PkzijkteYMQD8NueJg3y6ZiyFzdt
OOkvVB44AI+RiueJxPydnUQmtURnjg2u1g2/ej3a11MRKzS8vXKr2Q9gLrzIt9t+i64W0+qEDiVA
9ZlkK/Th+xcxW0dGC6gZonDCETotWh+s7R2kr9FQmegRuSTQY0iTyCjkP+vZg7HI6XFJ02KuLKxD
dHNTsce1b5VHue4LEURxxnKsmN2p1btmDAriM+ivxBR86VH7X8J6ZsmPHtjzJvvHTKCn4gJJjh3y
61f2l/0XdboQ6IdTnxftTIUowbIEFPEKKwtrR6TRI8/qXg8XikATrF9QiG3osTP0KzbxQHowftvd
rDzY7xciNtnzfBJWd78o7CLk6rVQB0E30OaNcbLgD3XeLnCLKDh42rIjdT3nYMtWYIw14NFftwuL
biLxBvG5cOagHvCaxfvfP5d+36qUNcwIpSrtVA1Yu8zDq5hINBxo//17tPSpIUGHO65X3aijKh2Z
RHRn+da9hcYN7Fh5QW04gVeth/B1pl06fFSW78n/UJX5BTwcPG5HlKv3BgocdwqftMAmQ8CRpr6S
fRjOCqF2pukGufQDkaYsHVF7jO5e9P823uWqWEsr+54JBIo9XFtCwn7+02pw3cmwv51YMsow1/ad
TDN2kJ0QQ4rTbDiLaeaho0bdD5ikTrTLx0fskubXoX+5nfgCvltC/WVC2zWisSpv5nQrDqWDD7kk
c1TxSvO9Xzd185gkecFzmgeupeIL1hQc/G66BnKA+kgbz3vi2iy8Ng6Uoiu80xZCs3/O4MR3TXcz
WEHDiUyf3Y5BcL+6Poo8x6d7nLvJcMPvuXMQ9dL0YJG2FAK3QVInx85K7OH5JQ4zP+pKHCW/8XYO
TN2IApe3FH1frTA4UcST6XaopjVQ2hV4IA95328sNSMhc4gE7DpHWBpFMc337b1b5MMXh7AI11qz
9nnY0kM4x8tNTwVutd+0XTfOYMemB8K39g8BdJVW9ssNKG8iPy8xpGYF5i+jjpRUyrCQN0/a12WO
7KbRcl9/9j5juSsiKP0ZMLjj0c68wEIA9D1S8RysXWT9DgpQn8BCn8kDAUPg3GIWZW3lql6sn20a
45JsbTLA42VPuX9XMvmQn3zLiAO52bX0EmdxpWILI1CRxd9FF2CB10XvhbKXKiA4Yoo0CpsBS4Z0
5c6FOlqpogYhGK4oy53W9sXX+QF7jlTWrazXBiht8S/2//rW7vCnzwgoUaLJt3J5whtX2I885EyJ
N05d0ijNfqfKjAUMdYvP8E37cz3raway1EhW6MQrNC9LwAScu08k12bcH3BZdAkh1wEOpjgzWx6p
aTKrjCSRengRidgm8Ov/5OQIuKouvfRqTX/saP5T9p2zX7j5vKnKirLdNDZ/Axn+QADq9f58gBBz
nuLGsQW5geJtB9JF+wHN9YmfBhszcayImkXdgLauerdwRaJ+pZ4mnRTDjQLLXds2DMVkELToR3eZ
603WJq/zjTRul+pz61w2wGE4zWRDAlkrR+5HnKXjxoaiJqV1n0vR+3qbHIEMzvyZxIzbmpZOh2X3
epj2551ZYRaa4oBH9HJgXUip2YnXA8Q9zzLF5ZKwAIKSZiQL6eecztc4NQNBjfSyucQKPIF2PZcK
65ntjdZiqyHhiuIMhCwKBLywzNE4RHc62IpICLUoKs5xFZAI5XJ9I8C+noZ0A6rdFwCDPGnS/Itz
OGkTUnFZgrNmld0PtXo5OhoKiBxU+22A5akXPGkj4vjje6B8i1Ydqd3mcQlaPgUNc2RU+5PzN7Nx
fWn/qR8Cf16OC9TLFiS8umcNJ9vdJ/oVvlE3ODVTB7ydiQHZtgdv+JTJlDoF45LZplaIWJtx52rt
rBY28L1isV28KertbqE2jOEoonuDRxaHUcr26m/unj+zny9U1vuFtKWNwTikBStH1XY90qrxAqIi
ZjFfk/Ul2ytXvVhOZHkKKRsfL6Cm+vm54zLnNgx48X/5J5sDoOaDFpN3h3ah60bS13VnWUSrpP9J
m2DOIOjtKIDbV8XPpr5M4AZq8Y9D5GCCLzIQ5rpN4BCUmA/7JPTayy98Srdh5ba1hsiVHlSa94aI
2ihogwwregvlfbJ8hwl1P7MVJZCe8IvchJ+r2FoMYuRLrxSiVczlJtb65emSiz4h3T5+XUCPzDrN
kRbuLbfMDkead8NNn39HY0Ul6qNvl2+mu7fgYCF7cxzqsxVlwXEuzWBDlVgV0zso6XPVUSSYArQB
OY8Rk17nxmCoM++dSSnfW8SaH0cxIu4D1187InhQwYSZj+i9P7vuB5nIBlOKsSPhBki6D4s+ouKL
j683wdjEYM4WwzQrpNXs7k4fnavmXxYCc5HJOYddYcCsqNn5E0odBJFZJ6y+Bswzm1rAfFSWSTe3
up7zDhpoA9uWBSsjdWS4lTqajSmLmghd20FtQeRgNs7Cfuz8FV8aJPS3PvUFLZRdDZqfeqw26bkv
oTiy3m0N+WCqOGxtVXVCC3MByzmIhaEONnaStIpO1ht4iHI2HnI9eRsMDn2KhoxFFkrOJZCqcAe/
dr1e7BMyNga6ZmN8upsoP4rc+NeDvtPCn76+DjALwCaeF15jSpuhbI8bIjFOKJAK0tVgN//i9X6v
a4U4A6CSg2FOax+jIYWRwaUL0WVnM82fhmM9nLL5GWRcKWvIgw9iHvEAa7FPmLsJARySFAgggfET
2Fim6S/3Bx226Wih6WjxQoUf6y9cU/QlpFzLg1YuJMsuuT7xBmg9A4gY+2cpuPnE2UjhQNJgbo6w
fzE0sEF2UFYsAz5sx+/eCn1HZ8RgMN1t8xip2X2lE/Yv/GB8muvL/yM+G6pLG7ukRqUcDq/rGV2E
ITmk67Nnx7KHojZhf9m/xV3zVsCitMvuPq/jH3hefl3LQdnpHE2+3bd2YzqG/LhvzFKj5Ia7sH7x
tL+rq7DEGEmcTaJ9qibK2d2X+1yunASr5xPFey0XV7kF0uCk4Q4One9HAiR/XFep1FLlIzg+dbe+
pUdLSR3yiD2+wNXdscT21eVtB+SjvnhuOsf3iNyAbv1nibrPUXkxyUke08MQCdzLkwE686O80CdF
RI4L16mVXOtR6mpLvtKIO8o9jKNQhp6t7FKsR+wrOGQPPJ+Dwyf+u5/1vjGEF3VaMJ7VOZLmwxJN
+M6mKamqKrJ65ETwdABv5ReodNDDGCVod+QBNPB6msSsnv1Q4CkFLZrcGAlkhJYu42UzR/RD3aU0
Q2+Jf3w+d7fSWb+k701F/fDqGAmfsETuOwwbY5nUchnsuVAgxQKx/OEEkwXiG2UO5khK3E2wwHke
1VdiSLs5RAKTTAV2CpJgId05T1WHPavNdJlD70jqZH7YEc6Wua1BXxMjDe8Pnp7O2+xhYYsYohvJ
KHV0LiUE5Rxej/DV56Virtc05YCBp7uJAopjxp1YoAH4eW+DeVR4+uBS5UPNKNa/BkI8ROPeO2kG
DftDLBIl9fi0mAF6cNvFT6lfjjyr7rp3b1iAn+pP2BWpa7fc8T/bNrXvZ4VIsxPnz0bFlztQ9MOl
px35LCbW3wZ6dU6Ijv0Q5fsVIvK2Q+qCt9orQEnYA9/+9j54CBAExTAdUqNqA6S6X//erJm+eDZ6
9Pxoufi47UNqFPVLwDG3JYGRYG9kI++JGw15S/BElURIHZswAFnejiwuiy0u5FKOu+lh+Br5WQNy
99dqdPo+26KpvWDU3mmSUVV5x9/0JbdlDiOSxabsbsfNTeVGthefFWA87X3uXfXk7wynt4RqMQhG
270EdU5FF4KQbXUBiAraN9GHiXyt+3dY11AXsG4y3Owuv2jKRI3ZOPEYkgce5C5zLv6pH7Bt2hmD
TjNvhscfEtLNnoQ/MeDM9/IFDhdj55e2z6iJp0PvykXiUko5jrZFw5mlLoVjoUFhh0xR7e1FG7cb
5Rv4QEOxW921tJv93/6dsLsYPZJ9lbQVN/YOYXjdGrKvBLceNO+NmlpbekvbHGgzNKWfDDZPghF9
0UwlOG/xbaZCgsKlyqMPR0PvklTI5DaEZVBBmRB1Xx80+8dPcOsXFcHLwa3FOVDaHLkDEL4//Hfa
qToCkgMeGEYn518DR78IRqDQfG/n0F3cYk2WNthvYudy2ZzTJE3MVw/DwSgcCUV5nF3BjqH2oP62
fPy0IjedtJ+3/vIimKpSgmdmIliF8bDUocX3dN3ZLkVHOqHTm5TCa2eJbqymFW+5i0a+wD6lu2oi
WIxg4hTmVRhE9YYone6VAo61H/2G4qyzs2F/uxDMWmH8y05eMkLZxb70uHsv54IiA0X8GGnBVEwu
4zK25SCIhJRQHTiwwqHVci0/cs4oV7b6f4KejjiHUP9TF/DKsK7vZk94D1sYtXirImROjncMs4lT
uD+vGnruE7VXCvXcA/5Qp1KySutTnTwo1GQ8/vargATBZbU6gw8ERf6+eKuMaFwVDWGnaVZ4L3Vp
d3/P81otCsSttSC6D2ogjk8/+bQpE7jyIjuUW9f3eC2kMRDnlESgyNLE0Bbm6fK6CsF4iG8DJ/8E
HjLy9NlboX7aOMfrGYQQxxmd6aiRY94ho7996/gHDkILRN9i63oO/6UkkWm+uxUpyZ1CqnuzNmt+
oTtRQFjdGZ+zRps/Eqv6QCp3yluMlJIUscP84nfJ/by4lvadfZ7a+M/u+6cUZFpuJE2CeUaLjcqy
7de6dRxVvIvMYhB69RKDfuevbf1l+E5G+CEm5MoCLGCgpWd3ewS6Kh52rUrdh0w3fr3QkBspSvkb
71jD0muqiJwMzOHBNLDbEn8/79s7BwMRH+dLbmIDCbWfV9JWl3QQxgO1PmQkRRB1ZkYig6/EJzyt
+hFuRTKR3DZ5sQ82Z1pp+zuJKDW7HgfPuZtEdZKDpAT2rsN5Qqj6r6ArGt8LIZ2P79b79P48zS8W
RlwXoaCp2EaylhrxGYeFgWZxmqu98PGGA7LkcIRsQEfPfu5UccBJjQH4AQF2Ir9WAYeT49RGu5A2
Ul1Fan0NRBHwekELjZaVklzwS7zTNugFKiGULRx8S9PTRelOLTkOv80N9DYITckOhjYCDJdJXcV/
wDYq7ExW6iKkq2YLrLggEMLAeJEKPNt0YsEyyOETkaD+eARldo7ZAo4VTgxHK41Fk3wRGehEx3eu
4JaQJV2GIzDCLO0TIQcuRNddmvxGWnAhZr+wkNyCN5dJlz1HLahmTv0+cXqoLF3Kin9hygtrjrUn
vEYtkNDBLpUVyipHEQFGeILdJNn3cHHsVefAFbFkunk08Popn8t2ssEJN/Mzp7gBGuHgRNZWItpb
6SuIMAx3DhY9/n+ceKvzQuzA3LRXGL+9hvB87WQoAcY9Q5SjSUQntqgB+1spbBpZL4h1/v+3Xr9i
wSDQ9MtCZ6SOml1C5jUNMlJ6xSw3OwELL4/V5JMSaXxezs9FVcQIiLgyRDrDlxAoJ6MirA1I4w2w
UVb+5cpxtSRZF89H6+HFq5JaHXJ66Skxrfd51QucXZLr+TetKyC7oxFZm5RUxkp/A3a5gWAWOVIT
/5OvsfQJBd3MSUEorJPJLIFjdsCNZgqbnkHoLSjfYWlRgRB28bsOytkuwoTFQ/AASsM1Bwk/sgl/
3Ek/A6TU6IzqZyuEnPAULeXrBFCJZCU7DU4FcDo1M3Gs1B2kACetv3W96Dzi3L6j9iMrZSaacH46
3UeBiD0ehp1C3P5H2rHtOtAwiey4g3P32kD5qx2HY6nfzubv+SHfr5Ysidxc1hWQQXjT+io65zKw
fhRrM7gquAsO+WjfoX7UoQ39TMs9R8wxX98IGIQTTzoiA274SCCwGrvq1vZ9QlvFSAIpj7AzR0Cf
KipSKHyJKvFBd17URTHRiqflYR4ECeSl7abEYYBQqenpkkE4P6yjAfNsW21e+tK/w1SEamarFryZ
J6NGgiUUmnLfxVRxyDGoSkEEm2FzOQQZYfNPf3i8UtWnUQRPtGCmThGfHNc/MtTBdX7f/1QCMawT
AltmWFmL7d+5cDmxs0o2R2wxEUu1K8vbewmFGl0hOgf/OLplSeEJYfGSY/r/y7ytIkXBNQUzAT6r
4on4s5zestrpSQc1jKDJjewTV4yJqciTLn3F+e8tOcPWbMgIuw0lAK68s+JuF8XlAa+3SlflZ3cM
LSfq/ObH5z4gfC8h/UuhCAuKEoVYwmVEDjfPcmski3usoLyZOWjsnqOsnBc0loM2P0D0bIc+c7nd
Oz6zOfPOHRbhaXkSvsU/VcHHs5s5HAlY+ai8ejN9uhUNQgDlBlIp83SOlOFz//m4VDrNF2/x8ZdE
GcRa/yLLyqYb0oMT0wEpDpz882nhplxahjFDuNMPGA+RQVLzenbuhFMm6OXHXSdh1jzMkhV4DV1O
KcxofJFgPeQRjVTC51XfpYatfZ2I0t0LPaHacue/eF8jflsM5P13ofTVoUn0iT7VZF+Z59xu9DLL
5jT2MkhZnrQ4+vo1130Yv0CCHbmok8zV6y4pCOs/SnhpXmZxIAcCijYQTTaqY6sInwSgLAtAWxue
H4ch1HUfzQ+S011eWwN0yrrYAV/P803Nt9YTdHNeSkaShhEx5EHbNMbVEJVxU/jvJOPBKEwfghye
eqeq06a/5RNHgeOLwg8GJYzIMjJJzP0Lp419bXuKU1AjnZWg5qVmAIpfpmYpBC3DOadZDZzSj3VR
r/13k/OMZNbgO9eO3baLqihX7/WMqBon5p8vcBTVi9/7B4Ty5aCvSkFZBhs6hjC1mH9L5HPFc9L5
Ym8Tw2BokKkrgpKwOCQ9Iq7seMcdsbhhU8amrTPiOMnk8TJt0SESufnYt/iI9Vt3+XSR/g3hpNVz
dR8PvlrGeoXIDCzCo9GDZKvpl3EGUIq06rjIOYWhQtx2v4AnurBg3AMs7qEuWvIYcbOlU8FMu86O
xly3aGu8464/DVnvBcf2vEW+IJ+1deiQaAUdDbhZjF5+JZZ07IrlcV6wkZEUCen1s13wPf0cc+KB
cdDHHni0h1IJdSQDylCZ6ulKq36+g/hHjZXICRcFWarMVAf6N+t7c2ghYmeTozfEI9bJo576dYAK
N1Dvl66JHMKooPSzvNCzERCgLqrQSM5Cs+EpjjwpVq8ogfvGc9XJHKmn0qBAhsYnc567+3851vAr
lu6VvrIECxNqRC1GBqu6lXmfemVXjtiUQH3MfsGpximT6ulzBmJxR30MZj86FbsRG725K1YS/tJ/
ATzP41+rta2FMknIPszF89r5NRGSu3QAICXbfizz/YO1qXaUwemLPwA28ptgYg6T8whtiCUEMYt1
hbHF9RCazR+X+EjPxmVZIevEktxQcYT6apDGK3ptCvFwJMD0EP7lv37MylluaZa/s8kQZpCruQ/M
J3k0mO1ThrMCNoonBbop5lUcmffYs3kKg8tYboNrEDoKO8rKkeB1noTFCBGWaLnG4U51cafyBmFK
TKrrH5KhGzFfVROOhJDu5d+3n6DIkc6H3yPWrSqCmgH/ZoQh9a+i13yNbHE4u/FI8DhIl+ncWWO1
DzujsgcNZvtNajtQhlGunF3gGpN3XrlMpN1sOikGB5WVPrN0582ovLYyXtMNXZ+kRA6VMLo/uV1b
TGdpJ1zyQRr+eCk2iwdWbK9pF1jvm5GWiO+RcmPWugFcmS8b5pJOk/1XTPeHUCn1eXgZTXEOQGEY
58P7UkSY/UglqR1U93Zt/A55KVI71XRZhf9Ujbj58F4vj9vXBXLBOHAnI8CIyyCZqTTyHMpLbWZf
Eilq63PUmDJaipSjkOQDT94vdPLOFrbSX2Y8iXFwSdTZutx8mClT4lCRIuf3wcak5ibiukW73vQ5
VbmH5Y86aC0XkuFEImPj6kYkSibYYcFTGgfeeYLBkDtTGVNLqoiFmk4UN+8ryEQMsu9U2VivhK2k
I4bxdhjLAJ2t83Q+lLUJxvbAX0o7m5u+6g/8hjkXBtDJ35DVbusf/m/B6eCi+V7gW/o4VZWOvz6Q
SO8BSbdvJrZoowaqAcGgo1qysRjAuVfOC3z3V1PCiOxymQpCWRT0pocm7pgGdtTSmwJu0nrePeX6
s+FvwXprHxB1ZQP4L1blNo+Uo4tlpVEv0nMT+UUwm3gTJFdR5viAA0zq9pSvUhX2FB4wRtnl+48F
GMr/na9KfvGOtiGdV+40WnZfIP7yw07RJvhJO26K//SejyJ3bRlq7KxZfYt+8DmNtN98kSWR1wto
UY3n1wLSkX8034yQeAsTUuqGY6gXLd9SwuRizK5DhNZQ9xJ4QQrHQ4UoDgujvfbH8wD/BZtrJNMc
t7HAZZoHJQ4yXLxj8HrtxK/jRjlj2cvJYJWNORSQUrGZ7V6yknF0lfKMgtEAiEV7xeM/j+oAaY3g
BMvbfn302kA0q90JNMJcuKAheH8jIhKReDHWPRpjXmkPZNpoXH9tuWRPQWW0BNPqZYPcOpz9vZHQ
XyS8OBpqNtBEy9oisJzdVq4T8ipjRXHmEwQKeUolYX/Vf+bzm9jq7ycVd71iq+wfpZXV9GCWAXtB
J8ucYExSCt9e2oTms0eMeLl0zZKvH6aFUtK7ymD81f4yqzE4+sb2lVqCsfs4r1jsX2qtSwywHPI9
HMMBFgURjZNGfLeqqq/tNwnZtsAD9Aw2O15q4cl5E+ViTjptVj+BlRGvXzKVIWzZjYACVJsdcPF9
nwJhSkZyKaW0afslGmQGJ32dTR9smQHTvxw+IoE7XLnNg4MvJ7g62G0t0UEUsLD38lzcJ34Tnnj2
3w92iFmZAH/iKe4vHxQoKwFc2r15XCpwhP41ckDWLJbPAgFaUyfKus2a0tVWF7kAbxbABZwfaLpL
vrfILnzGibuEDih3X4C3wHjdok0DdaZYHH3L8iLPmV3cttfau15lsupwmQz+bKIApeEvIE9Zu2/F
AbwQSSfKmF9boE6SSg2MWZy9/j2z2YAeQEJoU0fCEpjQuYffuOJ3Jjp1N/LjWq5BUhqn7CDlm/gk
iJl0SEpcu1eDxcnP9f3GRUnOLytXJpDxdxfwGAIujAx+F+DtjAVrZwBlneXx4oRY36mtwtYmE49l
lN4RgpE4MNlVULXyzea2wr7Y3pBcPrBhntkjbpq9gizmu3MSfMdAQcK+2rX/54jSbirPliBJ6Hgg
LDJ+jHQho+vBFHK9bOeYxSX6u2lj3NcXjuM4Qlebtv/kLAy4go5RIQ72ctoU0WfqhepGwaem2oDc
J6Ml/l02wdwd1T6EPuEpiH1xxu/pho6Yux1Gwi9pex1GXOD2ceExqGnJMWaTWc6JzcFvMSV2hrRw
Xo7CmQERzr9nPp+V5b27owOi74TgLltzn1Hllb7fJALvaCZWhTSnDduDMvcU/bxt/OUyvOeNfpMs
B/2eQMD9+Esbo8jjY5LXYu+zKUwrCs74FIbPI9EozfrCP0EuK/HGa/ui5ToVj6BN+0uUdMtza6Sm
IW9wbUa9r8VZhxIL3q/KJta8STKLYkNU/zWk1iYczdEdcEPosHLg4Vr9Q2eGpKHJbqK2oucmC/LU
Hc11d9pMNHyDWCz6bQqnNbNHucGdy5Q584Ppk4IvfEhvMqxNKeOqRSlXhr/0GGmUDOnNxM5l6Si1
9hn8XLNpo0kBqVtVqAoBJpQB0/T0yTKMEvNeWERMTpen4IJda/ws5q9BsOGIxlfs+Rb2y+xEfvhn
BFvVaccVGLZsFz5T5oCOq6KJK+3dwEk70nFXmpW696Y90R0nnZONPRWs1tLkwV3iP3YpztNlIyv6
IRLYL6zQ/3MUt4gNWYZ6WOzX3knno5RmBi1qA3rlKwBrMzfF8SjPKrAvr5o1nCFFZ87f5EzfHn2Z
dstp9lguBHOPByQjeTSN0t7tU+Hf7XNY4tdXzHkfLGSVKx42nMyKwHZlY8/iDuAuIul1Atyo8GWh
UQYmDZ88FgPXN+iQ/YpbUyinnMyCuXeVAOALNn9WHIrPLdzIMV4DkBTs4FoibIZbkS/1D5Ww92u+
Mt9SeLt8bwxEt4pdQmezeBpdgjUAJwA3yWSxHfpuYKXrYauYcM+2akJT+NEP10NpWxzDWPPRnZUJ
XDSqaZgRv2MFIS9lqsnIhda3S9SWQzFvVpZiM+gyN2QmVXe7ptEufCDp9fsZ/Y+nSEK5wlzJ7ZtI
+D8D4sbDShQNscuso2uOuX8ovUYqoueI2fTBzDc8U5bncqYOMwbSYWkg6oelV8b3gqbBXS5RQs/o
RdAhAygEvn5UwxNrD0WAFdaOuLlLtLo8RuEDuCPfLHuPO+2DozXRhr+fNNxrWrm6TQxCgehdUftk
wFb1vgaQL3UX04i7ikE016UdhXrx/wHEAVVrKlXu55N72zh0gHCrq/bJFW6lqHE5ODa5dq69aEEv
lajPi8A4vXELs7JNf9pLqe51JQUOHDRAlNMV+OACviBegVRmVNmY2n/rUR7aA9UlFPXRirl+o3JQ
8KT86JOWLYtEIhjs5I4AsXT4hDykLslgC3VvdZr1/Rzu0/Wid2A3C/Sm48xuUTpuzpOHyW0ATnW2
e6HsRC840HFsTdM1umEiQWsi3/lZl70sTzHYKh8IQzbEVDDz/zIczcQ19IjeKUGwlS+eDS7bye8k
bEgm9sI/x+OsAkjsIWBACQiIFM03YG78YkGOUk+ePtqXLSt/u+JYkApmX3zPrpYrj8xyHjH9iwxq
ykSjTjQAbiyX15z31dROfJ4VKEGpafKALKZZXYiaHd6w1ox7HpnprSDnx0gqjFYGKs1MWZKCwXIC
hKO09dc+ALcDzjSvCsZXZgLXCDeCTihnC2U/WsN8eV3USv2IViKpPyKLnZy0kQzIwh/Wu26bhA2r
UndSnb7Qzstab+ZPn4P+kHOnAXsBY1OyUxfZylHqRnmYUD2uKQ4CxK04mgpdoo7zar0CJ4ZeBOS6
sAy0D5eEYeZesQHHSixUi94KKdgsA5tEf4qKufhEM2iVH+6WYjf9t3YH99Tj8Gc0vMTCEoo9dEgT
h5DO9gjMxEf4SvBSyHWpUxTg0AIeWZK/fmzbjZVgsJHIVrApVfEyHMAZSZSlMHjC5ck886bTWB/4
0Ks0RoaIHXaXUGf4ZvsdM1usTg8mY8P1IkxMt7C3WrOYVJIWBt9Kmqd8RVUq0zn96+zL+9Gr//1e
uRkQEUC2JACQxzzW6M46jz6utMWZH+rOSTI3Wa5gN3FXe8MdqXme+w48LfatwdhDVFsLKoYW6qns
9NvbJGlLvlSw6BeSJndHKJWMzM51QPkrv7mz7KO8eiBn0mXiwGdWU0XmKArXrUMhmDOVvIPRLqDx
5Cu0NrhuENQFNOBIHPAtBYvfQx47jq1cNwwyZfUSVdbkAKlzP764QDlTzg7FRE4bgJ7NhJ+X/H7i
f9fNfQnbwPcE7rRUABdo2Zr9RCPBR2olC6TfmEuI3AXbPNeR4AW73XBNBaQVq7U5C6jkr3oAl4H7
rGKcV9UvT0g2nDkScEtfeG2SHL4BkGoKwo7K3nCu9j0i63SvuljMmZxRMRActLeea9xNIgMZGTT9
RyfXVlgLhvfofzLoBxQqF+t7XJqa6oDloDQSlqezrEAAfcC1nD+feufxXOPZpaBAJzVi82jyxFdW
ss5wbCy932rhF8f7XahIVVPxVcfQ3GCIs4d+20p4UG6pAdBbbnFU+kN1iVsLe3Mrmf4h8a502Vs9
UC124O4ysg+fcxRsVQxdGh12qYyUlPKsvGHC/k+ZeHEsVlvWpdETAboWIv5n+585Yx9jFnCZVsV4
a9B+jglS/DdnZhu550sinXs/Q/o+IaWPiukX97/hNr4U/s7ygXtc9YVNm+DF6m250nJuCbQCm9Lg
v1zVzCHFZA5H84EFtDtRfFYmbEw+8ye0j9woaeiaFXXQEdZ+pInWbHT6I3nULGEBWjhp+naDZRjz
CkZN6qpAOuKv8Nk7CrZ1uHaDFlYyep3tHdd/q8tUpn75JvcY8swVU4WKClgPDCqsxt2k4zeLArFW
xcv0/g1FIBlJ8YJoF6jBdlax8pCs7PA31c8wVKiwEap1iXPPt1KNsHZdpwyKlJHDn6qWerYz52ch
vIqcQ0iO/R0CSpYS5dBINLYMmDt58v/jZz9uI09zAhbjkGF9bC5zbzGlqLY6R1uVbsXKCs0fdSWH
r8NRHF7nt9cRA6mKUYfYCeWRCVegAQpmG13HiH6L2JqDmu6X5TiZLUsPD8vcShS7RRerfgFn5qZm
7u2eQFAZtRSrsZZnTJFEdVDkcYMXngtE/bwgd3msAO5Tjgv/fvBNBQg0oQMjUDdoZADzQUYehbEO
GyyAtpKwnC5uWbbYE/d4xq8xJ3IwUblxWWrNT/WYjtI6QzF6FSwSDRlEqt1WIj3yeG0aksm/qWL9
u3HI2WzYDwh8CqGOBE2BPGFHooADgaLDbZ2ZE5lu6lgeRu/NdGtPtsw6gcLrTweo8YsQB7l2kAKZ
tnErsO2wTrNoNYhXcjkgsI/X0u1Nn/Vgl4/oBCEjwrSjgLa6ejJZ2GHZ9IeohXDYMJVKgL9kT4Z6
p3Htyg8vadNXSjojNB5Zx3wOcMY+Q3/M6g+K3nsZ73HJs4NgFwRacoAjXxZO6wNYJSY2lqnmzbnL
22k/jcgkisj1jMhq4D5YYIC+r+uEgDbMJy0feWhaiG3SwAOuttpSds+QqU+ZOcaxsVRpjoSIXytV
tjeBaQP2vsbxYsupxzl7/l/x85gtgXIO8N+p1kT3/NAK32fuW7C6FkJhakNdHbRLcG9BSEogZcp/
CkdQYojekvh6es4OynANUZHqD3dIxWCigsRrQw+tySpQ4JFin97bGgVHoKeNgXwzLJwY6/lBgJSD
pKS+73i8er7WA0BC0XPNgnxpLkMwUcfQrBWQ0vfNBNDbLiYLb3/uIb91hMatpH1YTgCeoTMAVBOP
kt4A3bDU5p8PiYInYU6KSmaPWsM6S8N3n2cT8ACnCv8YzK0k4aEnBIlMGDGtBwgTRqNe/fUGHz5D
J67t886l021dr8UxT3qlPREHjFo5vLIAkeBdc6mpCgyZdZ/AojIDY2xuxq62q64w8fqumvCn7FbG
ld+PgPRDjW4ehuvQAdQ/IsUHiUsUZ35y0ZXoFkI9mzkZ8EphBtRCcMaFQ3iCcpdd6qT6pAH7ytVl
sKpSC4WN3xrnLwZxM/T2YXh97T0CYhOomJn4wyZ4ILiuybuuA2yLBeyYTx3iHrgzLDyuusRfpqSy
0RVw00qR7SXH2NtRpuJG4XhuB27ukdj+aB0CvPydytzjCx28Bdu15Ke/YJpl9fOODlbMqIAHTAE1
lY48iS8+eD+7wcWB2/YvnVo00oD+qCcjkM6NsTODfHIoUkAV9u9uvDPwKMUjf8RFxwsqCOZ+ohvG
WRmBnNVgn10Tnn/vQo6O9tCyoCw+LtPQmNtD7W5ncVn2dXJamBmnUnbN0+xWkI64h8/OxeAWIW/n
0hRf9udAXMNoF31QQEBleCF0Ln+OuEHFylS3K4URyWEUbWwMvBtKsi1xXSzGVqAENE1sDMj/ARL6
+IofYXZNxcRwLqdaOq0kLUjHO2CUEBeAmYK4/crxv/KWoDIBEFWHTweVSugM1xRe6Ckt0ShLehYq
/4lQGr9GjxsMv8BIESyBJc2y34GLgSbUjfswqyf5KSjCZYtyM2INSQtbBscCQsGhADiU6noOOI2w
iBvwQlI013ar61SD1I8q3Pbl33qo6FEyh72ll1cX/heGsFhkEhUGYPC8F+Mh7RE/IWeCXQI1NUlw
zofxsvyjFFOlc3qoY7++CnXj5ejYp9bGCJyqz+upM03kJvyM4nN4CxcJjPt+aYX0/b9K6waLqcId
2tSFTmg1JVhs3TVlA+txz1DdQqSkZCjSn+BsVbBCwUI20NvBN4hTPKL395EVy9Rd4zwXg8JRbwJ6
vgsI3WBtXX200Aew/jehl4R4nD2oYXM9+r11DFFBMqktZaC/kI5svNPqYxxXukOS99QlTuIAIxBM
gfuo/54Mg6xr3LW7Reui/MyaSaPEimrzmo97Br0S7DRf5zruQbiI/OTSrNZO7nGGyXHdx534mhjp
kYqOLuWahqRmbhxDWphwZ6AoSuNVbMPxwKmtR6Dbsn3XNXMRAZFFZzar7kPA8SRa6P6MNG64+ARU
WMAeRuap8ZaRSQcB0dfUPWSYN4x6gt2f0ho/DUoWB3t67XI4kP73nQjUxPNCwM1rSuWGQ9t1iLLR
9IvgJ2gYwrC2MjlS9+mN8jZKCi4NaZ+8hq8vTdY0iwWa2n1kWAdDRoB/Hzpn/AApCytJKRg/AWBW
baJXUpsH0gE+kAacgeIHaNIBV6IjHYFXk50b++DpM0xsQzSsfwH1KFgHNSNQAiH8SQpfAfpwRMdF
rIS7AnJ+hlTvDfiUaroHJm/fPLX9FhSXGmWclXbB7ceXt/J9rlw1WEN9foCWDeECtBXuUgwEg/cd
koLliw0cIFTBmXJwH56QPHRdTzlfINq/TPAbWij7vWgitrGvXy2DOfaEGrl9IUB4UaXUQzVbBbvs
5WRCLj6Hxrfw+3syq5L9oP/lyZ+3srfpqnUArzwnWgXkRvtl/tzku/qjO49v0kEWOvFKskjCyq20
FwTduVSktToUUO29MugRgPQzNPi3L3cOY3GQeTmQlspvOw0FYK05hOxMzaHJ4riUlpUtXMps7IwA
y9o7krW3/HinrMR8rJuj9cOS/4hnMOVJm7R/S4rqQJNgFAd5oV0iyfe9EbvEv6DDzAEx5VDyJbSn
qyNRT0w7+jBW1HEPct5Htg/d632CF3fTzQJTL4kPBW0tf+Me8Q7ft3GrW9wyi5PjD8gaoTS/+kFq
LyTbaYS9px4RzPDYKN92IHhaI476UDiteTOejFZoYeRzNb4B+LGTpyz/p+vZsqmprKUEQR9oTtlM
G15bjJV9/P/Z47r0/sEyCX8LJzHFunst8944sAuwIWuTO/s1ysvE4Fz7tYQ7Jq1lgQAb2itIstPj
ehzY0Lhka8GFLcU7ZJN2GDzuvWEGIiCmHuctSSGCh/eKq6xGfyJSlL7MwN5MkXt+ar7C1A/bXNGd
7oN/AHfUDaXoTRbx4p6+rIhRceIaj4ep32/AyV8WyZf4W/MSIvussBPfabntr+pjYuzsQjYqIZHs
om3cRmyXdHUB0pmmgRlnUNb90dY5vj17d0mXfRq2BwTJXqK8Le32+avIoe8v9SIRbg+9SMKj8Scl
w65F8IDEJV6m4cpZ4DtFXXshnEzLb1nJzRr8BJQy36N8zsoxtk9FMlG/deU28uWHHt0q5X1bHzYL
n+KUoYF6+pAnviD7DHWwIpEEYvQAkxwvMcWZlMP+xsUCqC05ROYZZVua9dlnpvHAmmWXMLxpKu1G
uY7qoKf+zJDco4exx14lnNMsKgoawP4jIzG3dYC72fKZ2xr7cQWz8FkZQDZbmnu9xcq6qBpID8Ux
pmfNlGyN9iztM/HALo/qomMJ1pmfx0qWbKTYOTk9qejmJzGp2Yq7h6zJPL+Zuj8rDCDePuUUipBZ
mzOV2CbaKc1uFsYinNqOq+jclLz/bQvTLPK03KTADyqn70RbTYsCEfEN9LYeAdYfWA35QEJbTCGV
PyyNVhuAxpjFaR9UKYbY2SGhhVNNVNhB/wac4QucDdqrGyL5kWBcJ56eajQuNihEaOAljXzkdwz1
uf/C2qkj3z53LLn0IVnrncVbboYFdRuP2/73WKkYLmzq+YG0TqGk4ILSQurihxIXa47a15DX5FM9
HYIl5eJifn/m1jVv+i+mQos2C66ucnDRObbfPsvPN1gebJOUOkPLCtWWN+PNvcWBJGLyqzO72vwA
Z/1FULRE7uYgZvLPtZNIJhxFFLab8SCT3AgmJjv9kxgTC3XeMUkvNgPnZX7JWZh4I4pgqnRythFr
nGOTT+XzLy3473gWATENEs0AOFpj4C4svJDCvpYObaz4COtGp8xWLAfq9qTEfhCbcrfomQrgts1A
T5ND3PhwTIGhw6iZpMZV21J9vYyQit9zQFE5+zV9ztx2xfJsghP2WuO1B6xReBTReTsZ8T2cHHF2
TkbO6KSFfZSPVoScY13YEZbg7wLwUe2AfU/9/i0CaLK4lGZiRfj+WKpqDBissmVm5v+NRLjKovmd
qfcR3CTfrZVRffpdQ3MeANreLAUxOK6UDurSUdphng/rpSc3TPWXNNlXtxeYygOj95Y47bsBtCcx
S+VqFM/tSggtjrKj/sXtQIVov/DjQKeMqHtSBFuWHv8EzC/Wu31VzAzqMHvtqJyr2noyWN1mH+I2
yLdbzyc06++1DiYS6FPXgu7AckUS/VHjgLlLD/Kho0PV6JLyIFQffqaDFLui0d5MjU8BkBXxjhx8
lh5XHqpDOpQvM4uo8LG7RSflhbi0SksT67/6NwMMWHKXVv99t7FhLgMWIcUMpv5ng0A/+nPkVxYH
GtafQ/BVvdzXnpXdnws2aaI+vglkGXEHvONyAAYGP+cElkHc9kTnsUdCME5qFD5VXFTPLYsW1F14
tNpBcfZIlHGv8/fm/6R2LnxLYcYSlJIJNYaoBRQG7hT8uJnZ5HLJ7Gg5fxYsPcbLnKVuMb4NLYcR
LV7b27hRBCF9rWQVI0C4KOuLxOB4MRFM1u8YI+fPMmyzrMZ/yo1aJN7i9FXRO+lNsSNC3tDZUo+h
DJ/pPMc3FSJWKyXjv5ubNnvEHzp0X1OYdPBYUwofgtXZ4GVxLwXtPb18IJvUdc/CyAZj+J1BwtxY
ZPIyMOVReYo75dzP4wQGkTS2+8lvNGsnTFI8XmdamPuw5m+6VEjXUniSpD43YLwLg0pSlWI9PZMW
NzZ6nm2H1LRZTxgaugwJfHXoPN8m5CrTKjdfq8QQ5MSWz/Op3hZY0BrSQu17qbQ+IlGWuo/lVIwG
j+wrS5ZMpQLmsYbI1AKfsJndVzF4VOihMddwpxLq7lC14nVyJmDELq/4WWHSw02eqCsXTetwCGkw
QFHg+NmM9MTHsezrjg23vy65+9XmGoPp1O9aEy05CbT64amlogmxD5B5HbFKVTuwS9FpxgZue0BP
JJfslcQRwXNfUsk9uVOi7PJgk3sG+JeSz9BPCwrRQEaE3nxiIoNQ9rM50TFqv/MXqeqUG9qChuJH
94NpdqlKPWrOFgDhGNMXwz3nViPr9hIwfKNmdsE+e6BW/68p3GTtdcAvXs1NwSVJlPDgwrKy4xAA
d1fSfQ4wU0mYDKSsHL4WMGaPm4zWUw5dVXZ94HsE/LfNS2tSaV1rEHg2ERuY91C+ajkZpH1YbTWX
TXRMsa+kUc1vEalqSqRWNZI9hY9HpFOJDK60ApkSHbFRt+MkcsZFdyeH+ApEn+zyvPHL+KlnNd/r
LZRWr7FQ5xxkYS9A/yQ/hUQWLoQBJUBAsjA8/WMklV8VsoCCplF9kSCRqbbWPp96y6zR2UBw9kA4
I0ojvMbRi4hQBUhGNlmiHbybbDsPFwDtSPGkBU9rSYOQ+mKmGbildFkpeatCYGpeeQcjqNuE+KxK
uPPZj6Io/LAP4gzY26bufjs5E6pZ+2otfpEZJY2rLkj0i5Vk2G8glZ8w71xHbABsbyEuCvG7ZmRB
31EhXwaV2XXT5fFDxpG5iT97LOp+sju7oaDG7gO7Gl5kx/+hx0p22VZ+DomFyu/UsqlTFMHMwZ8v
s8ibUgNvnbeeNddwbClh03MDIH+AlmIjAdbSQp2LJ39RgNPM+1Xj/ivAmyU8WarV+YVSAe119y+X
ZxbWmwfGvUPUyVbeIfqMuTaETLzvplivKvr+H3psVulC9ULcYuCIxMe8s9QOFAYBVjHnmd18GwUm
cjuXtB+ITicZ26mkw5+iEKTio8Eex8B4L7mdyX7k74jkkYMnHutZujg03TZotEvkaZZggq88ZyeO
qCvJzpcHPlFXfwTFz2JxDO4hfyInUoZCXmgUVJEE9N3j7P8vUTfKOfgYcPhWuKQXoAkV0UK+AGSG
CABzqr98A8AJK/jPc5COoap/G1EdcAu4wGx2dk7mLpou2vd80v32ezw8nDk0osht0i8yag5uiFBJ
TohJ94qCvn4BZA02L+CU2Pe5rIdzwtfzE0iDte9tK68LQ9CLfyKnevX1XgA3GAW7dhGwvLAJeGDb
a4S2Y8w8kF++quxPuNhcRVkAxlIU58+Nb9mrhMnY9cFN6Yti+YxIObZzLayT+qe6joRdB2GBc2jL
rjjXAM3FvsFgYcx+QbxNTC7N9TPOr6yKMfQlYiikYdq//JlRg0qANJMFSa21Sp96wM9tA2pToFe0
Br14NKYoCts9FwB/E7HUns2wgkLSHg0uizuxL5wQ9Z7DMRIkg3iN+/BYnrMejm0T9EKd6VOBXFG5
+R/1klPdChR2h8eallk6ZfkHpnjoE0Hgsc0+qjwmZO9bZHztnbydlkoM7AyvrYdLHoC1RwgDVBmr
nrei5cvgFNfWzlPvJbI3JRoqrIK7rZpUG5JWDZlFcRH5pC6aMb2XaPfp1Qm1uNgqbTI9XnViq00O
2PN2j87pxSi33tBZOsZB7K+ZDlqpaRX7owwvz9biJBvYZR0dh8QEldoIK5Icb2W2cIkcl0kd4j3C
E57DI2qsKfk9AiIWTNbIbeilnN74Iz27lrOBU3gmIZn080YGUwO3MBxYw6E7J+2FTJK0WEvaX09A
JQKYx8DJgSDNvhZKTZOYQqTvvMPfKQvzdyguFMxxoLmuyf8X4csEaAM/V/Us1uVaAyoQGUQR4zyn
6CR/cc7so4L7oKqTGMvW3tRIAmImr4Mc66QApze11T/qJ2egtO5QxgitkavNAYpYuNX9ZJwrVaCl
glJaAhbjjkOjfl6p+8pOWdi81sH3grh+zt+SweDtRJR6AUMuPmppjE0PscNNj70ZOJ0cmQ9sMFn/
eBnlOIosSze9IQYX8xoehGKTqibvEUKBe2UHvZTqCrrhuket3F5u0MXTdQC0KBcgI9BM/r3zKfMp
BGzRRG9W7n1R+41MyX5J3EnSvY2SuZ/guSlNn7c9nWiIBFGIwBYnr2xf8cB9gn/8lhH3g1RMdwPM
jR/yDvJXlcjH0ME4CNy6GJbsYxCUwCnk23duzrlxhIGFzpPv77eAzC0l/qRCshn/Jzkft8KBqDGf
e+Ab+7yH7ol16arL/BG9DbqJBoXKGzj+0D22Yoz5jbBiiSCn/Rjun397ADaaLsLB/yNIkcxlsBrg
1ypDvndlB+kfj+goSxYTrkUkBw2LnQXgHqa6nnMcZ4HCE1hpjp8WGZAya8s3iUVZK7j2JC1DSdv0
zLtJIlOonnm1OwBMfdYji+ZMB/G4bt5wp/ma2T1/lpDj4fPEEA/qGIqkWwoynLl/nXkRk9ennt1g
medG6oq24nDpKaGqA0HVDJgtNogt/eIVTczPPGmWUihUsmBU5qP/f/UEQZoZ5mtCbUsgvuTGyvk0
VSX+WCGZOqKd2/xQUz1fVN0Wj8yZJKNOFYy/jMV5dWJ2/92KXDtFCInUYKCmTETNlukq+VHLgpNa
10MIrEIek60aLfjFJEbitUn9GnhIiJibEKgIWtKr7K+713kIYQhNiuhb5hRhPc2MgiAzheBfsLnt
+WMVxUAXHeuczOJ1DPr+Z3uHmTmwiJ5lIza8JlAWD39Ne2sjOpeXHO+K87J0ldhv55203NYQUqOq
duGtf85jA84NUCGtYD7MaS8XmTlionkADFJ2QFZGL2zSdUxz9zIyrYSAai8Sd6fHG3R0zP6P5BMo
CmzyqIz5z3qXkZGol2hs5nP3FKSamMYTZcRX8ehllH+lSS4jhtAT2NJnXOC/lcMpMuxllLQWaFqs
yhe9ch3lnUlqlMP9h5RZyWWT4t4RJgICj46TwbVdXY/Qa6l0XaPaQjunFxiaadWI2BDUQbaWuBJ2
XdRuzmzmzK51qHsJipeo3hZnf/KYtdxRG1Xp1+jko2Ld5563tdE2dQpXVYaqjOlVqm5q+nYyPRle
kCbcm0Tumnk+VC5psmwfdiyTmurogAaw0ciRVP2+niYmBg/W0Z3ZHpLDTpyVIlt16GVw0HebMa4h
9IZJ60TMeuTH9oeo5Vu8yU2Ayy7Q4W0N+/95HOYbr/yc4LNzw+DcsZh9A0W/WI/Zs/IRrr43p6tV
aEG3dTfOk7CoJ65f96HFU6Iz7QdKbZK0js0cZMgN0S2UnmDYOciNASDIgfGJy78lNJ1S3miSySg3
077RGLGnTun9TZ9Dy0FBfni8aPoWLMXtl9bgyjhrjA1YcFuUJvs3atzOPaF/7DeWZjj3ayGjmOGl
FvxS7Mhp6gXFv4P2gJwniZr09IQPYQjnjgHPeWU7mnVxyAObCI4JU4hbwN1wkbRZheofO8KbjUBF
LZYnD6kGvjQzaApYnfLze8relYHmY+x6tBQghxmBaTscjzF/Lsak8I8JZmh2bLQPQEdh1xLKNRDh
+SEzVn8toKtKwi3vxFomxjzHVKYvfFngvvQ606dg854e+vBXNVAOEP0Ab8HUzyVrolUrzchKnjNd
G2KoTu2GbOl28wmnPGq9yQJmZM7gJi/K/TW8IgX6jebuFx5Id4Mc08IeQcdUUJ+irv+V921jqdLS
I6u5ZUmn1LMetfhywKCPdjEkEDVaTj3x4WnLm96Hw+oxQ2feSQ9KRXI9JEd/ZXZT99jFJe4HXXgp
vnmeoyAUVwHjm4EGSVg982c1xj+EpihXxLLok0Q8VseoojAVwoC+TYriJAAdcZj2UMn0++FU2b1i
T3V5UVnSwlGqEQIoFVDr7pxh91w6AtkMQcJ8PIKai3yV7CHgoqo218xf+6KDmFNJZY3WGtdszxdk
54xD57HZEUzF2E+ETouxYq0RtqQcGGrEE7qB2aXyiHglPwzJmXCOf6KN/cZfIiyzvzhJLbjXsHK7
WfJIFUxd6c3xEA+UjqLJtlq87m407HhURWXX0ergjpickF8psV7AzZl2g7VHHCePwjtz0VW0Q/u2
TlA5rIhiZ+O7f5T1t4zVTUG54TLewXkmtkxJ4fxa1ze5nDlJtrD+7WG83BglLX69/CgPgqE5uJp1
jEkL33eIMlIWktam5wCRAedumityh9bIgeBZfKl0Hxa2yM6pah+K+eoUJBhc6n8loBQWIB9VHr1k
y6DqDpmQhrk3fBXd/QBp42fxC+ndV0j9zqNSKxs5Le+Gzc+P9FFrfGqCUVUTKpYb0KrEN+D0/SsS
NFufcqp354lng6J3tuC4jKUphyIm9cUz3XgyK2c/D+VKjIHHYbfW6Mstr45paMPJ9M/k/LZ4+H/s
OrvIGllEWsp5fIYzfFTXzdGiHcIt6KjOMItubjdIGGX9MNAJ6thSRHKpTCJdj+u3iF/k2flmKs/4
kSbcVKXPUtL/TJPATEFheVluDkIjcOPvDZKzG4Aeokxh5DIWEWjuW7+UoozM2XPMyEF+s/8pf/mT
bVwQxJyshtS1dybPt2htkBBImo8qxx+AwwjgHnhOp90uvirD93vUHIOgIh3H6L7IzOpnzxXK0+i4
e9uxNeURKwwu0Nfgx0ReW202ifv+QFDdpmg1MevfvoWrN1AjJYwQCE+70FK+FClBJscWQHY1/MVV
NtALU2jrryG+qUHI1wfohuHjOOqLTUj33Ity4YK0rYPl+wMjgr8yCIr0VPE2KwH4E/KGlLbMjLH7
nW20z8Ac5sDV2s+zZARTt1U7ThioroSf5GvfzhF4z9hggvI3sTVjk9R1EVuy4X7QHUELVVE4gwFx
8QvYWUfVRgn57SGDXMQrKpOuK/FuS51GXML0d2VenVlOHJM9ZjqX1H2nA1RKqZrfFxWtgdxSD72r
UkMY7vVDKteB+uCOEhgJOEndng2Ge+OJYVUNDORstRgtGHUuYY2SlUYiHkw/c6Et4E6l1Xtlf7jW
rfrb9ftaADPju3W8NYy9ZStJIg5M8hSUbAaYqPUxkgTg2B4wX75KndjTxc+jGfTbmHNzH2jvdkPV
mgHqSKaZK5cswyPY4ScIBXrgeSuQh1OHVhs4/A6INfIeYjAQVfi1QIEfSeFRU+8uGLzX/BXvNBp1
F6c1g8oG8K2Q5TE4taoodFkGDeBlmAurJWOCsD3f12yYJ3r5ye9MwY9AH2BaE5YMW3Rap5khbwjm
adVOQ08FbeXlYLqpB9nbgf9nSSq9+EuXK7rwoaX1BGeiQjy/nNc1bnQRwBPp7x4KBHOJlbUx2z+W
0A/J7t3pmvjz5XYrUUBhORkyufxUECqrUOjk2EUon99lAry+Uzpr9LmM5zlML9SiyZs69TfSTT3o
TbMNwAYfvzkaEfCqeYVnIJN3TBSkGRdmf94gr1q0F1izlu7kqqc0MKHQG7l6QKxvDB4cpwiL2PQY
S3Br3QYJuUDxM3nytVsJeiXmqCv7Nks3yOjFXYxtOcprDnFurYwzHxytJPPU90BmSCPyaF4pbTiI
/wmf7J+hR9yTSaFgy67xJoj24g7LdMvx8MqeDqbXFq0Sn003CrvDCfqZZIP4r8Jb8pfIPtRfboOW
6LHcjbJ5YsxXdIs1/FwzBqL4Frzh34FbiDz4SZ/IoE1x5QGCF6M+2hwxSQCwJh7zoGwsixwaaVOK
pK8y6x5vaW05B0nQTg09INRSRoToBHIlLoB18kBEykBM4PJoACp75t7AmC73lXd0XqA6iETmgRPm
/eyaTERbstvvDGVr6BANulSQCum3XO8J0ElhXaByM8+K09vFHuO3u02MdKM4b7Y0gCmXY0eUuprK
Elog4YAitTWFT8QEtgQbEXLHf+kCe2oLxrmz85Zrr7C0Sj2r7QV8PZmFfg01wXRtovveoUatUJv8
FqaRQZqlQPUJ0UCPB5pI+OIGZOTReuWcEXUt8KXcF/6ShFqSw7mT24/I1tUPU8ttjln62FwFIrBT
x1wHmvXvkOANZ5P8awLNRD9iRyOquUB80Vuhas1oCULGQxBuCQW49R7xNSsoDccSGVvC+zKaNG+K
QMuqs60rQWDXzFtNqUB7cbKJ134mUeTPgE/TYC/czZX7xI1GEcqlWq9BBCe2KMIWe/nvMVsw4aUP
/17s18ldbn4E1KIsXAppoSYRiDZxow+MrNg0/8MBJwf2q81LdWs6RwNS4wis99UizjHxfBN1NRWL
Y/MSMIvDBGvmcSRAeyNYZyAeNzBHCWug548F2g8K7ur/+PVJWvHsa+bSS6X3dI9XVqvnCTXvuQ7I
Hy3i+ULXCVV3siH14GItoaicR40OFO595lhgkRlXE25RxCLm61/VkB1LVtB/VPgrhydK2y1+OFM8
AWYkxwPBA73iyswN/QiL2gM+LraOoalF4Ne8GJrqldeKxgsea7Od+syEeEB61+ecUQ/M88XzrXDu
9MlMqo1PLsb3mMzJCfIVoRrYoS6TrIs19Ch+BdoGquDVSmRxCHKk0jmp99AfefKgb2dsyXxvtjFG
HUkTCFXy5jSS79kJm1mV2yjwbiD8qRufy4FP/01Wj6PJRVuO9O42RdjCWwNYgNWyWxML1XxTpZQG
A1+5bde3JGLgMnHH7rHi9fVYIGIe1zXYFjh5cTyKZRutOAxlsi+0yqbm6JZq8EVTRkNyHJs2Dtz0
DnRd24QZArilDSftsgO/27hOjStpKVfCg5yrK3yHJ4S0SAj2ErCGOYGgR5FVCuUw4EHIZvYQAZ6I
O3gt10jjYRzbTLSJy2HXdqGgWEQUlOs4Gpasej9PINOZhgF++atKnvKd+/xEVEyINz/KpPdRHrIG
JaMpL3nvUlpUbyj4UpQth0Mb9rwI3My1HeZUdMnN4dUuP5/Fq4/p3x8d1zhNQvKh5MNAE6au5nRM
IJ4MOcqEsxcetLLNjvQ1GdAzsrDeyKlquJdyYjxGWi5y6ddNI3XenJpJ754/q6wON+CVnXqGQmYl
LBCqmu/cRZeyNRN3zqUwGGMYIyrD/uIyoemPH9p/+erlE/s5KhMtcU0n/+zwStc1ivejq5GJySF7
ZqpCRZ5SigZZsfhTGLGmzZ14jqC36ugfAGXcaarh+RPRiuc240oHVZHrEq+kBLCym9dLoGyjrzcA
jWDP5YQUQ9tw3Rbs72R4etdqzT+2GeBDr2113c3kiIyeUS4WtE4hpvGiSAciD3O3xpTYQD/uF721
sWMHfoj1yR0UhHGDsoGPunuLlQrbwy0BDKyv+m8APSu47qVDL8QBHhg9Fnanws8J5LDCTas8V7Dq
WC4xLiSJGn3Q0UUivDVuf/Hi/SSE5C3v705ajDESK7mRkXfZmy6Sm8KNPIusceHUNuMaRUocBiaP
nu2E7ukpfz+YGPQgYP9O6lWl1Q6ALNxmMX9YPa5DbyIAwQOJxHmVvw9bAX7lu1KtqNXSrYsqTwfO
M53xJ7j4fFCfdUdpk8S3eI89zFo6tIbF/1elWNBscOWM9EXLanIMTZO4CKLdVvUTrHbA7zhFoqrv
bdVncd5aeeBdKY3gw5KSJU5um9jbUNysxMco1jToePQgULtLXG+HUh2TRe3zhct4SYAGnymWyZXC
rc0c0IsTK6eqyIgNDta+o7noe1BUPS42fxOf+xnRIVcRLW3eCr8wi1Vf7uYeed80IixUs8tjRbt5
5TH28CbMm6/eLmJUEbkOWGiq/YVdPfjbuPoc6ndFp5iDh8ptmORWAafBzGb47dJqjE92Of0cE4wt
DP6Oh8NkcLaoi3hFNze00+NLiaun+jDg/jhgSz0GJhsisSPILcTsBnHuMO1jFl+WMKOQWHLFDmtP
ZyGZOKxmNQ3RTZ+B3VJ+q4rnEC9Z4kguCVeaKq4f4BBMWVeANCohM8Z7kRcU7FOMtbeRzEZsozDF
zIRt14ud7ZhrjlRe5nPMhUyIecWTGwKJ1CqGf57nSCXxll9MhvIFDWelwTVSdxjJiT/FI6077jaL
kzs/9oOAlvoQcYZP222NxAZdjA05AjYVbPaNnvpF5wfbI0ifKP1XhBRoyD67Ym+wJdYoyrGQOfzz
yociEYLpD5N/Fhvyk9kD8lLAlxqMXiprT5elPoDeDtDk7duigy2v2G+4tlFcUxBw0QIg1NCymQvN
qYGwfgu9xctyABDyTrG5FlKrp0CBdDL0h1j2DqXaRKFPcMEHDN89c6CA4P2RjFv+MpSHI/pYnhlT
bH3N0dt+3Pm0aYk69+91KZojZn/JiULviTpQof7TQm8f+prrF1MVDNRXDEy6aXPQDLxG64l/7vUu
qhzSzLIjNRQr3a0SrGgbqpRhFwTND5FHIBGZNOZjiGV+P5tSq2UTj9q7esyBoY22fzT8DEPqWU7p
g0TCbbSxJ2pfQ5jcG+/v9T5eeSwFcPR1B4v3xLWJ6p6WddPvCRN9krKXZl8eBdqLgmob0N9AfZSr
7hZ8HOCFCBq0tjBA8qbYNkH+Eg48YayWKcDSnSB19GAZoD0bMHPqLoVCbp1Caud+2nTT47nt0fB2
hNdYcDaR4HODozwMkeVHbQq0S9Cm5Q2iQRRduV2lRKcun8xLexA8h0/RS63LIHXN8OTa4T+yATGt
2wYGnwPafs8wTMNS196KhmUGTmdup21C8+BWkX0Crpz1r9W+aru46zMajuJNYQgGUw9QT/RWKkQN
5qpKAj83h7oua0UC4puno1csvYxWjZ76Wo0VRsDT6mo0H3fczHOEBelCsfbvSuxTi0/2Mr1e5gL6
jEChDMXnEv83eaZ/7kQejQRXfRd2qsX9Ye2gUCuzBk2L3fwzJyEa1LeQMnWvehKglO1PFgRfQNyN
MGJsKYbwYzvKBBiOMg2HBn14drIlD8XgDAFQNSAkqFkoFmKhA7+0TIkxM+TC0xLIFCHVg0PN2prA
9VGg/v/d6afCZwhOZPi2u7HWdgUZg/hC0Ce9VRTNolobdSe06EFXx8v+GSgtNSaauiHMfLr7fS2H
vaH5huB8FvpwRh2roLwNZQCALDIcO8NVco/r7+cM7G6n9jC8IKlly7pzyBnGGEk0X6kN8xxeNezb
WeAjQKJwSjoGPzpyul29hMB4l0AiYRK3p9DojsIlSjfbXrXrIc9NhtllM9ZjTc/CPjhpKWM13QPT
9uWxb94NNXFfNE8L2jJ0zGnxunJYFHCtjkAWWGBUl/X4Q/qChy01l2sOzZGntsDw1Pp0QF37ircb
0hnKbH5Gb2m/JOXb1a9LKuhvZlo2C3W1ZL1LlIse9Q6Lc1q93mOyWQeBad+k17y/vfs40LSmfCDn
0GehePJzAqKQC0xHFYCsuYmBVflqY7GA9To+WP3M3gij13mgEoq8QYNlmjGZ5Hf5+3OuV92ZlP+g
PHVZfIULocK1J67tHQNTgHNiA1DmJrcbpQtSiYSv+U1jTytYPivjUff3g9egMComx0Peiji8fiD6
dgV4aaUL05fO+o7BnftHnrCDqwO79o8v4keKj0vAgzOjpCsS/7cA4sh/FebWrvhEklaLkMS3U0l2
qL1go3i9pDn3I4CYVbffQ9nRWuenbdFHgt27HDrEATIkaoUt/oB+KQrVbEGYHXQPVA3U62ESpR3A
WUdjkif952c4APwxYst+vKkqHNLnEbphC/vsQW8fz4QR7LI2P0+Apw/Q/lFi7a0I6BkwLJ/nGna0
6ne63AOvzVslwEs1bycAX0kWnTDScHVJj96TI1/WHzACLTtuvtz9QoSFWRM/jFFzUeSen1SNgH6d
eY7/HKdAu64CasSc7At2kNdOntHkfMYELxFJXQZpJg4D9q5Rru5SdQB+g0lPaywirCCZWdn+IeNX
J2tWmS3yXzY13FGb2saJka1xPqgcH7em3QADmlbNK8cynTSGa0bs7CCMxCN2ldN88rV40hZZan2D
hiMXMAOg1unFx15tIic44DVg9+hNXLO34nyPf0B3BoRXtUdeZmmZ3PyJdQCSBJ8qe9XGetLnLVAX
9aS6PRxg2OyaTueo0qUq8TsBaKX0eK9aBLzQkSzBrw/Z6sKKm+ofiMbdXt19jgxnKpUhE31l+9BT
Mq0joRqgjNL0U8t7j95cPq94/6qInWYeZqEuJES59JGksYILq2SaoeuBFSXBfYt47cRNDI3BeW3G
nltGcyx5wcqqJe+Tcg7sghHdhoFR3tX3Qx661IDcwvOkWCnpcvG5QSssNMAKp1cQV7P0tfAaTZ6U
qp0G/Xo9E58jprW4Qwvby9v0xzfbKheLeN4zjr17sTM9xpOMX9ikY8ykwlUvZUhFDAaN6NSS8RL0
3jCerWsbSPyybcTDfyYI0pvZ3fUzBUvokZv8sUxmWslCBC3ZfQyWK/UZ8lPftRpOVWsmD5xjGywK
dVdLOr1UE/d/uK/X19DWPHZWWqfvO2dH4d2zwnyBIW3PdlIyreKnYHF6/L01jDqMZZjGWbDGYDJW
KmUYuSOqd/GJGBK5YgEUZSkHeJSqnqFh74H5UHy615bl2q+1x3PZwyWopAN66wBFkxTmOqQy4TjZ
XokIv+vgrouiG1wPMvsIPSxuf1FP5PsA/4qp+AbMiw6vSu+Yx/2xB5TVzc12D7K7ocmYE7VIrMwm
F1nx0viAtP2f/YqfansAzE7/f2YMY1HipgK5Bkq0jq56oiaD9if0RU4Mzwu+ksRZNc2iTQQJLg/I
oYgXKNhbnJymZbAp+x9pSW2zMpJAaCkKEcxv2PWixNV5br952zq24ygtGvK9wsvZIQzszNnX2+bL
yH0SAxe7d54k/+3H+vHW4ujeaiJJ0kVcu11wiPx09UMPLgCT3PDis+5g0aQqIX6NTiB1VhRFCPnx
TVlKgn+qdMLUmFTP4M6bG0V2ECyjx5ydbSxc/8ZjvlmGyb9lE6pIpzQPGNtsZiYjnLcHWSzjR4Oe
b/cRcUjiFaoyrC11fz8RB4HLYNdiFthTHJ7EuSo0gJT6KlUHSwpJBospTpst7U/MWt4tVCsOrNgj
DzTvu5iRwtxPIzJG3cz1v655AXEZVqHU03RlVvyDb7zNV6TEc2V0fNdqPsmsm5UcokHbORIAYSvY
bvs2plYcddTYxu1kKQ8YFq8/dMyvzV36golOEgqZQtxuMWd2or8T89ZnXMYuUnwzfHSOlnr7wSKz
oZv8F7PVUH0AmDgc5MnFyAHRwhDioBcPLX9QEeW3aCkPxymUG/v0ba1xuKPqBTM6vLgUmh/QiOZl
vgkDxG2xw78TyWbcleKKIO/O1EY+ARGiyYzBhg52uFZ6q7rbkfkjFgQFBx8+1NxSHl49gg/18dJG
XKzQjkZRg3xhKlX19ZRRwcKSov8lFp1XaF844Q/5gqO6k23mPZA/0mf9IPvdgwL6Xejt7DyLCUYB
xW6XwRYqGexoTSgdna+IsB+U3IAotBKzVMb/RRFEQ0wt531ycQ+Ws2vN7fvsnJMfFlxmBLnaqRyN
4XzhsDwkVRSiKPSC9hL4pR7BLHOf2l9ucehHa6MXoENELGt9ufr/TsEGflCaOgQIsE6ZZEbZ8Ous
LuI9/MrRw1OYH3QzFSwlPAkcKHfoZF6K6xOeE/wqRwOK4+U4HnEN/kynxWhNodv2dYgGEV5jcw3X
dE+0KUWhEEdwD8ptFlih9GQBudh+SqLxZ2Dpa9BOI/yEP+WuJJIBPoRI5vOLUksxIQcnGqAXeqIe
+Kc0OAUL+z7keVimiRBWuQ8Zgb50rHDBEGBuL1P0EiGBxF1xCfRqeMXjnXDqbd/vtf1PIrDPAuk5
JN0ftOvGRy05Pt12qm7GQY+WCbwodmkBdQBkDMxyq8SWlelwmP6qIp4fnHfVmCTzsf83j0mRw+B7
PLqSTQI79zSrgcAnmor/ku49k0of7SE//+7wWbRPCdE1W6Ajpobz3oEn0xaT8xTCBUj9DaKyxJES
RRyQITeTKUd5flnjuRjaxUMCPv+GTEtkz/kutxQxUgJjylVgTec9RnEa2eln1tuj1frOpxF8Q32F
qSrQkbPK+juQNGHCs1Kbw6zqzSPqBBBnGpUJ8GTMko3Y/J56Hhu1TTDJJ3Z9dc56BZ3oALlhw4KC
5e/D6r2bM1826Za9kmGro61OqPUc9TwshZLiVQfoF9eai8wiGHnVa6IsfQSG7yCxlEQCcbxlkaGE
j0rM7yolhInQqQmesEiVF233F/aexIfHz36E4bTVjgkSxj3kyZU0ES6y6Egk/SiAr1p0IXjSALTW
gjKXZ4IXk77NgxnkEd449zN1FpGLz92SVe/bdlhPwufi+ysq5Ab6lADOGFqh9OWEqSN7J+7W2eKg
TY0KqgAf6YoHQi9kKj8Y2ryZ6GTG73eRd/c4n4qwITIAYtJ8uKhhumqr9OZYIedSOsznhNhi/q1N
NatMTEsmk2z54WonIPmetxZ79V6hV3XWQNQUxeqUIEUP+1Bfwbmui630Y12hjTavQU/Fsnhiotrx
aSk+3WvZPgzhl4gLq9z/AgPPRaW9d8esBHx5XO31eXhXSbJ6q5OBOaN0xNgLGr6+Yw5oLyTe6EHe
41oohQlG+UD7mDNZ0efImHWbpod0L3o47kTmtAEUIyWpwMCMLJXOKuYMZfqXE51ZquEkMiwKCFwa
R3bqjLdrIMGYjJaqwmim2HnkPCsqhnhzzGv1ySmTR88m+Hkwm8Rrd5C7JNe7VI5y+FKWuUg6piSr
06awOUoFWvIQmNqVDFlcF+Bd3g1KYWAjveNArFrBWywrp2Uc1iSDJvJNEjiaVur+dTDddRP5lq/w
IkQPSh3ENIMYmFlxm1EIL64ngrf6AWfjR1oaZvhdhnE7gA1v3VAMw76phmwDZ+ch2lAjaT7g5IvO
xoG8KTy7Trv506sFlFbzcWeQxMhCXTFyzidPZH2dwmoDuAazRqHnkgTPuA2BC1SxZraDk2x8hZGa
9xnYXyH+ohmnmGiYjPqyqgJ/LmD84kSPRsZc2aKA9lmCo+ZHAklydXa420w4W+FDqGOrTzR3YAtr
zGQZlYmQ+qazHNIdctZFwbwlibbSdNEDy2H8Vw2DZ0pgmg0tZoZ6HqV+hhdZ84Qal3Dq2hCFdQPN
oxnbmHgz9dz5p0vo7H+ssJmenTZ3JW2vs0F4c4XvfHumGQEtK3mDJtCKoTL9qHEBkNEpYlnWaQWO
Jf9dYYHRR9oV6b9EgNGy59MF3Aqk5FBvpiCXPcBPzD1nfOi6Bqc0AyVP7PiV9JV307hgrlep82Hp
zixROpYagvgKc1cAf7wabjbP7JxOvUTsR2VRqycdk/q1nKMbS5RvKVNxc/cKFW2wm/Fazi1zAir0
GKcxGnlJ7+ikwkWujWZZ8zETRDaHrBldVqbiVckCCLDBamYMCiKNRJOHEzjyBRnIr0V3CYCiBKuO
t2CiaKseAS6J7OOoynIbp6YtOA4s5lRVSmjCi1xJ8/A31WPdQC/rrB+xo5TB7yfiZPsjlohsYdC6
Dn3fW9QLIWIvBMB2RExSXFiZdPBLczEj0uTUAC/LR9z2lSBjUQDVhIX1yuzeCDpGqM3CiVCFLDme
1lZhVrGufl6CuuCTNkuRV5YNyFcJVs37rrCHW/NQCLowBf8i/1RFexQIQLS03R+NpwLDs000dhH+
/nkdBIJm1Lo9k/fG5M/G9Rwn7WL+or3tIHmkHt6EUIGh1j1mA6yOoY1az+DoqMKyDxyP1DWBZuSl
eodRFjT6O7LxYP/e/vFz+/duJ1tpcQEE1fU2rMoII4CP9YdOCkd5ieXX/oTdJodLm9ZOe/wBYKG9
zJkddwRavVn03op0+5TgEPUSL7nEyeKjddEFz9nQJk0MZnXktFt+nBuzN/69rTkVNatdOWaIe4qf
nQgkDKBCQdtw3TNVsgUzMb0Ck1uvbmkPCFfFICYOgZXI9iYgCcJe1preGmpgHMF7STPAvlYIABiG
I89D81IdVbtWuPOf4SSusCRshRFg1e+a+rNCaFV0IE2omzcIt8haSyYv+lm9WPZq27iB682RKkUy
yaNPAJHmPFhVrJ6/a9bS1bm6/Xhnh5trMKDCiHBitAZ0/dqCIO20LwGjatGNJS9xuhNMXkQr+mYW
Xqp6m9fi09EwRM/yRSwOGuYeVYOS5Jqucq/25ad8exf0YnvBYi8LbKbZ+F5HUobacajpnsFGdUap
Ow1ffzx2j05NtnTYe4/w8gROcJFjOG53IyfkdAZJU0jzwHpDF6DNwORf+drYAbktR85wKKq0WQhh
G8vS0S+9PN3RSM5brwi0sNXaFzw3lWmOqzwl7TVi+GeD3EOX6aplbiXcJs1QgiPjSVz77AhhB426
q2Ed30ivJDSURYyozxEGnq37d8dVhR4XNtvsc828BzXJNQdieAcR6Fxu3MReZQ/BBbTj33W+45WH
Hv7n82NYVcprJkAxelJQyAVPs5OezKtvZs+2B/T/lwHee5Cz2VMtRuC1BM2lbAn+J8ZM7h0ZBr3v
j2FgYQ/WQf88dnmugkWSWKTr8s2giFkPuRWLEnq1A50EijTIqzS8o4N9L8IdBUzxjI9jKuwbrZtu
N67kMjU9dieCUf3TkePZZ0zLW+/nimA71gRK1kPFcxgVVvd+OPzIfMaBuN8klYxhG7woozb283c7
EHy7+dd7UzkUn6FyIPxIADjzhOHSPNrih41rM/5WjJSYLGA2enJKNpEu50CikTx2eoRfQuY40y0o
r9fifKtuy+dH9QdJ4laLGr0cn+ndG4+1WsCpk9HkNKcae2YskD/tqssnFZYaH58w9ylaC/s55Uqn
/HF+3GzD65p3ghljYI1Y4I2Z0H7BPBkUCTRpNlla6u27v5h+/mGNJC/ZntMlRw9uXwP7Djej4ehb
EC/RnlA2A2oc8JgHOc4bDyJjmBELZ3QMK8Drzx3oNEfsHH04CYAtxMnsg4GM4hRqveR/9ai345+C
K56n4SV36UFTHR8pk84ZzU+FJ60Xp4n4TIpsNTgP3gnGL9VPoT3D0ZFDVlGf02v4AlhFmR7b5a29
+6rET8EgsphvLda2vgB2pvkPh5tqqwhoSELbFxMIyzHeQKi+fwS9A5mV0kDhygQNS5YlKmHjA+Vx
zjDtEvwQJkcuuPSlD2eKWZxLxk5vW3HGg9caXWGrvwUL49xvc4RTYNmqtxIWMWeqHz3C+Jc2axp7
8sjAr5Zfmuz6AaLohGYa164d65LTbTC7kZM6CX1d3yM0UaVhKyzn1vjTp8jWJjjM5kPOSHpP6Vpb
0BtL0NKldmgcEI6Y3HqAFEhh/wQjIhFbdNdZ1iZeRuTdI39bM5a6w3uguNwxDUzvbIcIkh2XFiwZ
8Q1wQf3m8XxktY41UkFxiAE91aNS68eCGwBCF2O4WB4Q7wjnC7u3vXtq6A0P2nCB9LK3xCSHyMiR
kXWc1rnAPXVhFHmut9qNzv8+4S7dQsSe57NO6obHbMe9tR0I8L2vxBrzaQF+2NyAU6oK6LqomeW0
8NYBgsXzvFMA21MDHVSIseHXG4d8HysBAnFIrpsuWY6GPviyKjbzqj319vevu3bdf3dUOZgSSA7+
9aaKyWpLURwaIMYt2ofa7qODqwPQVHKaT1iq51E7bZFLjZKQqnWJkmyQTW0mkZt6wkOwtYsSvpRv
OMfVHZ7y4REf3GcMyKvcLyGwvWlj2rXGZBetgSkdpfVcXdEs10K7DpACckhqVLoQi+b2y2xr9EpB
niKWA/CQQCeYOAmsCjFj3yPxHY/83eZ/zi+G8v14TlhCP8D3qB+xVawUdmDomm3nvUCsRvsYCc8K
DGyHYM346n8IVEu46mG9eBlq++dJPtyQxthkV1Zp89ZZhGlF/16NsYJ+F79lolp5i7z1ZehBUzp5
WNWuSOBenSLpcsTseTgOq9XmHwMsaOmnbbGS4Cs56nxX/cVD0Ib8NLJQXio/4brOzMp50MAy/QLx
r3parYPKgFjMxTtI7MQuRyBhS+p0f0U+8DM8KgCWjZUvMRQvSgm3caWDRbrzOiafDCt1qmDcrbQq
Qg71CurG3fFK1wTPCO9cKdiavvdP1cwXNehndLGOathCIeI6Dmu2UsP7ndELqJWAelNI4ntFrHTr
/YW1h7p6LliEKeHw2760baU+4AvOFRKqIYntw6genZZLgfZFiybG+M+osrjCGv+C1Wj1nJuS+XoH
73cY8HaVB8W0dBr64fOuwI+kzpziiVBxHur75BCBy5DqnR85pYIntJP6lWbm29bcNyEBfCHfwDCV
dCZVns3vW8WTbzHdleV4MPNED1ESnbckF7EVDLYP2UGxDPtO55t580nwRwTjDQf8p3Z61c9ST2X5
F90kKEJ993wqmYTdW0DXlaXSRaYAJFNvD2DDdkEXW1wk3Eif5dDlRxa8UMUXsbbdvnPkQN7R/K/T
G4OCVs/aHfkW3SHZdhXN3bxx9l71f1Kf2RvlzJTq0xylLd73Y3h2Ng43HZX7NIXzUU4M2zXHasNC
3tCq4YRaK2VdbAsgTp+Ko9k3Xk7C3hie9P0ZE4zyt2e14t+Olf4Od9g/k3y5PRz1M3iuhCY+rEsV
k0ktt1rVNmVsMPdk4rnmNJptBDBYd7CsOTF5pZuAtxc5sSGlVO1yKQiVcJkaAYOuandxOwTKywSy
Nu8XA+6+cOG1DenB3lOFDPxUilixNuP1GS2Z5YN2YwKx/x7awVyEmMrkOR6C7YG5bZZX9TJhHE27
Nte62a11htRrEH8fc79+d6hFizZyLGMmwjFgfwRtKLXLnZIvuBAIfXITkhM9e4FLDNAjZhFtkdPb
3r9krtpm+FpqboJUNMqUzoMdsysn6IySQj5Tjq+NRrW8BCNY+GpWBb7whTjOmMXxysrNcAUAQBFR
HrRJsQWE1EDS8Gge8B83L4at1DjzdvbAxwJk8Bpg8hlmAzwtdAPYrKR/n15ajlbiiSP7wzPJmyp+
3V90IBXVgyO/MZTecjWS6BRTtpYvKS7fZPnpiqJjNTfqe7UJ/VPAxvtMDXhOXRpzB0bJf6g7scZM
yreeJmXccqN3aOHUb+ZFvwodsWRVWvy0CKa4w1J3/WqWexHWFxTD75IHSyvP5I9DJLLeO63PI8do
5shWgL4w3y8mwrmTFFNp2ampASpDZMJfHDRhCbAZsbdirdQFpkxAfvdN7rSghbjV0WhcoQMuvIrf
mtY86w/LoHOocdo7kluRG5xKNmaCQczRbEl/OwWSCuyxGDpKRoJVd9D9+VjyO8CKS/QectCkV9H7
EEP4q8jeQ2Y52kMkLlUFVEKlHgpbVdxVyy9e9s5S094S+B/rWCpiN0zzjgkhP+P8YMR7Se2u2QR9
/N9llCjStzvIYLKteCimTikr+cV01GeybYz6ZjBKwIvbAA1hnIvV1vqTCnGwihhhmfQU9DXiutt8
BcrTJhYBCEkjf4Xy180lHEiUiyBBNnmvzWxSfVsXHfybbGT9L081XoCqhIg5k8ZZRg35a8i9x4xD
nA+1WuA/KqQsgzPmWRfGWZEqMvNaZfLhy3xNPGGR7+DRaFQLf1NdrYdzljJ1S8csUfcjhkJ13e2f
zyHNUQrG0GpKtogN89cEBHmr1w6a3uNyj8/A012suMNx7/qEQWaIMO9QVzg+UVjTFe2tBBvbsxte
aGX61CkM2F7XDSoVNfi+c9QBjfk0jOEqwGsQJ/aoLK6u4GStXC5Aj6cobCG9QQpQoGPPjAYNN+BY
d2kiskuqy2FWggTw8BHE38lTD45NF2bAX1SsaenMI3Qbz37DPHcFZGJAr3KbWODLYhJWHk28sGTL
VNxmMWPGsBfAtUtoAO4WFHM0/SZZYZoHSSqkALAOsHhoXPfvtNZ+CJTzMKqQ5Fs2XQS4dAtzX+l4
M8yZc4dI+xngU0/vCPWriwsBY1WAfMF8DHNuvxK7xQh8DfdsbUDJWVM7yl6DB+62PlkmXYryZv3D
DhlGnT/XKsdVO31G7AFIclKVfX/iI5SNKklLf4EM7EtWUpyOhP4sNRVnpDk8iWhKcHb43RVAZ/3i
8Q1zou4dolqZ9KYyrFQDWcCFTAlwZT+OwVOiZK2uqFiCutw/vWKAI9wGU3o+fdGMHjDcv5KOSs9K
hokHE9On/bhZN52bGxujBxa3Ntt6VAUygqzF6ZfQvKmgLt8N1nQ3HxKQVkgEQ7rd8/9EPPPuIpsJ
AaE0/5eIRsd9FCCTj06tIcTbb0bpVvDRCDGCXIe4nAWtGPcl7QUn81marKkv4niA8t6dwNfKHuSG
CgRyUlB24ZSBgN8zJU1LVYH+TZJIjzoGtDD5zvMlWox6kKndFTMm76UPJ/4CK3TJb50mGDiT5lWG
nBhXuK4tUcSptZinj32OWRwBJBJdiUwje+BuA0Kg6ApIix4p45CjGvG0+tzh2GCHX63F3cbk42h9
Sekj4nOG8RDEvfwjQqfdeu9f+hVves0F0cYnua4RPKLvHLJz6/Ti3HfAIba0OC8DUSpD7K5b5yLS
qz1i2uYvadCfHIIR/jB6Aug7adkbsvZ/vzl+mhQ3+urBZdZabbeMSmo0h0y3ls2Cs5xLhmxorZVc
fi8iM6YAo7yxsVRb9/XCcna/9x7inskn3sE9VgPntSGVGFntI98/Hri9sF3u8NmqI37nNlPQ9IQT
kWhJM7GvuathykbcBe/TU+xQaQWBIceOcJf7h4Tnkg46idcIWdU/W5rYO7grAMXxyUgsrtif1qEw
9WQevrg8MhsGljG4ijJKTjCBnrhSmSm4ztKmprHPxCCpZ1fMig1/sv+EzHzL9kdMvEJerFVQHl3f
+TZO/Qccnmc5cvugvpxMj6LcdoU8Y/Z5w+r0xrjctGs2U4xQBW1zsNOO4u+E4czk+lI5gZr6Zn1u
MMTFOuDtx2XZZxdx7dZj8NoCetQ/M+bkN7l+fDpo04dOtvDz4fHmQcI/VumPrJmVowJ3dI+c3OzX
Z4Y4W4cFnjnfsY7uCqA+hhoyEu1e7md77JCCKzGtfVNaHKWm7jMvuR8mtAuzqtZhXVIV/QZegle8
O8JR3SuXXsMyGB9dHcdEDf29V6oehLragDIgendK/JJiQe7N7o73BRr0xhHx/F5mkaWf++P5DmIR
JG4F1qLXl7dB3V+XNFrog9lltzVdFzbknMVyvQE79/tVyXgxuvLxGT8qAEQlUMWAz9wHCbASepjy
NGHHv8SIxhsb9yWQvCZ+YaTHCTzFkCVmHMqikTPAylaEt8DQltUWgU1ycio4CThx5g3K+1W6/hFF
YeMXWkkvDFjQWJDK5QjDyXXjQG9SUCpMT3LPeRJw3hJMvFDTLzvFxQUBkH8+qKS8FyrYGzcbxOV0
mUZ3IsgklOTYlVqyMGtP0YF/V9922JaU/j4FC7nCmXiRg/oJx4GEKT1Q0YxShhKNE/zqnG8G021L
NjnqdpI09OBaHvw2EyV6ijaUkbDBY9Zijjd76jmjWnJnnePVdg+4dh4WtH2/9OgGFvySRfK8oD32
uJ20MkIRtY+TeSH3OmFIoVZagJS/I4fwJ7LsO/PkFcy09HlriQyVgyUvqEEnxQfsv+G/NwiDrfnH
mT3IsUo4n/7sFULqn46KVngU1OXpFOHKpGrXDUPXheIeSsTimwePVh0wVAESdu8AU7JPZn8wxgn3
CuE1Tv2mxjMnY/EG19wrCUOkryRUdBfYwUkJkKQg2OiwutDvpsVdOkFe+iDnHZibRKcz7TvxmFB4
fYHhPHqRRjvuPINBoS7bvqtkh/tc5ExueLnCB4WxTTDdZB6HWqQxbbVlT4P0mEHQXHbaX2iS3zwc
XWXaFsmQa9Ny2QHTZK/XU7AxQfOiaGGj+AfyIBHQMu21JjlnI3rVeibzga9XqpMu7AMpaYsMTbcV
h7FhcdSrvmAT6QZUBYsywHyJ1T1N65b1vEel+u8pX/vT3io7rGtrxejPii2kYFJmjSWKL3ljydtF
jCLnlGQg47sYDL5t6Ow4HjLS1K8r0AF31budha62/qE9fhabpwwZjneF56RXKUMoZQKhGCaqfft0
rvYowijUBN6eAQrTxAJyM1xUz4hsbzKKXUGMGkWwAI6aySNMeZG24uy2SiGmjBcutbPZiEg2vk11
YkzzmNfJg8vYGl56ZyQwIVqaBbog8fjuveFxT+a3a+E0jh2pa2TV2yBlERnqt8L4MV7NfcWcCgSc
AuX8pMsv1r1P4BnKm/avWZZoj0ojrC8mZVUc9/QokOFxZB26fsAySDMVqOUthes+EEwRo1qqPfT7
tXy2n5GGU3lKfeRWcpAj15vRwHdZ2RRyIJHibLVDairPzRsnbIpSdkAco6LcOCDHXACBOV0wlmPP
1C2UDWMZEwRTHBIEtKKXv27scOpkjwXi1Zo0iqv8PbHwP+oNtDrx6uaNPT6cJ0cLXgb7Zga8HMlE
os1Cwk7lJ+NtJa+cVurlGx3KigBVSNwnh2Zrlr+QbuJMB0afe+6yTLxH3HMCz8F3V1443PZ6NQMj
eFN4NNaopvX1io4qjSnjKgL8WrOIiy/38TLi87OGGarw3/arQP5zjzm/rt7M7ouszTTQora9ayuB
seyw6YrerfgqglxBEBtMS9ukhuZ3oJqCw1hT3zh5wCOqZXmEc9XjShGJNeD76s9DSHzFcZeuldzv
1r9Ahlt3ncwIKfhOX5Y6RKARRXk1eaWxBQ0SYPY24S8nbMDO1MynmTVzq+Xf4I8ymBoF+WRI7esP
X+Q7haNbPnWrn/FYIxM3D1vq2dWZQqRVWzf4HTD5e5RpnqvTJ/mhAdpl6BHG/EERJCzrBdtyD0uj
TGmaPsIRjblrOA9Qb4/8Fh0ta9E6K7VYo5byOQ2sf+Cls+YNMmPUS2z/2F3iiMiGSrIU2xkPAX3N
eTelBWqXUxhz0yq0pIrHUjHA5Zvfnfg0yl5Zv7is/w2Sccm5O+rJhsAfx4gko0Zhmc7j+3k0w/Ug
BWNkSHz4x0seTbPsV0BakOCpN4m6uuqwUkRhSyssfAuInZd3y5dF+7WZllm27E0/6iz5ElDmxRB8
mf4d5VCMi/m2XvH+5LTcOGDmS6qy2SZTFwAvUoa2/lUbXeKzEvBYcQ6DYoIS4LMqT3BP4qfBcfdU
aluTseU+7eLZ+tkYXDuS7Z0rN3cA/7cfVkAt3bf9Y/UiSPMArpr66wPOwSxYBU8sO1xxlz9BzQgW
QP5LMmVb0VBY8wxH6HGs9/oLPLnLnYglPYqegCUrq07ZaJblkzMW+fI2xDB3p/+dmaqAFDmeq2mq
mISVmoa+1xlGQDUGpq/MmpJMfyWWisWiOWUUNZNcxGP7oot6PG5SzOu3LJXW7MvRgdmhNITGDHg+
wmd8eeqsAysQzbRYdCYtma4gq/21qWwBysqxXjDIS0qZHSZgT74GgY9bSH23xR66EGiJjm25LePl
urCNgQWl8vWsdmCekm0miRXB7LmTTs18uwY7sKheRFp38kZmXAlx2FdJrtiBx5DqYGeDeS5rTcXP
zpyDRUHtN57YkaK1Misg4BNn5qjy0iIE3e5rqzQukrvoFYt8KM+2QPWvUo4arARCudxs9Xq4qjdT
9puOeSeIR8OLrdGTg3ZSKs7x3zQXQQQ+DsOpj6cJIiFZFiNy9zs2pswX4u8L23HWQhbhmdc5UZP7
USpQ06whriQWqIFG4T1u8PpSEFBgRQEVIEgcaoXOcmw08hmR3eLbidT/fNAhSxgh9oEcto8aADAD
/kQmHrf4l+m2Jea/DjeLImk6fnnHtbXoIhJ0lwsGpM5Pb7qKbWOeIx5wgnPM3Toy9Nv/ffLWVwer
gtDEjb8vBWR5uRt8x+Piv7o0UJOY2LSvrDBVIY931DnJPcLCZBJ8QP4TpROK0hOgMTKKkpoX5DwF
9SQY/5QG19FRAF2VdirFyLkW+Oq0rmJV+18exa4PiIDLZGmgeHQcWSk5ehBCOKfVLqUSLR+8Zuz1
gkHNXC+W0ZcxaehCfy1ouNJI+WFaSdRaszQfXi4YZR3dLJDW0uWK6mBAQO7Q2+jigyT4VvLPxe4c
5pvvF0qPKjfHA4Is56DpGbqIz/sIsZ3rfjPaZzVpxzNBya1GCm30VTDv6bZC6CKI+8TKsowU/oj4
Qh21gQNuYgY6uyqo41GEx0YJDM7m9VKqPG/pNrhnCAHjVpTgftpz3qEY1cXrY2xGQnJYNEZtblDd
MO9QiC2d9/D28jNwp0yb8kEjeizoXjRBbgS4CHdZPSE0s7QELtWuklpVagqarx8j61lctm9NgFvZ
5J+1kRpM8LoTAMifOCKp8kRw/TIgE6j23pAVGJ7MgA1PvzwDmjub8oxARDfUH4hzR7KZ7ySzR2e1
sgQ2u7NweVfGPW0dBd2g+AEito6QDSj1uro4ilKZz5ZzDvhnisjugLATVp2Zjw40U0XIHmrAFcOc
DXaKiv0zt+n+syMZRqAXnHQeSOSA5cvw9LH9X53OqQiybwuOLxjGmIQV8OmLrCsCfZm3Sy6c93wF
v0EqgRDrEQt0OtPCWxDD8c1xYtMVjr1c9JjFdffh3C/YJ4g9gHsiSMgW3JcjDq5XH7izEpnTs9G6
lHFcLIkC9qGIWTgkwhCgDJQL99ibR8RWBBbahaFgnzLCSgIDJE1cLkzqeJIXQQ+QdGVKHuVP1KW5
MhrBGMUM5xeZE+3Z6F2nmFCQcNudHJAzHwKwGEM4RzXj4fDCL3jdro2WjhARr8SuzCP46ZnGJ038
PM9nBWC6XMuMSlO2vYrTcjJzWfvUUGdLCiPFDAloJ05fCd7X+mNe4h14EuTxhSm0NHa4XMlviNFS
1CDe4/9n01sBHfDZ1xfhL2V4zSOh3Bof0eVoLxyBPHwtiBpV9M7HQI92aL3+iM62hLAcM8fbItWy
17We2++mhb5lwBNO0WYHyMhfIr0jceLBJaNPoNTF+BOE+PfK5VpJ4b34RE2rmduKPt/VjA+tQGdF
JWNnv6pXYFL71can4egDmP3YG66AMAaNLWLTnVkEbbv/LNfp3kSz5gC5D3hU8d2V98cng7ZRwALc
YN5Lz+ZYg4zv2ajkmbFQtxOYDrL/H9vsC1RJF4gDTBFrENqyKzvBfIMKj66wsRloSXOGvTS6akqT
D6FZrMki0EqWdat5fpyNTU61YhRHorScnHLMKh5jppn1piIrZxrxmcxsN5B8vJsCfrXZrNQYRef/
xmAyGlZCf0IP4sS4W2XhWoPgt46N9K3x1mEBoUEJPyzpxWPUn0jUJJ4OGgED2hYGg0Euw/TVKMdt
zV6H+CVGIJ0EJKXBmQY/MzmMqHRXPMtW3zVZMC6dmGfuZP9N+1MHxafQNng5iIUiqN/544RxdY1w
LuMy3BhU/9+wQOQ2QlkQ7T/7qmIjLZUL/HmU8v0yZkurgT0UceBvk84dNaWXsX4cnWFbJi4Y+6q3
dkRL/VuJtN0JNdUNqb0YJLLOobKoI/3uYTYMNzXXiry/1YUn9Sd5V4QfYAyJ6LXeGnodUWZ/aHk+
hyVKNYAvlRLky0Sf/Nf6FtPhzXdBMw4Fd8t09t0lKLztGOG9e5CPepf2AJTHisWHDUJF1DVJSLXF
AksUbi6GfLLfjMne0epECvQJGZPSwJm532TGX0Vf1WVEoBTXLcimYb06qdxPUyztRFjmf7mw4kmo
s5KA7PK+CK5dhF6kX8EkH2NZsPAA5tYT0iVF45kRM7U5Q6vA34FqJuO1FiTSQBVFK/sy7Lf1pknu
Fome8bAQrCPDqipUeB+rgBjlvg4/1h8PH3WZI/1mYcQgPxJbxg72NOGjxIHPPCq1axcoKJ06YcGQ
Qh76tgPoElWO+FFM9oPcDBTqPp55t5+9cGhGphCgwRyShuFraRm+0RBe0BjfA6clA51g70iI0dNq
ouT0hH9/16SH9kbemuKzWnQf+5PWDaXfnEOH41ErY1GcWB1Fv0WWwKaO/+SGBO+OfWN/hRSxZaB2
z8T3d+22rH6htmDGViPR9psTHEhqgLwrEVv4GHujwXPzK7Ih58yjjxzY1qPZfcZz3c5ZatNMCvH1
lRSEMvpvDTuxFEaJ6bbeTAqfwjfaQuBKkNmEpq/q8YjZF3mHdkYX5x09qFRpBK0Hz1paucmIriRu
mF8/of8CEtXVbA6JhfWjZS9t2+Udjuv+cw8yxYGsWQfzTXfSa3y7pfksTiIpCaHX9wSTsZ0eJ1Kx
r+22EKrsZsbAaii27c+lKvfRP0Ew1clZK+fwpG58o1deyMjN5xuS/qyB3q7scKlI3yvoCdG4M/6F
H1hu8dzSxrwuAfDOepvbENrTr4btphWdufDj9Nb2ZFvp2FROGZigOuByg/1QTP9UMIdBJSrl66FM
YgDcShtppX7v1Hob28cM8VewxgMoaFReo5AEnW2WH+vDuAJsOWyV3xBDlNdKj2SjbOHcOyvx3lYV
1AR3rfWLuBSYSXxSBktksWyPGL1Ttf9K1wNUIt9ec/LpauoKuhsuBwbNFd20CINMrNl74+JLzdVL
f29J6t7U49mOaDJaUeOisDth8sRZz5e4wj4WHpZ/r/tmd9HZEyf5IFwshP/EQn25MnESJi2VPddI
Qku/d8Q/j+VVlv0AdQDhkZHqCsrczZCDfgL1uBGo44iYAWsyTCcVqocVbTJK6f8Yo9qTjr2cMNzm
TQ5skdfa1ePTDBJ4ObYOYtXrYF/GnlsUOrH5Wi+EIt1NKH1HqviQMpibnihipmcXMM2p11+engbH
9XWAvL0fgMvyKEDO5sl29jCZ7o05bU6I0goI+1dt8BDd4s3nACqccrjFtL7KGXjBcGQComhJlTlS
pku0L/PfuK6eSj7tA/X4F+kohATk6deDuqTgoD4INN/DqeRvT2X9YedOADID/GPO2HO5RRf2/Jdy
cFyqgjFEKc47nFL5/guxkS+iFngDS+5juiD+vZf1SaSu8ncRTDfU272N+bDW0XwkYQclpQm5x3Jo
MHpgVllxiEddA+3i6if6JKEikOinuepOXCLMCUEHHiznUOcmi1o/fA7nJXofNFiQLfWrQ2OzzcWJ
NeTv0WNsKYEQiWDRywHyp4+3ijB969QLc68uCiBSUTQr+/k2N/Iyt+McGCI7HOIvcs7PpjRhF13Z
9KT6w07P9bFnXK/arTFiryy8KHYTh58uWLcJ1WIomRVWiotaKVXnEZ6iPOImNRbhFW3GHdFZfbhh
qIuoLArJiWbBr68Wz1yeaVI40V3fff9UV21z86SRHCCAeba1isTNmLjqqPfqj7hYFXfTTi05QbpC
zDq1Vu/XlmJ5FYhom6fAQs+m2iD/l1JQWnwN6UW5ij7nVp9EsXrzWzgAKkKe7pd29BSOO1UtdUOl
KT8U5MVUH9PHl67AGpF1e2EHf5Tgzv1AgBXPzo9/nsjx5Apf0SCREd0ccZuEhc2XkKyj42T2Q6vf
gcWIPzxUpCXWrGNmwmGJEBvsLgcsMmD4X+BAVcLqQPuvJtG56YCE6DTrHY2ORNVNlFHWtqnAiyYk
MoeCgbw8lJCFzA+g2xlEmDFu0Oig2M67XRklvE3Wm+v4bGRU3oPU+Dif5v4oyxUN+3SP9/uYq4aV
9sRGL74Se1usQNfdr/t9nS/r0db1R8Gh0792vGrEiQdm+aemzJMgq+6W8ZPR4Yd5kazZiuVvh/pa
krqHFHi3+w+BvDaCkD5zdlAqjbe40f/AcnFEoneN8vqgW5V75YghRV95m44JyYiprZATnc3co9Fu
POuZ4Rwdb/dgqeYxe1Tfik8fEyOvEi57lRoQvksGZoHkU8dT1Ui3vvfKBch95lc9RWEGMmhwxLry
QuL73luLTSe4NyZi5HuLdMSbACSV2O48ymH+7QopprWKAeOhWd/gn7cXjsWvpDi3uYXrfOMOomnK
uIxiRmzywRKCMwHPOu7GJk2+aZSdTWvlgTV90uHsaVYRputnz3NUYfSwEXsDp0KSTRj0RQ1frRcp
XcOAYokwxQ6RRAclWcgYCTcXemb3GLXs5ytJCyG3aO6RgVYOnCnFyrfaBZ3rgT8QxYkgSdvNhYvw
so5MYfmhMaBGsczBw26N35AAG3AN+FCrHUCyunXbKop0qFXWOUcezhgsC6hdm8kgN/68uJrgC7lR
Rstnt5eAZklDxOTJcAacho3V21pZhtFy2mZlaAcYiX9N1kKUBrnYr+yVMil9YZ4OMbsHVy9Og5rQ
YUMxUUrcaHBLZHa7LZ/qQ4TCvZ3k1xXr+RDIXurGALrXeokLmHyloonacpoRukXyaQXBiVMIdXhD
/eQxiX1SeSWLDThSyMhO7xT7thzsb6TBfzBQk5soGfNNcurm1CKT/gcKTDH8rWyKCgbuWl4tyAGG
T14HqIJ9+NY09/STSYBogHA/6B2pIzYQgUWXcjuLWKPrQ7Tk1dPlmYl3e33dHxnoet1NUaKeKkjd
fFmlyuqTS4+lRKeY3yycO88QIxfjdTc0zvFCmL+OxAIrSbNssFO5Ujtqhb4A9bFiF17mLeH0mY9e
xFz8zGP3dtcWL9H0HUaZvPbUvGwyw+sAnSvDelrRakYRjc+6mqxXogkrrv1wGidmw38x8rJm7v1R
1jJ2qSRv43kNytvQY92CF8CIAmXpvw8Jhk6IfztSq81UgiLV7JOVFPtP+usItyugUxVUxEcwgToi
sujs2Vq7yt/drHVJxSaBD9hSmqa7SR13xjsRUC/Kg+hUeyNue0CgFX+EtzV8OgN3ARLwb4nrdnuB
/wu9PrWL/5QtEWRdt+sYuOqKzPXn/VYLN+GbjIAfG7RDmO+9Qf/srTkaCasGrUi3FJlpvoFlOF0W
fRryc3x2LnpAMRmEpqpyaVVyqwXWMJ1mk/7sKdBgyWk20T/rHyu8PZatDTd1i/J12BOJQy4TzkDy
8qbXHlDvSSddgA3Mxtvokdc1Q5TUysbKUDogjxN5OZtKMAdi2XLItkVCYkX587FMor/4ZvOlAd6v
ZG8TnoA7O8Pg99vMzT38n4rjSyg/z7K5Up5pPEywD+c+Mfg0KNF1kD8ZYk40qiXnekJoy+o2J8+w
sPwHOFO5qH9FI5usxtZunZGczxq2C1zT5xshtucs9WbwT4PVakg4ZLF7axJ1kAC2/O1IQWyLr0bQ
PpK+h6rEAsTlfTl3+M0i+U81jpIme507D/jb6MVm91iTlzqx1svEufZqMoO7ee7KmLVHXJdaTMRI
C4L8Y0sJ07/uGeVGyzcHhZhPn6RI9tCDrHohM9gI8n+Ad/7InKH6Jn+20dA/zdOjvJTbETLfNB5T
06QISyscSuRLBe7eIefn1+oJrVQCBuuGJBa/q1h+yfC1rowTs1OUt5qkGZILXnCQmcITRBO3WZoZ
QW7gBJTfkInitgHt59jmqv/iCfvG4Q0jkTVBwO/bqhTvJgeXB21+EExw52l9HAtY5ScyOT4YuvBs
kIghURu/9o8MjjGN6XOroXR9Ls47l4gvIAFuPHYptBABzJHHCIAqSojcLyBVEEAazk9mvXjC589S
+9EYbnMXM8T47+4ChPkBjeepUbzCF158q/FnHClVLw4k9hpdbb1zRmyoir0B0kcaavzlAlJrtiuo
+bBlWFAo/E80v3Zi7CQXyywPa+89eFWpfQ6e2PFB0Q5rdoKDv+LpKBHAPbS9KlHIxkdBIeBIAEy2
tJvhjZKoteCxDB30KnpH6OtqCKA464K4d9GA3viaQwR9IMwcxTvMs9uo1FgJvWeqOE0OUzD7EJzM
hDIXZEo/7JlP501MisLNJZvDh0p3axr1IpThBVgMoHiyUs0FF/SpQcBCJqnOvy93LsIzodTNdaPV
s9FncSswKcNceGGnNIKBLYHbvpoB/08IsUAqFyR2/C6xo+gAiMU6d8oizjilNJhzHYOjMP2zGVJr
AmfV7IjEFMWws3qzr9z/jPouDFK8EDHY4s46T7Yk620KkA4yT78GyUC71p7K7vcHzxZHn9vMXQ5B
+MGxzLKS5l9eADCAYFr6Fm+XSMJXfJOWwIIwaZ0O9wTye+X5JReJLbpFdd4UfnNMYoHsAFohvZ+s
rWZqzgpMzgX8W/sG1qHVJTabY61kYtZMLYDFdqqqYLYPGjTjYClnVk7Mm7pOtSzwZTa25FxoXFB+
+rJQnt8VgRHWfXIVddP2/lM67wzTLCqh9mesIqyeYPFeOST1dQgAM1zninEW1JezIkzUn8VJ6mNP
+RzrAyiqLzboq1ra6KUjEHwmpo51DbqTWr97nxbcGj2mPjAxd1fToTMbEn9UU+T2cg7hwY/GWl87
HGVN4tRkH/NBLgMTMZ5Qdla26JsP6Eo1oqa9TJjgklaZpPBS9fatf/W2bVsMdXsEJni53UV6t/Du
Wb3ZcyZ8+xnDenE18rAlngf+K4ldruT7zJGt5UDcNsB7VwQlGZmuHKDsQfRo2IO9l09tPhK/lWyP
SZeoTBgmcKsDLyo38BlI654MP94CS9aVt5fokretVckICJnG/KWkX3WuCi8dMRSOYUoMZSIYf5YY
7sCkPmZL3dSV3t+QC6XGZljkFRy3i7T3BdBQnY0KzgtKQm1/o4CwvT2Z5eabxgujwOthmV1sLKHc
wS+tUhCn3F+amRpdMjcycKTEOgR34gmSMIEMXyKJcEKvRedizNUBtNsxwkVYzGkHPlNoeIvc4WKh
f0rgtSLgfMjkqtNuGTb0y8OgEwqkLvmDcAzwQ3HSbAyQNa4xnU3zjCpD64uFj5uTXjBICRqS3qA4
CIi+ndW3yKSvoXbfad8T/Jr23d3CgQ6tcldQSwOnNQs+22FNb3JERbMEoG9glqf4yJOKq7L5FGCr
TjcfqinBrvA+61fpXL6k02wyDgWZ9VjWz/OYOfYmldjQ3zvPkt89g/Uq7iZOkeyouVUrUs9vz0bI
CLOB0lfdtf1B+tcAju80QfSMw5J19nfDRzVLIthYGG5sZV2HJLYBl3WCKhPgkkn45ELpBnUYiPT8
2FoXwxEDy82bOS37giwOGYgrLBdCgSU2Wu25Gmkd/a78c+NxD0hXo+mWOdjLtFT7ecN72aBMgjag
ZpzS7j1sKGp7NwDPP4ltYRa/w5/LLYG6hGDoN/yv9C1xgOBoGADmUsk368dmCRmKBhCiKd9mKSv9
o2VG5rl6khlmV79KMiKlyR627f+EHmNXxO4dTFYsoOHCigVCFARxRndcmDls8KPn91u52cWEjjfH
mLAI7jJD79HPD7usGsU+nVrK2G3V7JhKud8NEvwm/kf2RkYlGqkVgmBC4FiHPDofiuReriMWcsvu
L2m7hPHiSfiYmqhMofGdQQXRN8Fq6AKN6cXQQSLgGWdwdZWTqcxmvnxPHkeoaMCh4agRpixhdA/b
udg+y0m8d0koRqiJ7l8q+9VGnexjpZKGCYN5ZhDSFnz3lC7YNtuIZROdjejw1vu4+wis6KmilDBV
KzsIBLGIOUqO3jQ/0e9oXB/OCnEsjj65iMHc3XeapiWrrRi4Rx9co/X3FDlrHhYOFm0Fv02hzxkK
dwS4r0Y23Kq9MjCtTQTDJTo7sKazU4nkoGJXYMsC4ZB+LENsyV+vB6FnEInsZnlmoxXNnbnXCeWJ
A4yKxcdPgLHn9oBXFvH+XvssIVNc/4q44K5foo9NMc9NZ11kM/JWDngYbOULH3XXeMwUQSL+rvGC
WpS7wFGaZcDN4fm/4g/MUKhCXvW8fP/KvXGMAzfx4Ft4jiSHVxWCS9j/9FZZbxiDrD9ySk7EQbrp
7juUwvjMhOvYfofQz5mBjGFXVsccHK6PNA58WW69jcEADq/PStlk39X9J7nHo8eJqEqZnQRtEu6/
yJWTOZt9ihkEcjGU3cAsTMVpwPLsS2Fe2i714dC7T2XjKIWNvVqOud5aARtS605bwRIGeFf4y0lv
7mkr4meW15r3S+n9QO3zRvGow6GR54RADSf611O5J8Sl11DpxhNr0BdTCoFJKSU+EpI+kQQOClQI
YyHW3nk5T3ykxriPm5lAssMA0nWytjm9VaglQ9KtCtX1X9b6rcKkh3nHJIvEV0LICj/rGf7LkRaK
qzQfAl478WdGwYdkql82inL63LSxMUgYEXjL7kQYga3mGgmlPF67WjZ3nD7+P4xEAACltd9IZbjj
tXqYmskz4YL9p1vEYU6VqBDnMIg2rsDVXobIX2WY7SmwLUgy7ZM604i1mbAJiW1j/JcvMIMDdoD1
dKg5UfIk+w/JjZCx6yI6NBDQ5jef+J5LQMMCw/qIECXE/DbI8REXpaHJ9F2u+l7dgISXle2Qi8HJ
dXcCi8xFTmhNNl8f/WT72ZyqvUefo0qf9yZhNM+29JNiitYB9W64SA+PArLuihu85yJmt3lOsI9B
ge2cTsmaOlV2c97Vt5E6hjsGqspfL1R15LBXj2sIcIkzTx/RjY67fEyX6K5AqJgQU6VlRijA2yhB
X3dNVE3wABdqAFcJgoZTvOkEHKIcukvEZcJTf4DLpft/SNWU79K0qEpLK04QGN3HpZPu1wQ0+njZ
1YyMZZ/lfs6myqSDMnk9++GgOd3YKeGqLdM05aF2n5llEYIvj9WJa1ql4d7F7qiZZl23Tel0BCxz
LMwEWUASMka6QPmKvqG4JwN4MKC190J/G4eV/9eJ96gpm119vwZyjz5gM/QArK9wU/ZQ/7AAUxY7
S1BuyGTTeZ8mzHx5LqjtNpPDuNUlsVftXEQGN2E3REDNyygfVukSWJNAHC+PAJ1cro+OSJVYjpjj
mqLmRsQEnjHECJlj/ozmHkpvvqYN2aYrMQM+cMUA6W2f3bQDOlWE1rRt4ssgoP+6nrcYOPVOVmb6
Bga9VN6ZmGObDTlghBNZ31yOlfSA3fRdd9TtcQwMBr7KLUHzdl5I2thQl7HP6CCl2xTks3lIZt0/
LSaV85zj9iAQ87gpUddmBv8r96oNCBH6uwQ5Mn8Hx2hpyIg/1NjbAOQQXHtcTHmCuBtVbeuxNPaA
oui7tCbB393bv0hJhr1mYFSPHBYIhUqdkxYSPlWoynBp7LpQGVq0MAyc4cFPG5suC7NKkK2My3Lo
rEK0YB5kZW/lp+MSsW0utv59ySxFGGu5k3UGF0VUyqIAXHZApV/em8mzCEc00TGblY/XNYDWBY4g
5OO2M9ARG3OtkXPo0FdVNQ6dkaD+ypPvTm3WcXb/ieQFOv18EXxWoH0J57bf6HevaMtbapXYecrf
Qxw+hZuzEQ2TPmDE1bYOvz3q8ov+rvBafMyWaxTGElERAE2j6AiBocreOUP2jlCqqwA+gm7rN3/p
YZxV9KcddvkLjgE8wWqEQLVt8UenA+V8n/bheWm4FtjttjcRhvVP+LHpGq/nVo8CUJGLgFgfIndM
OD4Vx6P04B3sIFTqV6LyMsfhrwuBHKF1R9h3a2hgURawTpcadWiu9tb164qvQSRA/ppR5lZbDK7x
gomsA9veM5VJYno5cex4AmMtxW+3nE7WOTq80wClNqlFlXnoA/D9MWgj3022zlMjjt+Nv1lCfbQS
PceFTevijNZZENhAnDG8TjPu3Zxp0z2TnW7B4EOv5ZDLP9Owv0Hor6I3Ww8J4RlfH4xrczWx3ZsW
PAVTCWii9OAH0+Ac20i9ySpDxMddNg4+JYvlaZgaSI/0BBlRUMYLO67DgoZg32SX6A6o/TRRPZNk
nQlVkOYdd3YmvDgTD6Qx63+rWMowt6cTraePuGNivFa1J8Pm0wXvpfdQxNwLgLekHEUmEQAD7mYp
YWUS6bNZWHlbVloQsZeeeKYf2TJa0QPURy+hsluRcu5EA0B59j9Nr7s2A11DYWDLq8pCpRxfV6wU
LpPCTO8gGLzem475W01OYXvG30H99415W4ODRO18guWzkqqWCRrG/sWcqDR7uPW8TKXxraxaqv6r
7ieidsYO8j0a666VtkVgdyCDiYJkjeXcIG0huV0jkdt/3NZ+WjVLcRAdqOhdjhJHTDGpJKMMXzwn
NUWiXnSttgC6XsQunHLFDEetrJD97qimtVwUxAvjbMafb14XqpWRTd3p04BjuMHhY/KkPA+vvZbs
t59l0Z3wE0z3hLwRV+idUEDa7DKWc0zuzrNtm48Jt11iRf4//clQzrmfyC3/itjJiVI+nFn6TFD8
x7185jpkLCHFy0AZUmW7uEh/W6RNc+43O+vw+GZcN8N2lT4YNeBgXNb039Sxac0uiJxOQDD2A6io
vdzDZ0NgLyTLhFMuhgvPb+i0s8nke74VXECtFkDf1pX6feRG//2picLZUKYU7/eSoG185pT+8G1P
QGm/lCUqu7K2k0KrdJ1kN1dllVox1GntdGqnVQLoR7IVzUAHbO4bdsuY+qIq9nF8ptczuefoiotf
7igFJ9xYQzFgVztOWPzXg8eSapWOgJm79pHnq7hq+KN4AmEqdHvDqnjga6u28nIZKZOQEVsdUAzM
Bzb4LCnI4yGpv+q6YTf7GuYZtGTBHQMLxVI5KGKiQQGzg1al4HZvrqANvYKXU5YMN2dTVaBa79gA
PZn+6EKjcJfoJAisibjfzZRzyuXM2yKo+UnOVDvogiKjIPOykZ/YYKfzYAf3il/L1lxbBpgB4M54
77zadKRt8cl8H5dBVCRvkKPP9D16zz86N07PIamMTUzSh1S5ZCXLgwNDvC++S6OKFJv090DUe0mw
hFn1/946NJA/p3VxSTR+VjXFZZzUaXOipxxs3KAZug77VwS1dEGBgKzFLVPi98tRYVgiRib37v+j
tp9aIIZl953sSAjOEcKa+QPy02fEJZoE1G8UjKfs2BnlaWfCaDc6tic06qrCr/V+Kta/noVYz7U5
zJMsANk7e3siRwNl1babtfTEVG8mJrJmMRRjtCU1JXHq43Ia3lf8AlD2QZH5ETNXqi09ygr+vBvO
RUmx4K0DrfhrBOWZ8SzsOjvF0xc1S0r9oGjVGocpulFJdu6XXLrXX0KoKTx/8waZ3cdNbpt6WmXc
V4VntaSiHwe1Ot6s6jmex6enokStw+99OCCxhADFefLxneUdTIXt3rnmiejQRyABQvRSw1ynoOrc
obeXdSJYySEhkwV31etF45UmpHoPxRqBpKhb3SMVb7H8GkwAR4iR3vawySMoUCHo+An3Tz1qGawg
SIHRdAAKGJ8Dx+p1DcWQitUUvaPUSF/cOKnmLDwfOdR++LG/Q8ljwaz0A/QfIHYZtTPBBRNFWayP
4/F44KCD/rJNJDnSeKLjcbZQWkHKL212FXFzJfBZZ0Pgd5p7hnMuUswvwNScTwJf8ZDksfRkMW/D
mLcZADAaSnuaDTHmA83EI0ztKkQ7Ey2pRbI2QQIo9YG/1VESy/tRlNx13KbezICF6MAEakkbBaVh
qIkJZ24cOWUwf0xnJsszF1fmV3vfuptno3QKZMQKBHVfoEuGduCBMJ/r/RH+A0vixWWj3V2DywIE
dtdh2FDn1z803AAsqC5+tWvlaG2Uss3kBlgFuUkbvaKQMGruO+YaYD+ykslrJKrWLlhgGdRNk2yO
hF+t6/kdDQI0o8TAHqWNkn0lbvl83NS9xQWZP3OmKfQkm8NgjxmTiV/gLY3vzo95+p+YHtxUc7/e
MxXOTBAouWcShGWKHy7Sklv8XS3imK/cn1J6gyyAf4FtHuj+m5zuCswOb9JCsF5UHxhjP7R5HE9s
FfOgRacsDX5S14UTiag30IpzPOK69hXxBoWGf7DBm1kYLdzUZ8z79bdOij20Xs+AqpnK/SjLWJCf
Zo3jSlmH//4wzt6mrTB4Bz+KXqSpufp2MpmR9RwaW+liWi87zIspoDcSSHZV37AY+gnjmB4pAC7J
Mg1wOpTlYcMhkuStVj2RaxqD/WYvCPNB/OtunjV4R3+2Nyg3zOtzw9Fy4N/C/LNzS1ThqX3Dmcir
z77ZKvdAaLZlG7Mi0bEtfs0BdRMD1/L93CyXFm8LdbgyB1npTun0kFqWcorjT/15ZOUnT0ddoCOM
YfIepfwtOBGkSNSa8+VoyQp3utg9mA+bDNLhPmyhlU6cVAPOZuXhjbpOBV6n4jHFh79sQHKmsrVx
7SFgFxciZZMZfcnpsGsm6pHBriFC5oeLoBOV9abXcSIBsaCuFNur3BSbNR4EPgxrWX6TYF+pptTZ
TNEjERqYUP3JCDmI3dfZx730oSiCUc0eYuA+q8+ZmDJAfcYo84BE9QrOwfk4ymQYiiobGg5MSMLY
lzJoVTL5VnNrD5dq9Ay9s68aV7otiyJ8kMThrfYS9bPLytU2MUZQ7/sJhXH2QMTkg63/oqW8gEE9
uJzXn5ssvD5MSTNycIC6ylUea3KBRvg4Hfq+PdDITGwgO4mU2zUTgAJSYf7FUO8vllNpUt253uYX
xvj4HBJHUdquS3HxfH4asWDPdgP+FC8Vgso4ANq3nK5pRSX3N2hmAG2wv8/ZCGtpFA7vmQFLcM8o
Ue2k9GvC4oi4fFB6l9szEFQjYhCEbWGxx1ILGwal1ssHMT5s7kJ6X/5K6SbZj7S/y5/mlJzFetEt
xe9TgPxT9PHJcZ3X3nYjLNqVMa0vxWN9N0Ko8Gp6XFjM1fCPpcPGLqxJGgSaZIE6OQnD2LqDhmxl
JtsqdfXEoyUF+2R+ZgkEXPDKMY/Fyo1O9Eml7DkIHsFu5nvHPDOSCdSI1+zQPPjrcACnDRP6G3NK
VurW1jvaH2/psQGhjMcFDIAYqePnAU9J+zX+srqLgoQalJivH22ybfpd7qjFPH+kwkkxxqCact/i
AEXpInMk7Or26vKa0nAZ0BcdZjJIG8X/IC1QryxdfqRdKO7GI+3wdWbIMYGGjdtlCuQARVeyAnoV
kUcfMO0GtvddQafGYpBdfaXQmCbWJ/Co62C34RcP0tS/pOdUa2GY/lWcvJlNJhSUM5Kh5bbQuJPq
gpYdQMgRDRhx9j0rmoZN1bhvosgpr1ws+wHMkd/eXB4GMYwoTzjuYMHMsaqU/6oPtA/rFBO7ROef
rjgKyfdHUMUVyIo0C7FGN5ayf5+6qv8b4RS9DCNq6/CgoFkKQyMKW4s3I9H51uNUEESVAPJ4X53t
tjaCcUpBdG2U9i8YAVVm7tGA1hbnlsBa0yO93SPNLTn5pa2BRE76QsHlpA572VTYvvDXDD3vK3/Z
nXJqsOo2Xy7H3nbFviCeGhtAxCB4NCMRfvZYr2jj1EFxGUgH0+Ril66qJfnKsvoHwkFiEWpoaYAF
DubufJ+RiqInHK4ZENjH4VbcEqIBoOr66CdqFrD/IH9h9EqzMcl5XHn364RtCcfhVaV2NuuK79UM
jlG7P7v7+JlzxT3uUXL9LbHCXOTWpf1aHKuLJJ9j/nZ3cRixNJsOReaEzxDyPhmYFMWDFXtg55M8
8Jov6iFjSQQ/U/9+Qsv500xWVO0sizAtdifT4ZGTqpjIWqoubH7BVoIFjLOShs2hOn2x6gAq5aG8
WStpXPt1tZyRx9z0iSTTFF9TiMm7Vf8+15tZyZppYhMmISkRHIw9ZWaTPSatvnidmDdy72lqZtxU
r0+DUC+5RFGJdXr6MTh81L+gXZ8N+64LeXxZ34QZd9pRG6/KTLnvFefllMkmx9GFArWk3jpMEv8p
xH3ryMuQ0V7FTYZfMXNWMERxF6H0rNrQWrs6Kb9ZlnjvLt6sNvJfYyVgW0k26cjF9vgvZv/o1ArG
e4Mm1zkjFMZk8OtNaxkOWLQOj1XAA9cAtNY5mr+FehlsL9Vb+ujPupeRc5YUCbc7TWqXOKRxU2AK
KH9KYOvK1KYfiDG+EBKJ0GQIet4VGZz9AfmCLXJL0ykkZtWu7KzbA4Ur6YfpdbwTvJ501khmIh0B
izZ4xcJwde+NBl2+mpiK0jiSX7gVc5ECPwKIQzb2Yw0/cTBll6WQL9TOuqjVSBfzc2c1ZutsVLKo
LpkQXj8ETA/UVqWkWX86sGlcaYP3CzqToZn3vOpBeqHSIrb9HlfxCQLKJzkd719GvMUmq+3fZ5ee
GsPsydIoET+fJdT/Q8k9WTZJdtJAQYWgCPxWnOeFrcqYRdG/XihDK4p5s6QPpsN5jNWMpQhndszv
Uvky4/th+oCDAiTCPrNbdNR/76Sdu1AnK289aE34eAvmwtfUsMU9kPz0c9EYwHL4o2ftEPrpExBC
JPAiMTqXRfELUgcdJ08AMWgWyHLW6QaA7yn9uPScmxvt0q8idB4uFlXDGIZgvbEAY48CvZrQN6bX
bs0Ylch2QsYIogSLut0tlXZ/lL1p+FvoeIO1mWagvfQu/oN/VJOHrp80acsqKNSCDrfwHy0CnBGp
m8SE3hDwoQCpMuj1zerK4w0DP3A2PRwWM2+YpkFzLsJcN/CDwnnIqcx68MZDunfsHCS0tZ6i0boS
fI2udSF1U+5o2LW7rgnDPDEHJn6M0IozeSO+zV8ks6ClD4CpPmA3Q9uOSe7PaqaKaoOZnT1cf9UD
0zSzZEwvga2v8CNf6Zm0O39lHwtErRXXEJm1oBC6kZmvrD5JzHB6GErltJNiufnUpCJgj+USPj3G
1ei/fLyWqJtq36eDcfa2BwJUwAt9ftzHpDo42q1fu3iZVFORI0amPxrwh3stJPvIYAje39iHdNNH
3qbanSd7hbjSMtvad5z6x/cdQw3hKpI3jhZE9/DnJbV88NBoPWPrvU7vavsbzTePXLLnFL0Q6G0x
Q9P4e69T/p/QQ+nleJEWejlJiWpBru5poY5Hwwcx6xETz0ypvBafJt3F2dnVrovYy9erRGeXqXD0
TR4t/2ECyY0RN//r5LWjtHQBhHVkXfCP48oPBdvcOswJe/62rYEZLy1G113Kgf2DZuLJtn2saNKw
JWzHT+tatawjp6lQOcf7h8gUum2B457VRLxW5f0vs4ReL8Ur5DcXLfXaZRMgskx30sgFJ7PEpiYf
WZGexzfHSTClz9nmqz/K9H8kPpUqIC687DaiuuLaxt4IaGsQYDsa+txwsNvma6nM0WjPWu7TOt1V
LejL5WpfClfWFYHOhyEj4FEzyshQAQer+DKsGz4VBWKntyA+b7Hj31uQcpWSkffuiZIZMr5qpFEO
+c9DPo+5HDK23pONkkwnqzat5SPOVyt4Ly15iPwsRUcDxi9rbh0ROJi1PXNqL20Kk06I47UIDlJG
wyWycNQj73eEpo3oZkMwiyB4FZardO4B8gETDyrxGhozaLJZLy3iqdGA7K4azT9I9tDVNxR2mPSL
gbg63jD/mPN3sdJZUlS2RO9sm6z1CXQnBemmK7avqyCKGbFgl3FChF+hsofzn9S01TPn0JDrpkz0
y2JjrTDhmSOCJ1YSacFqZYzrJAbZetQlYQcNqI5pWLJ8sFZxVMuIoRGwMw3qM1feF+vxaIxHB4SW
P/wplJcK4rij4XkpYk4nhYalZBIFN+J266ZX060D7wBgZhAK6dNASc74sJLCOjaWY0GEP32WKdL7
IJJ49Um9JlDbsG9z+jz6zQ8JI+mGutw1XIndFXQcPq/X80i3mn0uwX/NVU3KHOhqf3DozWQuw84I
bsH9vUqOkUpRPpyvUACmRHVlMmstlf2DZASyf35czcZNiiNUkcQrpVEus0z4M8HItGqsAqGN5eSS
xO1Z6jx3pnEADRUyC/yHKlNTEnWxPm/Ae02jc0qaD7fcRgn5Eb1mRishQHHcVTVvyAZ9HtQ1za3g
rHyW8h8BpMGsCgvbhpb2YbVvhet6OJr0OngwbBkHLBqv91o4xDyIPqJ/aeas2fbet5EW7xWWWlJR
Xizx5xJHnE38a4D8oVNSM5AQ/ygccA+wu5znNh2jHVulytbG9bsgxgNWJBvdsxuUFmUzBtMYK1B8
MKvRwbzl/HBwoIycubsotOyFKkqsPSrpD4LJHKK9qFH7uKP3q3MR4pUsEgWcTRBighmqg/pflTXa
Hww31AQHQwSgcpw1XX7JQPFdAgBqZnjdQ4cfTt0NR12+EnL65i/pmYaFRqSWDf4D+oSqI11+tmrB
B1ZpcE7CRo7lxQu9qx86wuCQN1EclBAqdrpfnzaT1pWbfh5egVCUapraHnnxRS1q5bjPvvFMk8gY
YroV6yOXBN66QtWHYsHEnLXD5ohJ+D9rARJbwO4qyNFDd5OW7uSv5dVQpZ6fAxiP4q/1PgieW9mN
3ylWN6thCWthbmgpAT8VSu457xw6WfGgJvo8/3oXnMFfwcYzvGS0uTMZa4ym+lieBYJO53v3TpTV
2WhYwztzKJFheY4U2f3VVjt+Rj/I+M7fAoPfPObexpbg6R7gPKK4fyoot0EMTvHXLEZBAYCPmWka
E54LqxFQW7wViQTFDscQwNDhHLbFnvknP6OrkJnRXWn4FjvKlk1R/kC6e99JW6H8AqQ0u6fzIkBt
zDfueMiG0gjKjTyRnzEs6NGbDAo7rIwO65bpxJ2RIakEsOQbwmpuhkL/wF/OQ1GF2J8Rh0LMb1/n
r9w5fx/11pM9PI+LWi3pwkakwTqwcufZ7i0RJunYrPt/k4zsPafQnv16RYOoZHJ1SRYoZe5gIoYL
6j0o2g0XDJ3Kq6rq/uCjiIlUAqBOtrkdZVhuUYC2Uy9brSXNYqDZQEz+qNpAF7pk1n964gewwEKJ
3Rf7Nnz3w9Ls+wAZvDRhZNeaE2D7tXFpGLJNRGomv0EmdNQWG7pcKPaBoaW97o33oylFnV7X7kLc
OnCiHA7EkZIuMgDmorTJ7Gszhihsvu0Kci9ZuHI6AflqSCWoZ4T16wVystz3LlWcWSdYL2Tko5N7
j84NMxatr9pCT4RHC76yarmLtvQrmnXKLn9atFn7ENjfh8D4reACFsFlbFQLpFo8Da5u5Zik3kKK
sOF+8f/QQZMwHnZugZ813cplokFCANWMjnyjExR+OA5Bk24eipXfjkSLtUFrQEUTGagV4AUNi039
s+5jsbaiNUVa5NIZ7mJTHtfMIDoQlTsZYDOTJgpCFoi4qneydbdun34s2oe/GBuwqZ94FHoQ/eDO
GgiJIGLGE1aPJTYSeoTBkL75C9LIYLUUB1MTHiDOg+nfCWlPn3bvMot94LrSB9KA8NPIBh+rA2+X
bcpchpuE/R7IZ0Dpxo7poXrNBX/YU8ZMdga8PzhVHwv1H9F0LaqqrtiQOGyo+voTwtZNLWe3fZ1w
7lF60r1jBWCgN5AlguAGjNF/56Y0IkVzqgbhiL0/x9LpzSb9zQ+go+IZO1culDduAJnHH1x/uDip
NXQJqhh9L9bfCbAqU1RbK8ESju+ONQm1BatDHIu3EwNYN1mz/LlVuD6ayEi7ewSmemlpZEJ8MzYM
73cNoMY2+3HKdANkzHFT0J9Ff1NgWrkO8lr2UdITdG+rzJ6zwMi52vzjXbCJllXyvUYvwxwVWW4P
81DxS9QfOG1jAFtU0D/CipbZt3x+38+APjZGVtxFESX8qLAklWvD3zkTj+ZvEfFE+jAk1UkVk+z6
f9Cbjqe4dWLaVBLHJc6tW7kevKMVsi3D7s3TGJAR7t+TK5RKpNXbWFODt3EWPAjPiigRGqBCSy7r
0j6oHKhs/RURWuvKtw/1G3ZnTCO6iGzAEXyLDq5qzSUCdnhaXa4mf4cCz4hpn0YWaWYcX0GNDaRx
jW5EjjyVmVhjw9Mmrp3lQghOLMSOmKl20/R5Gudi8L37UUlIrO8qg098DlQEWrBOqmtpq6G1svUK
Jl2Sr3lyCxGTL4Wuu+coU/ApOyj3CurPdIQs4tv+A/JjaQSJ0TZtuuhToUa74kIzHs9sefhgQVAy
hQcNqyV5DOkxXlMV5DzG1QCFGaDylfD/iHomeQsrlaTgoXQiogwbBnZzS4/nsOOob6mPp83gjC/w
ZoOooCNN2xK6+W86rBHyTw1a/01ojEgA1WGFRFbNwV1Im89O7/3wQqE9sLelozOMljDL1yEmMUST
w72TGQz+hvQRpzH4mvM2yTYJ/+DxfLpL1Oq0s3L3s8hWCVz91DkrwmNlOaHmEJaimzLbBTk3t6aQ
oAhusyKnfL3NiLBnaeDB3ggsr6wu6fm9WgmhRpAjmFEMDWtWPurxr7ZJPoxzrJa5n+Fs8328dWEi
Stimk8yUTsHCsK1zdJ1qRXG1f71WuP69G3IvZugwql3d+Uht0erBy/zfKKjtJX8k+sEeUupMkreP
r6WSGWb9FpY//jdislhZvroJ5jYZLSxNQpOmX1j6G3EDu9FfKiSL5A5PYe2Fq6w5n0KdflncDcJy
dOsBm6KVkjAHXFMVmS3DMnmnOCBIJO7nO5QQIdLXm5FPu0WSL+uqYGl78fK+/hO+5BMmX0e4MQNQ
WOHeHEboHsiiVLwy5HMNXj2ZcXpWU7dd1gLuqDmm+RocDSgW1QNBxVN//Hs7AP5ZQZqhqDDjvmU5
e41dSaAhtfSPwgzDaaObgBMnDk/Uu2JwDALec8N8DfZjE/maafDEVgs384UAwpHlCxAAvQFIMMiX
fiI7a+FTHCC/J1FRQ1zaNcRL8msmMiy28pDgJlJujWM3uxv8IIkmTEeCFfp08b5J5bHiLWNnTMAI
pRCGa4dJe5YXQuVg0SVT4PAvpSEScWjcGkuaB/PN5zT7c50+GWGlvVcmELJVoOQzju1unOyVBqXJ
nuOmqIMKEJvBfDBtCvytwnssF+c/Qe0tFslxi7E7DkyvqcmxJu3h7vDIBEOc5qEJ3wE8pv+sIOWr
G1ZXJB5bBOgT/s+p0+AJpWrQBPrvXnnGzerWpS8sBSoT3R7FIOfEuZKso9jCcJ4S0NyUOrx/ceN0
1cBdlBx9LygRyg9FJGcbXGNpcTx3PaDt+NeneR8af8BCOZ0oNdDkZ1AepwJ/Gy5a8/H6F7ms/cx0
BYOQt75PcPg1IxV4agwNQBBdjoH1IUnaUQXWch7W0HB2T5pOpxRn7o//NRBeTsm6EHSc9qSlSWhw
TwIdiMYghUFPA1gQ3399rywbg+jNlq2AdhdXI2PfKvwuJVBUjnvEVZNiD/SAO0fCNLEtK/nDRUNO
cyAXbeFgdbK+lUC4kBoTSb/mkw23uJ23gEo+lv63sKf1aqbGmmRu/XhSHPI0xW9kXtsZiQVhub6D
gP7TREdcjK6ygupydU9tV9jm8VHLt1/PoRpKkbYGD95CQjmnrpQN4Ju8R6WV8THIaknx8D6YTNDl
d/zmoIE3V9cZmI6VEQllj37xm8bovPLspZF409pepr2bW3BLFqrmD0W3sDI/RTrfR6/g+INxb4r2
1DL9TQ1lSPjC276J7miINaDFJ8BOET/pNDu64LlxR/qq1zVDqwihJM3EBCGnPN2eHYjdLAdHQB44
3EQ9aRbH3HMKklXMWdKrVEh9Z3PlojSYNHDExr9ZyLwE/fJpDr1QXKxGOpqN96Oe4YRcfsxAy85a
rLeGwSpHKtiedX2tJQ4yXs0thjflEG8s0LeBNIN2P0sZhT+ZHhx4wZzk99KSk6W6WnfyxqBnsy+s
ITrvznF6ECLN2Udpx0z/ggG8+y8CcmJw3vdcUvyk3U7pLDZoluURqPTntAzLu/zUw+59wwGMwrUb
vi+F4IA5VEvCiyO4Zj2JNXlKk+ySJfSzqQ1Yp2S18bE1rEASkDEWPKvx23t8PiYMgtYHQrgcTv/K
E9fhPktfKjqvuYaRpWvzQFPi2QMxEQ688IMqOuP7HH9y5eWz7+fvHDKhlKb8M02l/OK8auNjxti0
tYa1blvNRV975+HITgOraF13smFPlqUawYiFZ1ALFZYqbccxHiSy6JrEXAR/7R70tFtkccWhr3ED
ieRuErGuf4diRmfleuk2EVGs9O/3G+uT5EVLzH8s6pr7nR9NvoDSYRGdMSnglB2gKMJZfc/S/UA3
ScLC/Zn8t3uKDDaqavAtVTx+OUKH30aQGBChnekQDrbeqQ+oly62AQZVPStUPMZ99DzurIVOAbxu
Pc55mWeBOFYqP/D5zimsiE/kGhq2/KUotXM+Xpjt9vh2YfcwUg+bVzj1nwl1jn15hXagG2PYpLBT
V2Y3IEJIKat4j1hoEZtSTovpSTHJPsO6QzbRE2fzB7+l1SJB+QSB72VAGjsWqyb7LXlc4zA3XzoW
Q8S5gUDBPtVCI0T3YkDCwMhLZvq5OAFuLqQISeIk7lJ1JSHNECT+wPbyYY1/JdQlsXmTfqSkXlwT
57yiJfFOqE6WNvFb7tzvRxHKSnmEASzZ41LH5++b/LUKRHluDrFQYwLIAilaABa3KEMVrdlI8fOq
TfgFef/+rYuSfgA/B/LqLKaho52DL9M8dY1uALrVPlnZ9q2kLNBZ0lISFyqXQWcfxuNqm7bP508X
//JTeGpL75eXKGWYa/w16ueoNxP6PD8MSnIm8W+ZiwhNgYzQymTu5SVGygOTV50Yh9Q4MNgBBPzk
rXqE54YdMVj84euZAJFyo3BJGFveVGxFjXHVpP+5yLFVgnGoQdqdtNWD/sjCPEUmhticHQvZfDlY
/1z0EXrDs6b1jMAXWJCi5eCc9zlS9lld0lyfmBY64wIf0pBe40ZZ5cMk7E0m8fsEUB4Ov2gEjCHu
KbEERV/f2ECalpm9WID2mhokAOIE8NEyvD3X7T/+3p7idPAtvzayujdbTMy9hEvNZnISBZsijRMO
oCclpSGZlSwrkXYI2kZkeAboICoz87s9yXkhVa9swoMwus47Hr8FZfmkRVFTIn92m+R1S7E2g0Rd
QPwEogq+8V+uI13ozT8NQDgBlTlFC5SR4yp8qAij7BYG8n9sbY3IjGKAjrrd5wakOYeNVJmUjpfD
zDqfraeVvUoUXw+qFPhtiwmBuxDahPuhGl2NFKqjkY4KWyC8uu06+3Yi79nGV7yMrK5M6X4/zXxv
NYTCEtwbrTcEmmq9A8y69AW1SMUoOhIAUGiS+GkBU7m18b8vUuVRvQcckQjTaMlPTDyUTPmDg/K4
KXCo/cgkNgctrSmbPC46pctayJ9/Gf0jJF8O3GNAGgeTRsyNfjLUiN/qNqKDHyBMgHCV17CqRydR
m2Af+sYIg8q8WtF2O+5LBENicSl3Kk4nTyKPceik7Y4R6RMljwOc42Hjjk58CbWW2+YcjhTcb2mv
lC53+DpDZoCzdIaflEu4oujTXzjCha0GyYCZvEC2Y1IJVCqRa1VyAu9+3iMP7/w9ETUcc1GsajvZ
YFgrz6+xjTA9b/wKKHDIfaHwvGE/pJJ6cQafGVGBvmdjp2NPM7feKGj2bzV6Yrz80I/Wm2CyBr9b
3/zfiOLvWtP10NrJ+mRHRudXJWJzq8CXunbolqL4LiceYyzCDxjaUGt81k+QKtWo39yrA+dNgVzq
pbPIUSybJpd5yUy0bc4564RnMJJ/VKEZuN641rbudLCLLYleumEoTJxLdbbPfNy9qrG41ROFy/FB
UGAPaxbJPAI3QnDUelpG0xt/33t4IKluBTeAzwS7aCAnF1RCbtriKbBtPLD9842UhBOu6hw7p/PU
Imz8SBviQAiiL59uennMoqX88QpNvEMOOAidlu674HKg9ieUIhcAeRs2Gnz2Lhri0WpG9fpJ8qfA
4nnXSh6vfKIukymFLwxr0I+GhNsgknKCsZo+S0PWY00Jnp4ATZuG+cYVpU8BO1SePOENrJLxBxSq
AVCYfVF2V2Qqn18x83kb01mHG2xOROtPDJukPI08Z3C4wx0VTHqA42s9ITLfSFUzPXL4LnsXDEk+
CqYHyxHZT5qX1wJ0EkHiPoZ8pxuBJPlA555VLwF8o8oQOE30ZvJ3U8TBTW/rsuYMB8naTPf3a0RQ
p9DATzfEPSkmzvhACuYr9hUaIP1LigI7xMPBPDrapYE/waH3FGQCF5CJ+MJuNADsABXKiWM9iUQo
s8SYAe9cfIWuWqSKcIQatANBnYcNj5mUs/w1ezSs//m1CSmyoUphpDqiUUgcL8G4jNtOkuwrVga9
FClgu4N3eh5VLeQZOiR+5bY2Pc7eplgnBsUoieSkDBLm1WIwuThPB7jvLkdGVhp+WEldsQRGFw7Q
znffXDoncXPR7gJljPSjbPsCtz6Vccd9bKSJ5CyTxqu/fiDIoybeVGiIS51/zhRLQdiWihqTsF4s
6dcO8DqNrIxGe/pVFu0R6VC9afQptPyki9bEp9HlPdRfzSagH6f1Qk/zC3sHHDT44kKnPPfcF7BV
0Vmivbn8TzRMSg+ABtdh02sQijP7MpQGRoe2iVXaJyhkVeSsnQzmdgoJdVkqsDuADz3H3Q48XYQe
FanPTXkGtooySMcbPSm1llfF89kA0LLmlM21iGJ5KvG6tRLFWZaA5eBtspCXEPswQA7ivuf+Jooh
FUmoq635OcHyKoRLvOJeKoA4qmyzlFSDd6vKCrrxsD8n23YfI8/yiKRhlExOxjo8iI4tyVQcUge3
yqaN1ckhxyWcEJH6N9JR/LiPh3Y7gd5Uwsnakl2ps7MizC/uhBStWNP/6f1GLuuK9gAR3offkl11
YW9omYx4JNNbHHfcG0F6gPNR4jQ9wqQNT3G5Vqy0I2d1kI8NtURimS1q/jO+IT2dAQLw3NHLcBCb
RC5dQxk88RTMZPwV6KvamDp+3XBRAmJ41LO/YbQEW/40oloYh1AM54dUhXAvcEwF1GK/C4XgC/sD
tyvssLHb9qZHkRTRWLqN05sISjVXCIFNziauQxyVjlMvfUOI/sg+UknGF5twREESKJeSg1/b0wMJ
gw5FHwNmGp0qU1dtMuEsr/fH5dHEWNeWJRIZSxivJNgsmJfw9MnzKy9y04Nd3p63U4A9a21oEkqw
dw9jgaxxNMDMyFkWEu5ivr8gvz6m/UpZAIDrQq1ujEW7R+Xm0fBuNkCufWVqcmNVhHKDGBPg+OuA
CAMrnEaso7z7u7GAZjhllKUgXvTOW9AwRzHudlxtHJ7bHZ9rgOhWBvWb4OAPiobBzrfIpZlnN6yl
mGfigFASWJDc1LKEQVh4SlbUCrifSFRQTikJt6PJi3WqmBW/azrHyjrjY1Byu7Cjaygs1S1ZqIQq
FBWRaT1em1RNIFwjFyG/Vr/6QULtFRDm6ssbFENawqA15DoYxYeknBStgY6aGSn2BLWsLrqyet71
yXcQzh+uG6PQSHtGDJIASxu+uMTnyoB1ReT+ORWoNEJUqmrQ7/qg6NR737N4MPmORSVwOe3TCeLA
BZbE/6tnOqW24vDUDvRuOPiDu2fKBTvTPPmtlU0w1oj4DyyAiteMvQtTZNQrYL0w30jMLkRSTS44
MbPFct0Z2lLe4qX+DsO2IdZcbkzd6Sde854aQ3l8IRDxz6SHX70HSaiAlCqJK2EdacCudOimCvR0
OCM5u7UcVnakXsTBJMasEzVi6T3axWEVVHmJl6Vw6SiV8ccN83PiaD+cWuvbiAhqwALXviO45ZPx
+0HYKCt9b/vYe/rw5yjykIg5upxKIn5hZV7dCcGUGfR8RlDzdnf3y8vqPDqYzjezY4u6uPVicLlD
xSHgoTpEyaM5WJooaWnZLvaRkjcjSF/HEJYNDR8tJ62MboGadbqVns/V46yP73fBiDpUJopsJzFm
iAzekAGlaIjR4pXVD1Y3JAMwd5dRkfCf+ikjpZD3L3J9EnOPOYB3fbv45TUmo3STL3/v7r5vxvHW
IXnkKqiPpKSsueF/1daVkTOAKHwWJmnG+WxGLNUNTOjFzviBEyNogftws5XwaGeZS39jH15sttP9
yE47pw9tABITLMXP5ne98XArgZMUF0fTqV37Wuo0+lNSKqdVg0+Uvx6mforuFMLoIKGna9jbK2sM
+oF4DrqD0N4zlV4TwG+Ok8mjZEZ6cfcghq0iozGJkS7rBCYQpiy1vcY3fpgLppsoZLiiN+Z/FK0u
mzCDFuV1xXoB/BELuFy8JqQT6Lg3cj3zFtSWXihfcOJkGwrX41UwcaSBm+yisVWAlpTVwD8Xr5ge
Ao1HvnQtL4YqLmOaYPlp+F4D0J1irHh6VA0fnolea/NgiF66cHowvDajWeKmAwDk6wt8h5nWrO6h
sGhRg8AYHnCIQ9NmBPc55KVUM8oPVPo4iRRXCTfkl9rsZweg+Onr7HOmqU+bDXQb9J25qrE4uL/A
my/X2eSzRtP5TyPvkqBRuIfrBRiKBN04eSp7lafpWdiIMGbpUCROvWB07J/D+Z9WNKOFoq9w9nsA
ccFrtMykD3k0w1l8sTD3kgvwrSJB6Uo3QMiR8nYyN9sG8eFboUhzarz048H4dfAKr4uCRYIVqDk+
RY8teKL32jGobwuITUY8GC2q1mtmtxficxYEviS92e/EKqrLTzACi6hHXf2mAhUD5otJ/L6iRmS+
ceEie7gfRM3qkAt6ryqVPl/qWFqOcpAPWP7eoC1OTarkUnkKhnSfP2tNIl+j5iev+nTXYV7M1+Rd
mjHlPZ/ajpe1GgGBmW2H69sa86JorjuDCgpG/oy6tsxLmizfSTyMoMvK8bWEiPdFXtEXqNmJyLb2
FfQXoUvSZGNy5IQ0iHbME6V4pPMW0cevrfrgBBHTakTu/f2plvTh/r40AZCQmX1u/dxZC3avoJch
yVD+olrHEA9UCq7jYnFOJEeFvcsjcxalZ46Xw1LLdD6aMzrAdGgEUw9ArbcAoVPyVoFfh84OqZvC
vEoyX2gXcqMhjyZ49jcbgY4HdGmRAYjqvPFlK95Sk6dqygFc1HcLMOOZd4Wz6qYz9MuKQlKw70pr
9xeuDsHD7Fe4qIt4XKu5+E148cLJMKQUQGdpYzc8vqNriS5Y1uMGpTNt52ygQHAJGf5Mf/XxD581
zc9Eh9EQoBdXvxZ7AeLCHiobPDKOPlFLbsv0q3OZ/p9X7pdGM169TOZBEZBPkLC6kh4tXn3lMXjP
R7N3LavbfxGYXvCn6wqZwxtf1RbwDm5h74V/5zg9gAdcIEVWLc0BFt3hEouJYJkUsm22TSWMFANL
vo47OqY3DD1hRx7Ou41gdNptsloBBxAfjYzArWU+aCq+/rsrwqn9zWZh1rS4AhwIhX0DqVGgnzXw
bmOnsWqfTbeMceAJQTHcc49NJqnksG6Y8JdzPbWZqn20XyecaHWlIJYdd6K/bJTWCvB1taiEcwy3
iXcErdcSjVybgX7D/0ZKUG8Czn8nx9Fn7xPZUCBLcnf+BrB8x5Ufjsh2ydfLM5BE7Qg5lRbGf9e5
TFQjA64xR//lKYx33I/GB5MR9JfT4QOOpBDqfe+Hhpkx9yzRqMW3J8Wd+ACTCalgDmiuhX3rJM6S
lazd3qXcxbWTLpID1huOSsLW+MA1oIFGyl65/GycCAlkx7UurmDMYCHWnxmGsdYJd/5FlrsyXgnX
ZQNm1ujyD0JiMXDYHWzqMkcjjW9UfI8d4yKWD3BoirW8k95tUdGIhiSVhbj7zKXVD0pWhIMpQetR
Yh+lAfsRrC88rHX2OLR+b8339u8Xsk66ZFD9TVrj9MLgZ2qPSp8gB8I+czAOUdPyP0+R+NtfV1wm
Er95HeQKz23n/carwlDngJ4YuFAO1kmcYcjHsayUqMBH5mJGlQyFKwmK7b4jmniCikdmRiALbPCK
G5JhMiHzabAP2+49DsUNVfRNYZrXG/lOU3Kv4oygrxl01Ki2FgiwZohrccYa7tRj467pjinWDPjh
bSLG8Qoab5ApaRU9iKaTxz9AHibZCrTRSeSuer+t+DacU4ik2uNVGi+xJfZ0VdgdZd+wyn69mucX
HNLYj34zHAEIYy9ojArC2FhITn3507vAz6Ior3XoVK6j6IEctUDHQPwZTa4C3oaK7sumIkul3Lx/
DnIYpT+lHQ2yUDzCIX8wTjogBGdk06FGg1rMW/78keqkCoSAh/ktvmGiXDBkKIBnHLxaLDKY2yqK
yPjxkQwCpnmHT/lxHN+1LT+BnofiHo43GwQjrKJwI3uPBYzXB5iqd0HWn8SrLbnLhKjDgod0DfEH
VHxQlMa9d2nYbG3s39klxiAZnBcqodF6TJwlWuPGvyCuxmLmeklKXipIEE3vDhnEqBhhBjDedPfd
NnkepTkm4okwMz3E4aalTTKkghvT5g2fziLU0X3LhtY1ATzIlqn1vqETytq/lfVVXB5ihJilChw/
BJXVrXo+2fUSN8PB5tACGlaYfjomzO2l56VQc32bNpoUEm4fFjp/X8L53c3g300JEmnybgkC74EW
hiD1SAstiZgqJfY0PILjO0r2HVzI+VKRg9ZiUzcQ9k5I3CPLBZcTnKfLnIkFsimsRwgqcKtrfTkc
Ymh7ZXQpD2XO3rXLpY55uqgOhqowUBsINs3shLUos2Lm/yzbKNmg8Byk5EnXx7F8aCCCSp/u3TEq
LNj6X1Riy5wLCK/Q/c//3YATesu/GeqS2XTp8ZFvh7+QFt+Myg5pYgbHAWBKVhlxoLxIP3mIrcG8
ivMAFU3S2SgbIb709LWrPseg47OKPSG/hErn+oQBu2eHDNEciearg+ZqD2OA5ec9HaNLPYGiTq30
BB1X9KSDxF5rRy4RXg8jlqjJ6crKHcuiFPAc4cDxMpSld344vjrlLfi9NppgiP6NoL/ERTKuBy1l
bYb+PTYuB2cOqivzYXz1GGc+EV+cpY+Uv5ETR6fAVGZRLF5W9oojqoCs9BR9F8S8nLMpkuXy3LvI
eZrV1AVkhc5U5nYNmEuA5iH6CDBkQ83lT5FbDLyC13Ky1zNuj5Ig6c3fAguacT01RfmjJlelY8Fc
d/UlxZulvkh8sumYbXdYY5JjATh4e+6Kui1LynSPHi3/m24TaPLeED/Kv66JaI/boUBZMmFfCMZj
wKDhqhvN1GU8x5xpn+JOVn3+MGxnPS9y1v7nwT0uZDf5nsWZ3uv+4v3rPySYZ2+Be6uiVRn7GcgA
WAhv6s+l6PlHb8NUMX5fpUjwZNTFFFz0IUMcU7f/tR+WcA75cDTfTUAmgQOk76OjZ0DXZ0taunGi
uPmwq12JuONASvD/Su61hn+JjdmniClMr/mRWliqLWLo0s8ZrXzraOb6ZMJVuX0E9rEU2W32pjzS
GMvlYBEbzV4fe3NS9cjnXb/AB32MXiYfsX8CU2R5oDHQhLMwxZWErkmBwjTgU9LWceqNE7+8eSAY
tMtcYuumxgoU9B4EgbApRxVMbUQk/adD7yDBKlTQBOtL9CvuOR8EEcFkFSGe51l10ozoKsgNc77L
TqwBF4RKI8LS5VHDn7dPE1tWfpKZ8j/jDBMxi5ybdtcZUVQzEcRfjuYxQ0dPvI+b43ebGWxmcxrS
YcpLkHIG6OTAAeC88FAwxFRHaGlxIFpAqM8VuPzUMYyxl5Oo50DaorNfphzf2s7bzHmyrx0TsAkI
XH5yUpi0Jot3/lxPL+HKExmFW8qGlslqDOk7H8bmCM0njB9lMUfsBKIO2I1X9KuF3JDg3OgFAj+/
wZg/9CXGHxxuHQmLRfGXoT/xdUKYl2h9DExeHrUidGfx2E5y+9THre9LtcvLtPFURbfqagdwaebo
8724vBz2ShxK50pc7KYMohDbcaKrcI5xodXbzRh9qvuOJrkYEEescChf8qQUClBuTLr0GU1hdhUO
/FbD53wc28opFw0jYMnxgTzN4A3fkFP6DwQZ39t47whP7lrQgp5Ur9o5CrYg8J1+Uk3FxiR8q4bZ
rhbHR2GyhFuEibPL0QtGG5tLK4XNB7xcfSgPNVczygJH+EQAQGKnFtOCC1M9/k4k8dWxfeQXAZf5
b25KelDS6AFJunDafJ5dstLBmMch0Jew/exCvxAXsc2JUvxV5oh31te3HgKeGndPivirpnA7wGLB
UxZJrAcoEthhyBzvRnZijuUBy4t5ltcuBDmWJ0IutqHRoQoxTrI6TYsIOJN1T22UVGcGWRAQjDCg
I1MQ4QgzOjE//jIYGOgjCYZLO3WPy2FeavVrPtgeebeJ6eAHtsNF2VwBnaG5UCLxUINHKww0DYw2
RwBEUEtjtg4mr7Q5jyPgmF+gL2Wr/3MBVGVzK3vs/NUn+I5wvkLi0hEd/JRfS4fGiPza7jDwutHU
6cz3O1x4mwGRD6K7DzBKMOZv8zH4NYMQdFaok8YaH6mqytlx9vJ5TIrqtbZmFN3B8+M30XUkp9I1
X5bzyC+8NSX6YyPTpdHNhcCiaEBB47wQmJPTSkc9gvvfSgmsnxnq/aCJuBBJ3zhF5aGHLF2mL0MU
ccZT0ql7DM5LAgWrHI8hf8Mnj+Zda0oJYxhh5t1yaOOtVog2DYqLyXXJ/VQJ0AWKK60mYhiqGKmQ
XGdkKWYzGqczzZpyn0h0Up/PY9pBvSHrVTj5sjzcA3dUbUpJIsiIlk4CqpgI32YrDg5Fb9ZSFTIk
WPQkOge4ZyadD64jKEynGKo/HyMcQWSOj/u/zYHAJg5DcEK7qQ7obUAAq5O7j1Es8F+UNvTzai0L
xzXoHrcopDKoh44PVu0/L3byCUVppFa+0dguEizxRmKfGA51VznW8yhjOYsOuvEbAypRxjpdnFZ3
+KTFm7DSFwEIKXO4weIRPAFLGUyIOSEq7WB9BWuzlK0oq6PPAv3j2ouW0L2m9Oe/UDe12/Pz+1p8
w3emkzPYu/XlP7fgV+6QDs2sXJ497TxcWCls9WYgiyZKV5gL4eSXbvbR4W7+XMjrt9RwGVfwnPye
v2EX4Aw1YtfsI4OvNmxMOlzPQbZ8erGW6V5WXVsOCyec7Z871M3I0PR5H2j+gQt4hUp86YVdv5G1
Xb3gq6OgL7LQG/dxB89awakppBySFQANR/XQiat0n+H8PwkVUWd2yJWtCb/CdWQp8Zn/BBiFNcIT
LjY3OgwP0qKfBqWm8FQxxSMI3IhIiqU9gArNpcC3JquJCVO2fhyP9onajnalXocm7HMo931GOYOR
AcG3uy70Ul583P4ByLnP/fSYuEhhPKce9j3ZWsQJsji32pOSjz+59TTmmHeqOqMXN9Jx/NFF27pW
2YT11CouplMHpJSL2WDR0x2KiUWAxftHkSJWuU/8lB4tzjvcz59OYgTLHd8joM/PPaO+gAxgIymi
9ikxcLoH4//slhkFc1Oiyb97bL/iFLXvkHDXKfyIOMwwAU4fRp+m3hh6vMG0rlwhckAnd5m0IqIO
G7gI9N3vOTQW8tnRdBDO3jBtfvTEQs7OXaxdK87vlC0qJVFBhhPfdyRwagw8hgrgO3pPbwjXPbLR
XpkmsDqfvsuM98CWUF4/uNZU3xBgmIoec/vxg2lxQyF/Gv65B9Uxl0c6QmPURO1UG5XkIPhTpYJr
pIyby42MUZKjnWy3QZlIplsuRKpTc+5xGDt/8DTiUHhqAnsAsqsRv/7/K5j5i1DGBCMSP8vgYtjN
T4qAnhMpv3ZQqoaX1/lDXc4Lw+RXxEXisnENTfDj3K+S4Ykceg/PGPVjNx11dj07QIWW0KOomSOe
ovkd8Ot8YpCi7FTBvx/L6MQBu0Yr3nkcOAN38qfDk1COL/jnK0zXZmoNE2G/lfOhkIwbPurw1GjE
fPPbyqqaoh8k3PMD2UPIw7O7fEH/TFxUBVWQXTAoEyzj1L4KeIEj8nbfBs+bWe9MzK/WLMs8Ixys
FgiQN/ud+cdt6FBsqdZxrw1lq7lO+yu6/5QIlW2JQHAWCBfYPCqskvaW7dlNHa+8GRF6NBVfHR1K
YM37IYgmXV2ympGDNNDiOfob6hG1DTpXDhlapGhbCaPKG23Tvt9hJtgEIV09T+llLU8HUJEvTT2j
6JCELSZFk4OOK+5oudrngI1FbEl+DbTa8nS5yInI3deZvje9c9l2a3DXcUiQC/nk4yUEgP1rRuQN
abuO3wLSkYsUarTOseNSWkNuBIOLeJGExXCpwzyAgJqV+i+MZhurkfuN5RutIWuEuhhaMsJrw1Lg
mOryGbE3RRt+nk7VWkik81BjX9lv+ND70gx66twH9KZSQ0PGyfFTu3eAAHohhCfATVSEVt22HAix
o0+ofM2yoQVVN4Qvh5aoxkHWF9mdQGhw0WqtUs+Mab5XB6ICuBSW65lQcICAB0k6B1Tq9rHWqEqI
C0zUf/mjEDurEGDsmf2AOz9T86EpO5RoKYGD4EmflqGx1+XJ5VfELQ4iHl5dNl577/rMrs6U0EPM
8W6Qi3tzb/zPf9swCO02+2/zRacxsLZFEMHw3gKQZ1PIjg/PHi7FJEeSa1wIEXQXNYbMwm7LaS5d
LQYG8Z6LwG3THd6Od4qBcgG6g1LYfbUg+h0YQIBFjc6Ay6HPVZ4rkTAukvLm9AOnTd3TOF4MiYCP
wI/T6JcrEIuSozSUlU3JAkrJTZyzKxPTx1ju2NJAZP7CwDkoKAtm4PcSq7fQXfDoSKoDTp7bkQKR
Jnapi7ya9CIeMMLoHMiYFd3QK+1RWsG1BaRBcT6tSIFnPz0DcNJKyEsLDtMH+geVmzM5yNwEOP93
YDxX0vKWZUKKmt1mtNA3jIOs/5FO7HlPg+BTwVZze0TB+TxA9mJSPp28UIr+xM8wG7BHaDmbVziF
lPznbaJZuzK3wAaxLksqSofj3yxbTFM77ZIEWnXQM4n0t5vkCNilmvto103OZm4pEynPrST68YC9
MmWs0sjkys6WaIXUVTNw4nFtHcLfdTfNiYlnN78F8It8mzIBQAs9u1qckrZeMHcOmf8O7HJCYjXN
1CkIDfgxsl6P3FfmmuqKiDJE7KNwQIoWMQEoVYR8Ry2gWtBfl+Jx8DL/kmyiIdISuYx3kBCiVqgN
ayiMSAZsX2QxyOisF2Pc088kUSZQBpsGWYQVzwuQaJhA4yHzbSMU6yHV3ME85zpdUmeDJhh6jaw+
dRHh0CX5/+VhRog+aUwKBfcCh70qc5W3XZclkidsOpF0kNDgY7MVzIePj7GaJD7TkKN5k+HFRHDV
Fuy1JPfOl89PIaDbTYuoWqJ2HZlmyyfn2sYE+FAuNNZRLOaYOeSr7YnJoT71cVU6PPh87hqaM0IT
ZxJOPntRfdy5FIw8F0gN5hZ0qiJz7SVQN5G6IVw2wteXDH/OS84U3AGHMyVFdd9NlppkIm7c/DS8
Uqv3d2T7/Ww6wXTgUznA/C2vKigBdPnpIj6v/bEnx5v+D+eSfpwCkw1WbIfIy0dA78EtMR5ASYgl
Qxmy00QLisoX6BrXk4vJOxo8AbwzEXGfxa0ZVJDGHiT8I7lJllqEN2731kgeCyDFfUE+3F5QhzIm
0+pTIc2KkoVgIKxDMov/QxYLgj2oUw1TXRr2VrbPbzu1/246yRmACRYm4xoxvAvj3kzbNkrO+q9R
DOVTMqW00+Oo7eSTDcsWW+EvaJ56gSrfI97fAdMKkS+0U65N0QeNvJlWPA8A6gb1/wVQN0WdZKO9
N9xM5+9Fztt91ne0B17pLiPtI/QNd7u6VEOSXgsgF/9Vwu4sN10B6MzLkxuZyKd5/BZQy+t+mWl/
e4TIoXFsRwEqG/XykfLmbWQQ4zTr6ExyaQJRF2IUOiU+vzemaWtul3GwoOoXp0b1kg7aZZeNKkq+
xda3RkAb9MHxniL3ujnm+d5YYjJsxm/BBNBnp8IWvPh2Gyt4qXxrr8JQ+bIDvNRuYjvUppmQ9fR1
oI6eGlXMcPVUEjN4ftzC/42u174B3X7VrMjob/BqLimSsNgD5Q1y1Lc7N5IAA9CsNJoMTPPRHV70
kn85RBVIVT+DYK4gP11ivEPsXMetFeBKpl25c4ZkShuMqDAWKPBy4jPvvQvhtdXjXpONO+fO2M+D
uOeYlOAZ9DDPlcMBT63DabEETUYoo/bz63XJ0f+rDa/+yw371JdIrsPNoBfIFNocFEc1ykVyN5Wq
HUlLc+UvBVLmhAc/Kkd1k88iIyTIM5qjBZSEWMXjaRxZm99L/kcaF2PAgAoCE8B0JYBCpV/3jMeB
N5TurN/trBUNxOD/uOYNiufyXQSaiFOIpXgYYpzzjCT0I1UhQA4QIzO7NbtHA0mtckIlkflUsl2c
O/WwxPQT5mLuLyeFj22jSxv1hX7B2oipAF+9qqH8IVSd6DApr81gA7VNI8xEF7eTp01K0PIoWLf6
2QUkKuKUiC/Q0p3NmxycjkpcI8ZypRH20VDDmtCMm+XS+pmiwH9rEwXbmJNZ/fJyx9H+zNDL2+4K
XzhPKSJayZRDc/P1QPlIvTH9YJvyUkDZANeHbZDLOSHtGhIjWDLU+JuRUhSzPbA4xyfNbm1MTohJ
OndSlKYcBinHoj6errgD5wfmk8+VL7TcwUUYWOC3NIhK9jyKBLKY79+HLPEV3jHjEbalSmWOWTqp
kQq2/oZnOZdw6Jgq+EuCHtEwjUbQrJFKeIt8BWv69GvA4M25LP6adIb/Ij2UqMdP+zzyNede2En1
AraVLEocImXCfr/i7zkIVYNI7klfC8/QA81GK89mlhZ9s0fS2oV/Kovh9x6H61jv1pOvqFBcMOxx
NmL6CZN8FD5cqs0BBknjxfBiu6PzTv5zzgUjyvc/Pbkm+GscsuuyEM+Dd1Ow1KxXSCAQFd/fhzwT
QuejIaNeRrNysHp+qggQAqsB7xqK0uCmJBMjQ9/od9urhDOjZau/atVaFaZe1Jz0/GoLARFwdfg7
hWzyr/7s8/5hwwpc4bhFoCyp3RLgWoycuYl2luB+sP/px7n26msB8S4r50+qP/Klq++jzIzXhIAZ
PRRxBxtBXXc4ncOfQf6yT+t/IN2xhdmNkUN1A7zLRL73OprlYkWmfJiKanesbUwv5pByXt5Pvcl1
Y8BzuIZORWFj5YuKzzPVjaU95p8Y27qoDPcPCiKY2qpQr8ihHVIMAVM5FW4IgjIK6yqu6vcqbtuK
TcBq9DeCYUDbDXv+0Kl7Gi2Om4GTp/+jNrKEiOihwncfV7Hnx+dmBvBZgcsfVZftpOhqHMjIK5Rr
MzPQx7cA4t8H6fyhqz37MSUyKd7izY0upksREWcokZpCtACQBtQSbp01NOQ4Kia1HBpMjD92hNuM
nordrNOgY8aL0bwcFfS87OddXNm/sX4S2w9bn89mWKQ/ZaP+TLuJDcUWXNds9ob/E7rqznSXUGWB
T3Z75GZbQh9B6fL+ydwkSRnJ3UBvWrKPReypYIAA+1A7BzkL+8IeuahTyKjoIDBA5FwpLz/I4irw
DYJzdbQsJC9YKpMZ8oZGA0SoErm8k2oPsBGhbojcs+jSe7cnv9wOg/XlfKgrzlrYKkr/qZkPJIEa
KO0mXIKE6DNJ1lQgECGvwKwjZyHFE1WfKc8sldx+k0qoanvVyaiYOjG4ynqj2kz0NDvXdQbijDtx
gG3O+L0JmUjJIcjRcy6lh92oirYRmOE4BCs3mWE85BoOoSwkQR4maG4sy8C/08zG5oJbRo4F3p07
7kradcgSP8PF1jqhZk4PMbzccZpoU5Lxu3NOjZCzwVFcH3I4oBR1QltizZ0aN17IsoUod8n3vwgF
WNfZ4H2eLksis4dU0eTPYkV10YTN7IL7pwOe6AeBjig2HPiLh9tEWqyckGUYYwwfaTxPFiS4sJTg
YpYUcjlZTraqw8/4iUS0JLXUNguncudlLE1Kxv5WBBaKpXe288ITPF2fHypVqWUy44sKjtS7zk9t
D8HJNwQ9Q25CZXk8VYcLftuXdY2bbQiPa8Hd2B5VJqmF9S3WEDukT3DcUG7/I/LQRVAqGe6SBcxR
jaZ1Fbo99wmeVLKDuInnsrTz8B5Ltg0zdHz55FrqkBEqaz8rP494EtOt7JtGVzI8Nioregs3OTfj
Fj8SPlKrDWWjnCeCMjykijgtuB5yoRtcIU/a31d2LcGGM6VsYJ52NMHnD90EXKtcwT7v9URtCZRV
VaXHCBh4BV0Bko+p+yxkmXBfIs7lfyfEI2AyYlKxgmoybYpRxsP17r9ms52hjw5entxb0abaoMOR
MpDRG+O9ECoYsMDDHVpkEmYqrm1KKMN6/doeR2iFg559DxfLpH51Th3Lx4fcTXaolcbYPzkuyI6e
QHmzO7/L4KYU++jb1AmXN756G3hU/+3rkwfAD0M4j22lVsgz+4boFXPpCZn9QT7qY5TFbmw9unUz
L+9v3tjSb9dw6ANseMhZBESZbeXjrnWSDgSfRTEiApvtHmdLACXQmW7l0/ZMH3/fodV0c9NmZ6Dz
pE9+9ceUT1YmuHGrnbQIkQHnMr/i3CWB3cvWO5Rl9VpTSEMIZGOEC1qWg2kGndtiHe9od1kOLrKW
DTWFSAmSQZbekU8aZGtOf+D29cMNK3SiD+2hJWCG7Bb+UYxrDB/dPEBYRdhVHXj8nxQDVpa2jYn2
rlxoOFb9MDfwGup+jqftwutZ1oRnMn0gK+zZVJPgEf4Qbq2wGwq7+mK3Rc9vdkqfKTXh991i6YJR
V5UnqH3k/lec5rdF8rKIUltSHTmYuMcTLUNdcCz5vYjdl/t/GDX3SozNw4n4w4j90fnOtDxAn0s+
VE/fZfBGiQgoIAIR0XJRGfutw9FIOW0OwHbMKD4fGA7Q8aSyi2PBzm2EOVQGZ7ZlGh1PkYHCa2W2
Ro8IQYCmiQx4FsEAaWMxBCigAyRN+Zae+YMYPc7lxkBVc7zYsIgcwR72xjc2WjYrEVaLsBs3kBCL
2snF+l1s8Y++9ArmTvb4sBT1s1RGfwj4g5T4hqJ/UhwM439Vs/kKcDgZHNAEjqUuimQvKTVTCAUn
C65wCCi82ROXlWRoqKsGGICMNV75PCBQOvHwVLT8Pi/5PlKUfbbVUBFSKIIC4rY6wXVW9gU37Y1I
BcrkfW/gv1TgIJNMvM742FL7RXS4bYS7YqDhg1vn2XOX/Za83r+5tcLoXpl7eNmjG0gdzIjqN8pG
cWxxA7P2a8SpjmN9hzqkCf6qwIrHBt578JB7mpVNI1H9xoTeV1N6g2oBdFNygGjI53RDxPWPyv7h
pghjWuZnhc32px20Yfdo7PZV3/pUKPYbznlKuV4m2XCP2DsUkTF25opq+Tnc6Klk3/Tx9G5oc5yJ
2OrlsZy22gwYCv1VuzjP0JeD3dMTowy4cqZwcXROwTYYgzCY/K3OQFg2mFdmWR3RIIVV2GZpLOzd
C33YSFuHe1OB0+KWVuRQ4HaNwvzf9K1YUj2EmpXA34OUO23XuVvtLrKm7vRVU/KbTzhIRFzFkBO6
3hnMCsEv9uSUrpI8CE14z6XzqojdPbvEHnlqIXA/o6heSKUbZiZ+Af/JFTaujQK86EkniF90JUux
jtlQZIqPZKAThdQIaTLVGxTKXjpfONzDenXDcAo3eImEurDlm5k7Pc0s8MrabpR2Tw4pae7C4ct2
lSXUmIzRnzF7DVQEVZGlIqGGhOJU6yMIifzVrxrPdA6FZX2hdiyZjfJXkyZZGSngQS+A9ObbipVh
MLEOpJsJHC+LfX45rJasfKLmCqRdJevW5dx6n+0NxA7KzqbrxvqkGEJ6wvfLuAU/PShlYtBp/32m
9tLji0fq0FD6dXNnhnyvujCITgi5WGqR5OYCsYIQiLtu+o4eDrwNAc/mPjZMLen6kK2CxPzPRcoV
s4unSzgu7bXk+vmF2rD05eGVJhNtW8nCLQlSgxDyKjMRjzFxDgtsywM/6cp6bD2DeF1v3zCdu7St
zC3Ghy1+Wl+MBXf0V11xj7Fj7Z3afSZej8Ilgtx3LbYf/BHqHBliZNDVNmRyVoatpyXI6MCSKsU0
nnjslxto9buD+7UhKHcx7mUcxkeNNWdT3UuXJtDAVMwKf9mQ6PeRHEoowMFyVuyOpRLbNnuuqe5Y
/fk6RFEi05h66+YWsKBDmX6GpZWP1mwTZBVZ3as6UPDx5fSrppmH8+i171Q3sF3G6f1CfeZz8iUE
O0KoCYPrwpAiiH+zusXZ4cCBAKU9U8bx+vc+EoXacHl+fAHSwTqlQ/dCp2TsynWOIOBAoFFo8j03
uatsE/zz0zThT9kHHKf70VeAmSQcSceU8upH2DhXbSZ5ol1G4KOlNO4hbsOER3TxcgY2d7b4/pPt
jaC8o8ulLUiC1y7VBNSYCzwjMMfV9IbwswQ9JiMdqrtTOjjKpzueX0wYJ1oWyLNiWCTPzDpZOuwN
d8lamobJhLITOtXmhOqLxZpc/M2QQ2yWY0oI6nmj/cVYt4LGbbfu3ep8r/HxO4SUKQYDXsJ/lG//
6h8jK6lhGKSz6nRgkqgVJBdrCmlctaEXNRMI/Z9Z/ytFZzspU/xMUO1ACIGFCn/6XGd4xZn4/MKd
fppJfAELds91YVBYEV3boeKl6DrUzxmn7DPDaZ1OhS2ryvKpUo3v17EF+ts2i7+VjuwzHP28MgmX
YRYLnCIirzI5yPVLSpRjvCpeP9SRvoqposhnLLROX2t3IUkaaRSJdJWQ5DJ1Nv5hdaN+w0G+wh5C
mNdB/3AiDd7b56TxLDewQM5W+XMQXIDGq1ljx97kDpxUs6nxOJ4wMdE6u8211VPk1npnJxyNtOed
KoK6XuGPhvXuJ5eP/8FmUp5UXgcjdJw+xsH9p09h+V7OEU+qrI6IsJycLGgPA42UvmExt6cyx7Wz
2kysBGRfWaNWYHK9uNVlLEq3NPQB0nfS15zt41MMsNW80tiLFmE7ZpNr5JWsa5AkoU9q273FCsuw
tb1chkK22V4MCa47JHlxHgnivz1WrCVGRj4D243givGLVWEn3tjJTIe4oTpsH8weJPfPtBSORgl8
Wa9YQbBz/65mFaEAZmStf2OkHKyEe00OqYsF1kl5XMwtUU7yOykwzfTt2kYk6mjQPVRZ6hHF/2ij
DV/HfdwKQr6tFoXfvymcYhJW98jaiFGLXj6QeXg1rOZh50g6/CQkR0RqZ6u2h3nNGqXcFBfR9GFU
3Z0vAPF8y4vdrjVZiWK1FPrRM8w79/Rvi0Isy21MM39fkusB0iehKn8x3bowVwPS91T3lP0xRAz1
MFd0VQnuqq6GtNnqZB21KFc4XFaDc3A75gbcyZ4HFzz8yE6ey5oncnHsZ2C1niPMKSGujglLVwm8
RSyz0KbQbCOPbRH++g7wjTo8RznWSf4Tdk2yhDOJk9LRHLO2CMu/V0fd/i51rfzBc3UV4U62lfum
BOOdoWSL4d7MINNDlUdOqrrDRIqBgswaooDpV2yCZs4nljBtVsYOLuJkFg3QggmRfp/188wsn4LW
B2Qp/M2JD4HvzJiC2MUxkLUpaFjtRmCT3PILl1uK1EBpj0EsVTepCLuTDJXC1aClVQqwgrQxs/Fy
KecgOIMbmQ7hUrotE9PzIoTheDTwsnOAO/If08Y0x05XindlbVXx/FDT+Mk6pmXsFe0fP2WdxLKS
Adzz0eQaH0YG9W2NfGG4K1g1XyMEkvRV+PMLkfpip49/ckkiS+WkOOAppGawkswyTYObnnyScKf9
Z4OVtJcNHgRgZi8uA/M12HSnCRMEbDfqFTSMF8ozJN5FwwaN/XFvTEUgXqT1y4chR0hX4b7g1Hd2
SJrH2Oh7HF8WvAP1us52EbobcwBZTO2NoxgqM+1Qt0UXBX5OHdi2YDAMEPddv8Z3DUyLdRKkhi0X
ORKVx4kr/p08/7jmS4FSSWTcmCQi6KAEjqvmgoQMxOidspXFzkdxhUoyi24j97hsgCiYq9USzi2M
aiLqJxaGPybcCb0Pkk2GfPlBZuc16EqXlwftf2LlmbuWw1sAjE7KW69dMxbrg+7vZSxFgfolBiPX
CouYLjDdaCs9mm0UNTrOUB6ZBXxe8976o6u7Jt6T+phTO6yY5zv4ZA2Gbwwp4GJN/7iYSVUpGy6S
K/eLoiWOcpcH4DdWUyFiRLwpGm9YAyC0VOs4s6wrHvEjlkeM5bAspJgIWX/7Nj6+3JQoXD8E0GGk
cMTCE0QG2UADTQzlzTUsooZ2wIe9C5ZwZA3fKNboHv84blaXRcbhMUo1BFiHdpjHgDuPx7wWgDcW
UJKblvH+sdC3oDly0ZElqq2FjCu2UXQ4vQ9M2ZtUToCxIrLul3PSu+ycoXT7AKrAh/uEbbzbhd/z
uaUVH/8h9OLkavut2ur5yFN15dOWiREMR0WFR3oM2lTlOK0TMAr0sb5fcu/RffTQdhW/vFAnS1/T
ucicI5SH9QEUuy7pkdeqh4ggyn1xzqa8WyVeme+P7aESYhEznjkIHJMJzLaHaF0pViygHqQ35FQp
ul4BN/FuLeXABrntZu0QLvuIM3uYtznSxHjTmAfLEFarkk6Vmpfc3hUQrzM2B4sx4J+eqzU4jmFo
o0YvGtkTWcS8Xah4sIWbzylXLwv++lCzQYiM1bGjMT3iQdCaw2IrakVZWK5R2CJqQK4PgWjC5Pmm
deEysnwwunwDMUrl76IF55uppyYOPrE4YlA4Uk/NUApFt0Mjxq3Q5i4TNIK8kBnxbB+I4HifTL1s
qeehhFA5MYUs2ptTK6akm95tK61KRo4F7GkFWulXka/0cJlr9ceS9Xxm7GqdLcr+vh2t7bdQlnwV
avoD8WlIP72hYXcI4SUECpK0ntdRkgvcOVJE4fAk1aMUcSx9ZoF7Cg83x+jsQcAfaMAbhI5QW/v7
aQy2biadmMTTHfmynoz6fgqOIs65uVJ+Byr5TePmZuDEUbPJbOnd2upwRb6tc7HOrfXbU73WX7s9
+NSpaBXvfEy3vF8mcrGvoazHnTZupiEtfDaOBP1GmVczOOSxaXN2RtWwAgDR5fObGPNOK3YxwTIN
3wxxRLc443f8HAJI8MnJP8W+vsjRxLD4oQsARqEHl/0xWxl1Yx1vfMgS+Mfe2p+LaBbiULgZTvN7
FEZ2/PpgLanIwHiyg/yWZ8OWfa38V/K8dle3jDoKdlblazZCpoZAv8clH6818brM59VBQfQkxNaI
EANFkYV18sPE+JlHC9QkCK4jt9IRMXsAU9SWvVwZismjPouD9RyzaXnPfTpFBSLnMXfGoahgreya
54y4caJQWoQukSazqO17+q5VcqVCN9TACnB28H4T3473Gm/EaRt0DfCNu7izNet9Hdgr2eY8WDQt
2EqpStbczGU7FtJxtMHeqGjEkfqRsI07EYJ/Hg9f23SUOIrHUa++lLfzxFjePbQCwkqB3gX4jqZb
qJJdj+hiBsLYvZJOKe1mpdOtnlaVJBbSvGm+YKPhR4t7A/BA3KBqg3Vuib3vyfwdAj6E5pvCKarj
y7cizX0u28GrC0sAtXehJ9yjfC4eF205R0qFdWiPfXz2zAbl0gc1MkSuVpt4sr5ROPl9tiR3WhGd
UEtc0Cw9mMiyqr5Dp5vos/FXm+Dt8iBMU2sUsYmMzDZn64xsgTaNg50e2AN/Y4vvLY4ss+QWQ037
UBzGbkco4OeGhred5pD88eG5Ug9Q+OqiQKjaNVC10WVTeQRhCynzm8tJMXloUshvZ98TAELaVYsn
GhBMqRU+Ooj30iI14TtzHEHxDfeKEDwllH19QlQZVkcNh5eFDiYfK4HTngB8zoxdvDotBLTr7yeK
gHtR5dStZdaaxo2X6vDEa19F6VvCzO2+gRG7cOYFzv8EBh90GDXOkb+n2T3SYSMrTnIg0M1RX+rK
NxHgiothAPLdUtTeuORCG0esvOPkNMxaQiRsenAwLLKRTdYqLtXe5M83N+H1yoLsuTdv+ti3qroo
w4aIYF77NlZ973Dvq/o3Zyq/mGNPLloow1XP+frC74cEqWy5Ne9LUs1N98hpuQ7FmkCVL2bZeMVO
J2OTtmgLdKuCvHlB4fFI85J8G+lI6zxGAcjhr1YLGVnB7lKNRtDoqoa/xK13XdIjrC8cR5NApkFt
XxJvbOZy6aoCbPDv0KZ9t+lwaUEuRWC6qPjqzhVK/2XWcJmAOkLTEjLahDqa2wplLEojpyWNTzoL
/PNTGJ3O54SIWvczjQhKALbxrIjsOni1NTFA37Y2VOFeKosHhR2pZeDsII1vZtPtiRBI4eFlcoKh
N9ijLeuPB969VICfrcwzHZkQp278Fy3YWQHcCw2977wWsy6hrf8T2C2UXQi6fWy2dEuBYIspLKVP
Gap4H1Hi0TG3jT2WZwhrYHDq/j+apnAoyaf1VGQZOEluKyu6mwKpM3PTVIXKmxferhjK8uOMlP7U
+IR9TgqSEHm8wCTzXw2gC2nXX3b2+bp3jmA42QYQJ2icHx7f1dphZ+MZ/RygzyOODwFSwG0+T2Eu
wWIDwCV/ARxRx2OUuybpQ9GEITvNzFTpncM615CKGcriU2LwMK4wHiQiXyVFZKUsNi7xAAT5v3X2
FWuujw3AbY1ZSeS6Y9NK22qEp8ia7td5g5ZH69fCZyOynRI0k/eDbEDvTXA0Crxxwuv7VpXMeGKa
7SudQ7L12rmIlBvaF+ej5JTj/CVBmdBB6HenjvO1eR0SUmUehcIVJPgyBQe98EyJROf7ZD270AYc
/ugNYE1rdTXukUcenLhMUgaSemV1YRlvz3qPSoK8kaPq2hwRmeG/BAtLI7DbLuVZst8tRIBZt6B7
EIB6BM//9IWxYH3qmi0XWycqpj65QuwnzJOkHdt8qf73YOm0fNKPL6cY8iujKCN7iOK1kLcwszcu
2hy2OtgurGJi/5WXVG4HvI532VhdwfO9ZJUxvgsR/EH/LrgL874aq044xHe/O11HjXDKM8Krcs1j
BiBvqbBuEXaLr9AH3eJv4RsvUyKneNkWV+hicuYki27yWcEYLaDyouYDxBvVWp+uQfmqLORr8504
WKd0T/0pA0nLrSxJnAKe7EWS1KfGyQFP2ThPDOWZ/YiaVJec2aKbFocSrYxMIvVAsOMSnvxwhRss
9PcWIKkphktZFTnH4pdG580mkQz3rInk7w5ExOmm/PHlVzSiYCmr4y9XXdY+zvBGfiBsjg07vBb9
ugz9XQtGsALUx0MavWVMIUI94aVyDEngv9nFiPr9hI+eV69gnY0yLpKyyuIUKP0xEIz1OfqmmuyH
YxSes0P4XykfEiE/dpFDOJ22GtDdQv03emigNpU5E2HGTFOdl2OppBa6WFuQKAprAxaHJR6NP8Jv
AWkJDcgxoAjhOs2FSOt84aRTqnMHPGc9i5BR+BCu4RqMsaJxhpkHAdp+AqjF1U5gufvokZt1hIFa
q7cRu9kwdCMItHyfCID0o+YIlS9Z1EzKvLuJk8RAkXCnaiac7MDD1labZ7DvzC++U69EN/K6WRoJ
q9zTfHmdOpnX9U+jizMm5UC/OhtTA0b9jWFFV9B0rB1uIPHYvYR3chgx1s/d2SELAbJ5FQiAEvn7
c2VtWVAyXG8v/mrjAvyG/nt2LWqxLSdRL7fD2H29u1MV1S20rpTUv/BhV5D7ZDFvDoPdy8UDPQ6u
y5aeFAxG9o/p+l2Y2b9rP2ymi18lFo4YN/JEw7sTcic0DB+Kmgq2LuUjLOtyVWkoTNninjjnOKCp
yFsXCPHeN00/8um31PEsUYCPWGDL9igzR4840N6MRrwfNp0QrwYwlxoubqb8hDJnLI9gnK/JeHxh
3nf1ynFmhxtD/KmteaNQle5nQraKcfvjbclz1Jjjz66awWAQgk+t/6HrFUvQCUATIaer9Wpo+k+f
TC/Nlu4B/DA/o6Y38jHiChOnI1ieg1PHjFgnA/EnPBoWB/Dss/cisC+ufGIeKjTcUhcY8+8pdJ3H
+pjVZ714o5U10a0EdctKwY2HS4HrOITPiFqTmWiQP31F/dqrYP0S+O7MiBdV60Ez5jfo4aXYroXV
25FbwH0G9ah+O06GoNdR/2J0IeIHplkhfirN8TsYWbiSr0nJjrIiYcEQ3c0QxBl0WOqXRiW3FNGq
vJx18j4FA8//fwCtTzj9UKDXR3ObPwr8PyfzTtUZq27Lb1x+sojOB3vYkoA+GguBN/jxQgodPWuB
mOYfOjdhbhIh7DIQwnb4f0R9c/60bYhlk5DZEdWJ6Xnn2LxxVfC2xMGsvFrylZzvjQOTE8SzKIev
IHkHdGqiQmGOie06SCXcr8SQ/1bijdx7Hi20AJexasBScIY5ypJDa+6m7+mqEo7L6oHWsB2hBUi0
oHXCn0OO9VgwO3/IcqVPq3U+rRJyqNjMJji7wJMt36yzX0t3J89s1JC8n0ldSiAvN6yAoDoGK2Ed
a6Jj/6wjprjB9b6z+icmeTMotjQ6Zv8nfrFPKLUzc89sSgEN9Q632OYN+0FADMpnEhPCQEukW3xy
iexuSMha7lsF1Q8eqhEDUGXu5FQQu0WBcpFxbCsQnJ0D2FqOUxVkrsV+WRDH81BDlbknFRT+sdId
HnGaauSJ5XIZOekbSjIxrEtHPsFI1zLjNpmzbnTMYpi6qBDy3xO68D2LUfisigU2T+0yoSPeapPW
FkQwm/G2M/35VaTYyqmOVV4f2MrvK4zSHnSvzrk55IxOIxn0SROukEYG4pGDR/cymtz9dTGoSOmz
JdnE5vCI46a1vQcf9gRg6FdStZWVARn4Z80HBpB290nZcIXnK2Ya9w75ZpCEI34h6IjAIb9l4I+T
MgxmoRvDezuDYILNjR+aSIACgrZDTAASIN5+wr+CqaQEQuFdP7jc7nZ8O56Q911fMw6lYb1CJPGp
JwxMbuMGVWW6EMsiYZpGN1i6pkrQPGlo7+L6EC7Q7ZmroMor1E67Z1RCfFYYTwgrcXKP/kQ83q81
5kcoTCeb4dOM9qdzZ3ltmhD/vriURVzu4VH/AumTlzx6Zsl9YcjAxsdprM6bIcA5UD94Z9xv8KE2
tc26/2OUsQpXivHqq+LGtdGIxR6qm9Aaul2FxeBp2M0vHRP51jqJoWxMrysOcUqxry9B6CBI7C9N
DAX7evuf4hVqJPhBRbF++qGTV/r1xYrd91iYxMej5NdefoFeMxdE+WFLfRqgG757IZ2k1QgzVg/I
N95AYPIn0jntcPvdy5vKpDDaFU5dKKZNKAZso4m4ynUgm7EITV74vMrSe3jmMBnBpBRI+QpOO7YO
ZBGdWdjF0vvu+YCljtQJXwVCLYCO7Zhyn/9MPYfzdlIcIJfX7aVbTRDUAlPgPMnsYm1A42zrtKAs
TpdWFBMOh1H6fexRjFcJ2QmJQpPapUht9xEblmceyx+DbYI0kXtgYhXwGtDjAsI2HYOzS7E+MKhR
lEqBPhOMuBKxNzAHyWQPp5ZpCRigeSDbLvdBo1YmCRRHIhqUgzWTkJdc/hZCapxUpN/kgHDcoPVe
axq4QFCTD2tDWkX9n4p9lBkfGTvaNh7M49JUYN2i4g7JS7yAI7QTLzGhf5OcI6xhnfFXfLx66Tll
KaBZ1TbBct10UjaT4nRBiox0T70UQBySqGUTHJX/unB3eEpPLMz7hO+thv0KbCGi8C4F4GzW54eW
kXth1TfFXN6khmTWtdjSB+ocmlKb3RVQOmrMTPZWzSq87gqtFp4N5zg0py2Wxfbh4VoqDHQL/w5L
3iP22rnO9OXhUIPF2TlUzp+3R+qDsa7oRPCo0pIQWhmwIFcWXzL1G7f7nlYQdS0Cav+29mgozL0s
P6PWeeW1uJb5fydJ0SbYpKcAKq6HO4lp80dTbEIUUOH0aTFElcVw6mYUf/95cB7MQ2AoHkX0QXOk
bbvXVu5YfqWStvNvzsflY5B6ljoNMGBbfzvfqXgxl9JArimOBsoMYDVHbaX0y358oCYvLMa3yMyi
1Ej/OROM1Q8fKbKjQbZpMU1CoWV/NemvsfGLNJ+RZp43CWhmuxpLDcTR8cPU42FkBjK1l2AEM2zW
oIxEasjNmRD8I4DMWCVIWOlx71cKsheU89C6YZDD0Clx7dUcEVLlxfvKtJEx3gu3miSFy2DpmCWf
0dy5yBzaEfq5WReLricDPPSt5Ql4ROP7dw0f18UuuNhTFEqtQOHmlc3qT1kPoARkWOSy7g7e2tRk
gq/nDTWmj9FLF2vxp615Zxw/rXWqa9q8u6088GxOMpt8gakXgkWMY1w2Nh2oFWARjZ6anx5Eva3y
2D8YpaRDg2uDChWlknTUQqNDx5T78RfEO6luJd37kZd0F/KR6OBMRkNklMCqohwOSsRhyCZuGILa
OkCeJZOm/AqKGOEJ/XXpfAS6mI3RuiOaaQM7Xx23uCQl/aGFGR8HgjfSIoIwB6gq3iesb3eNNixx
KpBmGnielSS1vVHjcD55cp6UHRVci2OsC7U8bMLPuHJVhA/aiUk8PpjCrQApN8i1n33lUdMBhROL
GR4nXSQoscsnuvoOgpTCKZF2cEPgkDw8KwhqW9SYd4KhErYiRUyWYQAn1jwy3DgH+4TjsXDvFtXu
TBtp3QoPz0dY5jFAF+4jlvYoCyidZGfnkZ7lfUxBe8dGMoYIElfMBMh3mvdmgHuvqkbhyezrm/UY
nvT31TgpozoT0DxwOttHdaOFDwni+8vUh/cPz1sXZGqqAJXKnsL67YuRoOIN543u5sST0o//Pc5N
M71e4M098trdOA3OCjWFNaB8+vbZREKV2IIwWRNAb6q66czjlgi8YAhNZ7g75fTTiYkyQI6BkSmA
WnazYpIllZcAyxUpPtRGRapGcqWbO4eGn+ZzLOY8tzEqLP/SmH/HKT1M1KUZELtIZD7vBmVYPe0+
NgX38cnJSL4WDGOP3oOdDHnNtYiCgjtJvLDiBcq+5h+h+Y4sAVNkLFu9pkNiSI9ivjzyvYFYpvo1
LnloMf5qIrECVEVmXeW3veVLes/E4TV9hpC5iXI82FVX6VXeU76O93ZBDf+qKFR3GHyUvWLtrJOA
qK7vMiVZzZX1OtrSP9q5ThRaMlFf245e3XGg/COUMc9q/SOPSCNAKdFVJZzl8Hlz07y0t/BAOSLj
sppxNwJoYNzBPvcL4hYdqMp93qQmpw317KmiLXbIGI6AuN++Yfc9tpOcOtFSfPQlTnEUmgQkaCIU
KS2dH8bdQk0k32nGkCDCI4b/kdy5+rqVmtrBWnGVjCpruwOsqCowSUaePKPN3pjT7gMoEEQRWUfx
h2B1pEUQlvIciqh/ZTfAZ3ucbxOPzJ6CxGkD9+Dup1B6EIe41TxjXEBnBxgREJIyuP1WIzgttpwT
79a8yD2rZubbjymHQ7spr5uRsPFkj5DpKR0qA+puIigy1FszU+Xgy7e6q8LCpAOSmAyzqmtphBsJ
cgcJA8gTiywkr2+KieG0DC8Uo3qdlDRbZfNHDvSmZDygAk1uVVU6mAM0ZYVrgKa1C7iI+MZaYyky
E7b5ixQS2NZKeOb0a7Q4j9EBVlLM1S4eGfZE5ew+fU1aVqiSV52ymioRc2YvcfiNNXu5M5g3TQiF
Ff7K6uygVzWz0htzxaJuBH9WebrtdA8iLdiK8IXgfgWliDQRakmGwAGod5loXDixVhCpB+xjCcSp
GCNNgDdvABkAjyhWSkcK4/7qSeQitgjqdQ9VTG9w3EBRVaB65dGVu/8GGBlAQeIR2o69aD+vC/N3
JBF3LwrXYGl23Sgbaa0J3ImyThatP7CrprG34U/SoDnw/8VK2lmEridUGe5EaKbC7y32CgaCU//P
8WvygOzQwJIO1IrxIgCuWCJk4gmIXbp4mPwc6I6Wg7P5kPAGY0axYDl3yXIq8y+6FXdQMjD0PTW7
hysMpQk91DNsN8RgauhTzmFh3KzLSsAT1rSgV8fPJ8Kii4/H/fEkk47pMI9/LlD28Zsr85CQNLTe
1x/3qvlEKHwHK2l+RCaqCBF+6LE7vP2XCvKI97GKq5g62OKMVT594MYlAMnU7Bytmn+2+46DGpJY
LvMLHsSmqcngndi+EVv1SwmPJgrCsi/ey5YW5G64DQh1sU7mYR2fL5nB4fm4aO6w/x+zc7mut4zI
iqNakEkz+Fq1iOSNMcSfrNU2HI2UOgaQj2Z07CkGxhNcE2Qo4CxUWQwhW+91aCIfCoSTLpGPcLk+
i0TMwBm0i4XjxRsivwU2HCgkKdUcz6/U91kkHLMjzUIC2+FcyAyJ1GN09rAHWteI3A94jV4sHrVA
/xNB3NOeXUpsAbmAnMBH/0CBOJwVu1gI6KoAvT8VyQklx/5YIsCr57Exf1qudNRu6MTq+NfjIdzx
LATP5GwS4XTm1TdVNvYXIEBlUA+hOSP45BjIAsQd7b9Ep0N9ytXmbFa2htCLTEyjnqrPLX1+Y83F
SLmIkFKA6PxVDFbLU3EAhE+IhXJb9q6fehiIrrqQmadCLl50nvxajszO8jxZacCBYWBTSTkbIvm6
ePWOwbeRW08HUAzRK28aEFnRfMVDr33hgrWmS1RQpO5kUxTuLW0jDperW/bLP4vRbnIGOHk4544Z
3oqIja/xtxPQLLk/IXTFOXIMlJ8OBePQjgscljeNR3I82zVjmhGXMOtwXr5TGyXiXGdO2rP4KJna
sD1UiJ6vPmQKS7qJ5fn6CsiyX8e3N8TE0wcbCPVSqao89x5eQzA87NsWp/d5med/4MT2Skr4b0+p
LXUtqTIpEMRR0nJECx1g5ymdjp/3M1vPZsJGuFIDFGj+eGLK8w5uTLmhpFqsFMi6dNGCWPRDKlTj
PRD8JIiolx4CzSVr2g+F57//qrd8CmB+UAcMoAULBfRGfEMmcpdF0yKftG5Q2DoMdWqiYI2ExVuY
Vw3jbBfVeMJ20SlPVLLjK2++qeYbeHo9HbBu9p7L1wBRKZmDu/quicuXC6+AIaSOOPUQWG34DJii
4geQnM213T4+JB03UpPQQ7+pJQnSjQqW8N1s0oG5UeNYn4Fpcgkm1kXagqkadiHYXcKOD59gPeO3
G83m6u71+MxgZeu4c4ULEhmrdTTG1A0WKkmJNIVrxv6/o6H2GhVbh6HXRG1C/kv1tIdOQjHdAtjl
q7HLUqemRJFI/la20YaqCrYvrhm0PKiVDwy7WXnnhkmI+Skwn/pteA/pQEKmY31794m1Hte3OOIs
VduO9ECWQCqLTJXrJAuwwFUR0L1et0xpdCDWCJkL0MomkFIzRgQe6y4uBcDKQnu45+H8ltoa6OrM
2gqMUVW9oCQ5bZKB/XwBn33zOeMhpc40CZ8H+xPCr/+R14kEN1oM4u6NiVGuxX56Q5GrJCXQ3gbG
zdsCO1cwcXsoPgeIGmz/Got/1o4OxyKMRGSCGEfxVmcYwZPCqFe7oWPd/m3Ap7qM3DMh25/aJ3pU
xq1olwTACuirZsn6bEmoYt3D0b1dEcMfgO0CaaC0qKVkHU8yiB+5Jxkf0DTAhU0AdLHpGfTomntI
acHvUlt+du5VyJ7RDS1dZ38nVA3ktjIdVm9zzB2rok+tQVGQ1XKctlsBwO5Q9ASQa6Olb6UhR8DT
P95MGJ/VGdDwoucA7Zd3ajIFt/UwAW9/Rw1oEvUlvGz3jinnCHr62B680pMh50j4FPIYOI2modqV
XliR4eJ5w5uhhea1Qu81K4Zwid0soFfcnHqbTcTXDfsZO16EcN7RJhdmFZCEulmFBT8kvnJQM6Va
Nq9bGCtdmKB/yNwSMCNhHLyybWGiryLOdQ7KWqDDOtUThJSyyqj+dvh/HvDdWK7OMIHOb8PSiUJp
1U/dTPyhAjb4LVTgAuuKhi/R1F2RjPa19/+n+BTEBxMubg9/nTHvYHR1+rKvirK/qq0z3kS87ayj
iNg3A/ONjIEmxY/zpazo0E0E5ljR/Htl2tQmPMkGxR+3nDFO2pdsIk7lT2KUdM1L5vjwEBoFzOtI
znDuM8ADdH05ZAXUxTyh2Z4HJzxiEn/aLyGwBhFe0tNq1AD/vumS8GUk6KeLV6PMQpJXNkSfrOmI
jyP27+1pXWOhWTHHwUtXDd68k2z49yGezLP4RcxmEzywLT2ZMCIci9GSi556JeI81SZWqYvcYQGb
wcT/tdSai6E48vVtPFjaYcG9EB8yir6/9EBM2ToBMh8KRzrU+xNWVtH4YqsZaLhmffSaMpIznAtN
IFGAMAbQQLxM8tKaPAmW+6tHOfkYfowHJFGoKqe0uibPj42XI1/he2TZ/h2fR8/YlL1JK7iZVF91
4RXAYqNImg8bsWZrF3RO7kfmvhfiuZbc6cOcwdV+XcCiQ8S380FxxnY4XwNjQEumaODtHaEufP8c
ZinkGfmfLqw4axAlvGpooSC3v6wgZy7tG3jWSz73DotlTD0RlrbTadqglPG46uabVJoK2zACgGUf
UzKilel5vHjgq68xTuLkdoiCrtdIJDZteIYrn4VGLKUaAXjYyNt9Hm2wSq7fuQ7g87VnPR+I3wzk
wU4CxjszABPDO/2c3gtwFwBXGnN6w/WGyFcZ3Pwyw83QVuK5TG8cAYH+zYU6vhSWnp5V4/ZICtUh
Nt8FEyXn6AY6IvKYaHHK8d0vfqAHuMebieoiVCzWtzC0Sga7awgXBIWOt++sOwKtZACu6PuYX3d7
8OsoN2IafDQyrUmTiwupX0IcMlhesKiBjc8MDSiRjjZiDOK/gz91R/q/zom4SGgf4hsmq3CLji4S
7utHNNHHLEjZkxa0dL3kaxkiTD4E+QKTp++6eyKj8/cxsGVSVgDNPUdtWGMXws8+jnouU0EYXxdA
WK+2K+IQBZ8CELnqZXb4FoF3OOEgK0QPIKOp5pLlX1nBRNcad6yn2SR3ZOHPt8OSgJS9ZsHdse+P
SAZC44uDAEFH0aiSXpRphrASKqFdl/UrXReqB2rap/yrPH0vLkrhXukAMxaexKN4byzBRgkJIQfP
N7pAzeOKSc9S16aevQKPKWA2JEQqR41yX9G4HO+TJiEt70JSSLE0hX+GiLjc6EwDBeiATvVJsXAG
fgPVI481ClWkELMyE10idSwEdYVNSNJlkA4hfQ3XGN4J6XXqkchRc+9UU2PARwMKjCIdcIKsMHRZ
4OW9lf0asw4+bso3tqzyI0+bw/8G7LQK+9AUiHx93VHPXcOYm7maRCcb1tU/XZegaNQ2HNWMXsod
xPh+BQhG8hNW6TvQ6K1eL6fNlpXquA8v3f/hYAeKjJfHc67k6U+ae6kycjDQr/1k6qjDv7DaI9AM
QpvaqqxIgMzwFHHScD5niEvpgwT1q5jhIhr1w2VAeaFAdiJFTbBavDBTbOJoUpb5K/hH4yXhKadl
k/9fhOOLzeiGO7fQZIbsOYe+bzIxcprYvxqcEab0qmY0wpO41rSCbBGjHlHHWxnwN1NNeTjEJt1f
7nhRdcWnjonpeLizQ5HhVZfx3ikM/fK9Q1Qb4jjTVsxOLvHkqwyx845mKMAp3hriDtcUeLYrhqME
/b6x4Fr7JMG9bcFusnWuCmZ09JThvqTFYTgvqtYHuTxnSMJoIxYrSzOf6eDqCwobiavzumZy7Syl
cWUjkX+bLKLqtO4w326IIzjHOT4B2HiNe4uMglaMVvXmGgYDkTcIJ1D8yr/nwR2F7o2pIIe6/KtL
txiesWm93YB40N40TVP4ur90m6jNrY3eZpbZjNdBX/nTz8crfIiFltTMMZORPGJk6DkGTM9ROxr2
mgaq+G3PrMvLfF97lce4viZ+5yE+GOiUE/9jJeMX3SS7wSBIYjuOq22sBKAOBWSEaXBXpQh5e3pE
gbQZrJ/srJyqILZZZTC0qwTmZuX7xRoNSrivi/p7O/+1xJpwZIOxEG8OYMY2SXIZqoLnGhnlhidQ
YGaylBuq00S34ovO8leL87p2T5LFgEuGy9mkucPzx26TtYQ29w202O3nFUyLxh2jacul3gRDD2rI
1cWz1P03Jy5F7PZeYWTYyNQ6tUA3zZUvlFso9C7wCynAlSe2ZDrrLe9iAUQzdmXkrZy7MlBl2X+f
6ea84+y7+TQGbHxA8PwIc+0//O3k//fMvvWKyiZvd/DZoCgMMdcd+P3rdBokTyPDD/bgGT2mid44
dPRvUxgAh+U06iCyfH7/VaVVJWQvl75TVNdPYs1HVhOzu13/iDdnHW3lbU4C/jNu36bMlQwNbUpG
kgkFPNp/Yr2iWrmaBAoO0nGfoX/KM1DTZM+bG1yU+Yp2aPfNga+6nn9l3ljOrs7TKgqbQNira27O
xtH9iZVMwegzaVr/N3Sqq3oLmRQhDc5/lbFUUvkf4YD3Vxmiour8nhx4qwhPXhP4OMyEkXpm0RcH
6gd8dU1P3f9UwocQ3U5OwqIh9QMWK8zUg9dKQ6FIBm0BvJVRmG4IsNKup8c2+y3X2IyUdnD3FW1o
iCYFTH/lM4SY6GFGcBEeVcpKJTrBf/1gHkPmsDDsPRt+JrAWyq6fUIlWgaUVF/dyRVWgG1HPG5qP
2aq25llHZ6yoj0vZBXQFW2nGLlVD6tsHwbXTPhr2pDGDdcEsjuoWwoQTIwyHJvDScN2BhmK+O0P4
aWEYKt5BczxKpEcbRmnQOHlvOeFeN1U8J0Wy6FjxZE5+LI+TJopghulYkyvNTEAyJtzFdyQdeRYU
wwY3FWdxFUx0zSiLFkp6sMLWgpRlW+UyQToKWjGjH3JJIZwYp31ENU0U4elCGdODJyaT0FI6h5p/
YKvkEBMBU5aniQUc1Mbmg9YPLFkbVp6F7mfgAfS5YFUcJbaw6VZmEmPvWjDgtRPHiToUddJaz+kb
CKoWr6H1GjHG5L9wAUihFFH4ro2iwb4nl/n11xP0ZOayQljZ9/tcDrVUW98OL/jrcGGNZqAtWlbW
dD4slwvimcP7tE7OBu+6mRvIw5l0jteOD0G3MMjCssPxqGG14rb+J+0nrisbMqKeDmXnwzHhIcpy
IeDvJfxam18oiSbN9ns9JNXtGcJQWCU12JhmiBwna2HA8A+NtkZpYhQQl5Jzep9J/IBWbeDRLTdA
p0EmLz4pcghP3ZnSLVY9QJXiAc1zW1DsSVG88cWNMjzl8hiRRAbpEx42FGMnJn8OhMnVTP7XtfYz
vRIXSBvordcGjsllfNkpKV/V/KCVBs1qrwuTbX5gryUIcKmwZuNWpnjC5HHU6DvJ8KHjc2qebFro
pg71kPPH1ZqEFw563rVQ99B7k281ISHVJCoau3m2efJ98AmntDlRhVeW4N6uVPvEWq8W2XGiF8Kt
iRc14nreRUTZOInfmPzg6PvA7oPEoq/C7kYSQT0/GGtXbM1jKDXwOuIiEYxSwJiE2WokiSbo6yfi
pO/w8IuglbvHNKUrKdFswf/HAYDT0uf46iiKGxLnm5R69zVUS77UygY2sY/K+gxZkdZzGFZsoT0d
bJumVN+OwJDNtpwqtla7IaWO6uyvA3nbt9rfWueQ3ngry3B/taxIE93NgQ/ccWcE8p0hvEw8EM7Q
kMfqnp3zLZ/nfMXEg9NDUqnR0u/vfz7oHBXoPffJ4Edbr/DX7ssx5ayEwBNRALTer7dEymlV9j04
fJiXFrAa8Rv//E7vhF9OOLUFJOPmdxnX93Vt9+OyeXnopOWOYCPnKGl8wxHIe0FtMJ8Ja8ShP6j7
mGxm17+WUgwxZYpF7AWOqR8SqC1ZaWh1MZ1MQm3rb3yGAHEfjgpzuHHQG79kIOQJP57DrnHuJzN6
nWMlKPaAnW1f8GtFkAhV3zE1kXKl44K1ylxHh1mYtKHnDLyj9UcWRvUOlHj6vvHCAObLuVH3WFff
bIVbC39ZgYev73HYxHyMdxOW93wnBGe1/shtF9Ha+8vwQEcjL1JhhvAoGV0woxuyXXoxV0FpZxCA
x0WH9jQmBPiZSV1CsP8yfPXcu1GhB6SuHy7PnSexjMDfdIFY5fDFDXLf5wqnMpp/HSa5FE0U9stE
YBlmUKTWC4Q7SQI0uOQ47IO3G57V1xYHBsYQRj8sFyYtNjqFy+NBSwejXtx/sap5K60xURXcp/0s
Nb2lu7I3xpWCD/RG+OZp0EoWhrebpicO5TlAzB9QSd99XYubD7nbqN3uY9vG9i33+jci2Z+RPClO
96OoJINspiXx8FJtQE/MQXZz/PcNy0gUuG0qPrl4VVxqUkRsxu29YJDmdtDT9EgYd24dC4NkTub6
jEGo8mZ4rCFLvKCWjPuROBr7TEpXPPa2Rtk5gm/sRF0GT5ij6FzaYyUzwBbqRIAh9t6yMRNFybAN
I4AWZtcs9dYJ0K/jF/X+taYyX1qrFygq046+s3muJTrLSjoDm24BMLCNjZeax/Li05wGYOhoMBqJ
Zrh3W+BauCSJL33xbA/A9B4Uc3bZA5kOPb9gaNmEsUUHC8JC60QkHWSUXDo3UiV/WJl/OYwQ5Kwo
n5UJYf+4NLZOvK6z0Wd6cWKtmd1zDD9lx7IRUg4+D0PTbrK0WnoduVQdZ2DM/piDfWvrvk75g0cr
2woAx1PWSM+PbSep4INJ6kw3YXxB54TrVBBUTCb13k+fyX75Xei+3YnIApJjrBDix9/JbOXLWw0u
QLctWM2A8nc0LpBQr9B639QRqaa/5iSXYB/HkeL61LWmkR+8nDlz93xdngBOaG0mNH+l0GDq13T6
oG2aCeBwqsMORr5aJN6Dvj6YK5bjRzikeztGJMwnf2jC/I/Ko2aYmBCKYdgSrmPmy696AWoxRplZ
YZtqMWTOsg4ClhKmFQV9oU6fmk45kJ3v1YErEM9kUzm+h1snXXNNr8APpyDUsjFgz8UXI/S2crJJ
e6+o7gtPnWPTPIqsn4xqBsncs19FUxcrj8IOHkouVrFI99Yt/uQm8NjoM0nVaLr2buvDj1Erjz5r
+HXrn3jdn/5R7A4v7W1uLiEffouCfKlq0ChXMrWeRPtIbBABdy5u42OhlXqkhG2SiAWM8iC9gos0
nuvGjtChrmqw205FlkaN3ybbRI45sTCIlPI6Ocr3Si/nStsxksgYif8oQyKP0ASnbAD6MrgIG6Ja
8XN8EjlkwC0NK8+jikfwTQWEc/u6LxYnx15n6qbFP/CQsNxJY8B84+dgNrH7LpL+NUQomNRYiko/
o24iv9R3/G7jB0JvLuOAa+leRwiQRlDj5TqSnVd2E294+5RE3nBDoGKu62HHZQKaZ7tgOwDMsGrX
RH0M9t018IUskUqOyue4izsagL6HfDp4fwk2Nqrs4O7RnpMimoMl9oWg3X86yscRAX3iODgnD1cP
VjxXudmi+TylDpbdt4jRdixDdwk9zJLmj7aMb3e9/zU1NeSGWueYsdtEc3WKKSLpC/C/5M7HSNMN
YyI2IpHWABdjcgamdsS6dmxFhd3qGot7Bju7hwGQXNCpt0RhuWuv8ivypXnhGrwapl8HgRXU1cnv
C6k+nVnV9Ia5E8TB1gcAoiD5JbuuuSLbQb3cGtTug4cX0hs+ht9OPcAKZKqnMbTJoaN3nn5ClhVo
4AGEs5bcUgH4IlxiAqJR9Qoc5D6yYGSOQlu5MtOu+OM3zC0FsnJ05DUEc4q9lhcRVThZVDDJgvr4
IVvOycl7RQYNN8fbD+/g0b7xUXwi28hUbfCTz6CdTJI/cZAh6dxEZuIDMgQrijhPCRkgDYM/gPZC
ZZBUhWv+CJ9ob4CTxk7Odsn01ZnRKBvO1Y5d7d+opRWXpifvVxUjvpQEYx1zEE6PqCcZgDVaVq5e
4KSlrJVMAEge1wiN2iwBU0PzsKWWW4FEj3zekRhDONWAirXMha5d4na8lrzlNMdYH5bUPLbSiYuT
yEoyRfMsNrXR51GemOZ/0mkPLsgJhMen3o20g+vHQJU27Z0w2fHKXwhyDvLwq8ETwvftXWRAYVKS
mjcLx9ja1p82Dkp/DqyunWq5j2zNs4iFjdhbzUXgsRT4OlQoWXRWEUAdwj8QBKeuz4c0KNDi2DqU
nR8QU5XGbmoFYVOV/QgGLIQ4zXFDGy7+yJw/DoC9mAXOuWZGlFMLZhctyJz0n3NGzOiQhWZmsVr5
Jes573Yztq5iFyjFszGAD4CNXjsK6qf9fPJ7oUz+n1geJ13MT9Aqu/RRBobq9B7t5KwvK5G0RfVa
AXXdPczEK9iEujWueStunz+nDQ+bKAGNJlpOgWlzWZJMTeLsZmmYYqmt+gOB2y5B4U41TKCtop+g
nA/Nz6Cg6zznii9in3kZJD/i8qWltT6ZOitbcERYuvheVZla5oWBhTrw58ZQzTDsjyZZkuAWS62R
XWm6bJAhlnAgAzgPkQHMzA45JGO5d6qNRcOKKE6PERQyJEINoPRTni2mDIXVSMzJz5pRwkTVoh6S
e59Sk9SbVw73hmXQ+EXBzqiY1ktcbQisFGGlLW22NWgAw7NVWnska7PTBWFw3pZOWzGcPmxwWMt1
m77+0LM6S2rxAbBaW+rXIP6ytcz3fJCtZRjh2AKX6lRYQru99bdbYIoxis1+e6kwtvfte5HrOHxL
pwTbVMOWiBCbxUFZ8yxpzbZ9aqRhNhNHh5c0LOnBA8v6XRoI0vl4IJuU9AISdxW+fRwlRoSbWZC1
nHhXn5klEK1GXX9TJPHvElIxjVtZefB0LJajUuqWl08ttccDDGqkMrlSmbOCV7PUl8lBPnrkGdfT
CXLUOebyTRvHejLmnLudgD/ppfvs8mEjP33GWwEt/gbKppJesntBxgSrTXH5yQz8fcPqYfesJmU3
zYgUlC9UQkicK6diziWXgEYb2XvKSmFQwbhg8rjAN+NNonwv1xccAiQ/c47ldCMmOSj+QzQHDzQS
QfXt6HL1yaau+nOraXYtgBJuZHfV5b+IqPsowzGX0N5+Ph64yuQn/RH82Gf2Bh965lgD2YNTjYyS
K63kLGoxxJ+TzxTRuwQkhN/gqM9NVUHx+BMjv/BYQShDBZvaDdHWxi+AUMZ4aL8jCw8HKxm286CC
uP/wn1h6Z+j5+qHlJuu0mAjNbo//xiyBZ5fa/Tn8jk890b/E8q0K5u5WiUmaXZYfdJVjwbuR+2fk
PXb8WSFdlNfKPgJpgZWrVGtJ1mzld34HinFI3DB57bihqR0OrDYKVUe4rJMJaM65Ww7evwZq2aOZ
KPun68jmC/VgxSoQVWlMO5jnl1BXU+4X/UkdMJO7S+HHxFG1pnez7WQZP1MVXQooAyjB+bn53hb9
kI25Sysa7TfSZ7uxFlae1BbfyaNnKo5Agx53ILI5QszS9OKp8EU1XbyYctwcBWMmVtHenBsMiiqz
/PZvtVg7OKHiIrnM5lQFhmGCOF5W0aB5QDHuenXZGtY9UefO2AYGuLpg5FfEJKErMd9DY/xLOlvV
uEoYmpJhJc9+ZEfuErA8V6RdCPXEv3Q4SerdT5/RnYSgNch2i8WUUkWvV1/z6wdUjGC5cGn2OLQ4
kmsY5U+oJRhzOjR0DK8s56wp8TC2hjvT6hIQc2OApmWcP/L51m2lbLp8crN9lbP7rRiy3dh8OuP/
H46zh0qsvv91Lg2pr0ScNBVYKlOed7GOBrGJOyWo/gaLBfJSDZHBFIFQl6ZUmwCnfmKBEuG5dVJK
JNrPhApE59aziCW9KXD5p8/c5kiQkB3f2wHy2EvoXPNrDS8vY9znhn1m4HBSA2WmHodGgaRHrkAi
mVZtEkZuJkokvrjbxgr4HeGII0UJuUgxFrMG9bEBSxfbhNH+tblyFrsGS1XToNHqYcqO1WgwIfp8
l4c5imCSU2jAR+i0MwfPOj4HsXTxz8Ck0lXTsdnUBrg+RxcNUkcUy5+rzAtinADhcJnYyrl7gWFf
tSf41XuKM7/RQyhxtBrU8HCH4tZVUsUCG4KXaA/rK9sTSdhGQr2ENfNL56yJJPpwAo00v6pC4usF
Mm6H1KeFsaV2uZ/V+/+vrdoppSLqWOKVfMw7Kn7nHsTW0MpSVqyDExj7bCQjE20Dn73FRgUJg73C
p3PinxXhnrqmbkrzK0NJEpMJvIsSXadV84U0BY+B6uJkwL1iT3wWH9YEwph7TRyk+8puMZ0rPkUq
AYTjSNrLAh1dNeFxW0QkPRejyLPe1HfhFETdlvIBITxrcXMgR/Kx7gGMw/Wj4poeseqIK9ch6Nhj
8nbjMtKd6YWRKsmJECIb68zybu5FQXPsBVINxYPIyXMWNZ6iGYbTS8h5b7KYHh7uGf2Bou6yNotC
taheMmtvps/aSaq3a+Iq51tnv1VK9MghsXJ4kin3m+cLelk/uRsS1KLbcZsaUF/z+HDqOA88JYnR
mYUI//pE4GbNE9jtceTiQ0NrpQ4g8ZSZ5IvLFuwEzFp8APR8hDuQygIoYMhECs0kKA9h6z088TpL
TP9qdVCm9OjAIuZ8Vk9ZnbSpWLIDazed4ajEHyPLBwYuu95TBXvBoJdHY5Cc0QZm65S8VMJKoSCc
u1FZuRUQlt4W760LOPEAd91s16NKgCwhno/8nM4Zw6GrBtaRCM6qggdjcRrxXF2N/3GD+uqEBD1G
o5l51cIuTkFBKy+EjJn/P34cs1o5iwjU48gHSkg9OopRxpvxVMFRnk0+/tpiwyJuY7a+Z40xVniT
cJjc3WD1ArVzxdpe01oTQkwNcO+JhNHapI/SLXa2Ihof10u+SEMp45l/Dgd3UzNZZBi4BoE2OL6A
NWgNjPx4iDgn53AG7oztl3uY/sZ2horthCmd0sBoFo5SatETcxM9t8lkD3wH9dt+8onYtpPJYxLh
9ntmvR/XwqqYhSld2j3b5xI4W5/AihKnsTrE5VvJTTDoVzbp1BFUlix8BcFumV4ycly7e23F95T5
H5kxgMFVIZlm0rkBfzV2rFDzPIauBye5KLQYNTSPva0B4HVus0/7URNf6zUVX2BbZe+5W3Ylwb3H
X9vUv0cAi/1jrwwxBoOPVPbHxCtU5MqQUIw5tYl1eq3W16noLH+DGAGcoEjCKyK7coQ77BkcVAav
dCrqOeQtvXeOiqMDHaHc0O1/pKLX4ilphtoSp4CaFb1l4i2S43yCuTIP55lauuhelRl/4OZUo6bI
oYwdGQPBW57rJsGix3YZ4RGmlj79lNesRALBUd4cqk6EP4ft+rU71DHQqmHv42cj8g7vGwgke2tk
AxgsDwuSVQ93bdHGuaxNBwJ2c5GkDyckYKf4NjF/EXWbYNa1LCi0bOZfifilUfJLu1MZRvsuhIgs
RVczSaZgOfbf4tlwE2T6PzvdsxzrJrl0wW9XLvagfIcJscQdYsEdeoIHZhsNRCMeUZVmrI5nyJ8l
zNC8oPLGoa+yNFg/5h5DX55esd9zDMi6E8ExJMSon5GBAudm3CUB/N8BfwMzhCv7EJwsQa7bQKeD
sBGQ70VO9sB3PQaKaTD7fIm/femuMQcDCblFv1VXxXNEV/ZNhmBVmtuw4PiI5Asumd2XHLm1xGoy
YV+9SmZT23viKtVX5lv7uHRfbwtMGqxtI2ZLpZjqJwXpwgzxTT6nTPpT3IrnOy55iSi4WcMIyVeS
uiFH+Iv5Hx7F0hsfo2qs7/US/ERraplntcebUtTG/xVYbw4E9kDBEWKEhedj2y3RGGYc7MyuDUvI
kUJV4OGoxKsuoF6Yl/FQem8aRy2rCaNWWWnz7dNHtcFOY0DWre8P9UcE+TUAoY/hFa75loIL+haN
Hk/vv+fC5XgDlM9lqvRDU501yPrtx9WhU0fFJIEElxj+sLZoLTNiJMPxWUZOfIwJpD7qVgovZ8xb
XIvs14bKgXUDapE3iFMcSnHfTG7PoBRr3fNyYT/ff6NlInb/5NTgJequdVqTKlvLMwOs0uStULBo
5dNQvDgnQ+9X1L3ChGqKtv1N089r7R4vjYeEZzl8lHxG+XcWjzgTtWZluUPkHcnT9mxn4nOiKF94
6OT466xBn9N8/85iMT0Brb+TlHnpm5oRdfeG4QJeAoM1H/Peqn7SGpHSPMx7/oCPM3oPvtvUNPmA
Xq7/RJOzr/K8wUs2Y4GF7X/H3GRsKAHcNyRnYcNhsMlrRsB9GEb0rc9Ygs1hSHpfvDloISpNTcRt
+nLGxzu8Mv5DQtJT7cT1Wm578FZsWsztl3BPzFgoyQDSdctEnXHB5f2PPp/NhgjQYAHn8On12hRl
/Hj/C1+Xax3jA/zDIzprWGwPZMB3s/9RDlBQCZBSEP21KPNg9KM+GycZUfh5zL0uQE/xthKUY+we
NLeWNew/OdbHk7H3puLGh6UtU8B5Lgj+/xmKsqo6J1gsYGxIf4QdmksDug5/PyMZ00B3FG5SyI5H
nqk2a0NK4L1nnwIZUPHzw8dYmgO4lLZ57PZVVe0Lu816EzmLmOEn2aTnK3b2OuYii2fMvZsN0Rz4
CQMq9WRgdz+YzCKW77jzciqsfkfzCj8f8B902+QAGK/wCyIb/PUEoyj1K8W0YvzMui6sbIdGhrKs
G1rykERqytKlNJcHRYg7iFlytvYl648+tZhE9YSfarzGeA0QzKwiNrE6OaO9Et7aB7/XmaGrElV+
7+fOOozeK52wCkca4yZ258Z/X7pX6Wpec61QRlIzfGF2i/RzcATLOGkZoz7ZZ8KF+MJGT44OdN26
DJlyjBzkhueduJtx1kjh+XrU6dMdWjcaZTg7IJ/ia6d8CDC7qJELimXAzYmeBi6BTYh05yujMHAC
7mfqUvj2HfvIJDkIz3uku0b5RxSlHRH6PFPtiu5Xz9PjuVEFfjzQbgZ/vswdJmGfHqXjf36QgJqc
lUfp6Wv0QmxbdpvQ/UTdeYgk5KSou0MtLKA2s5p6+eByBYmAUR9EDYr2LsXGzC7bECdMjhjsc07Z
gCamwDREzImTclNbokxvmADRgwwPNrIdmK0Fw3IF9XZMhlGwS+JDkms7PNC2tQf6+BuTRLr9STDB
/Z8mECsuuwm/w93tA2Sqczs82CwwWRW3ldG4t27jTimW0ctU3NH+mqac9t08bDnZoYqg2R4/mS7g
Fr/tduaDy5NmHuph0JKPI7WOCfbs0v7Njn+RfZz5Pa03ucmDajggf7ureLMAJzzZwW4MxO94llDl
QGchGjIFgFFukj+W7f+IsYDfshr3VCl8uy9RrG46PUSWtpTlUb6Oylxl6SwCFhsLOn13NqJAwZ7U
DMirYL6YlxFr191zuq696k1fmYnlK/ovMRMj3E+tdFI2NLdLA3fnrAYpNEU5AeJ7H2rYITCEdRBK
s8P2ZIEGpkrVzTWM2uMl3qmn4cESWjJGTFDgSAIQeL/ewbXckZosUIBMiBTPhm0VptOKG5miAvFH
sM/MfwSFTEmeo8gLzI4W0dgyt+Y1cT/DhAxgsizzEG/or+IB4xevzb4n6ARwK29t5lhT3d4OGgms
/Vz5Yi8PRyz4ruUCCR+j5C41c3rE7wBlJBbZCZR9QNWzC/MZ7o2HH5uRXiar0144AXEgeX62xkJT
pm6DTU7YRcD52sO0/XBfcrPwiX3RopQOQqydNbOL8h78s65XGn5VMcB6AE6ToE73Z/A3pKYf2YbX
/O5NOJKibDANk5pbup0Tk7LBhkf4svPGxfQEgsyYmBARD2Tw2b8x4P0UTXBbv2JpNIzTj+YWoYN8
Bt4+O0ag2vLrVjEOWqGRSjTiu0vbBOUGAK5CIWcp3yMFtNwG2VX2x/MDpabT+8zEpGbvx+Z6Hrgb
fBEyHlSMOrN1KX79ouwu6/DC5uDsDp2Cj9WOSajFPCmLe22/uZQGHB10SSF6+iE8QLB2F8mZHPxd
3evLMRgbSxgWCb1iK+7x7WfmFkHS2xlUICv2Qg5bSUUNxp0oA5DLh7gZNv4qiG+9ew8/d/A+GdwL
F+xg0hjdbQ9h4VebIHd80HOkViGXH/7BX+GNZREOeiIm3UZwkgkqDezhqCPG9q1yauEOC8mUSpth
VNBiFkDbF7mL1GSlzz/i15cGwJmxiNUCLSE6VqPM4OAUceCcLb43i21jzHy19tEvKQqqtQ8k8Ksz
V++/qApV5h4ty1CSkgAq459tdGd9qeaeBsqnJb78TYEn6S/K5uL9lH1RcMd3ohbGGcvwRfq8ADN1
oW4NW9xeQebkF9i/1gmLsfbl3w0rOwj3qhoHZdBN0ndQIoVpPgWVQWB+M0hFkzycaqMIVW2ZtdcW
3Cq6BBJDNTpVYbfmwguku3rHSV/EkW46V9hnJVqaeyoEu8iSQN7er9o9aJU2Yrb8i13vHWvE9jpx
bDpeDsHkPkYtl9MZhWmuc1A/aeX59gERA+sEHFmakphlt/TWNWyh2AqMFYs1pS07HsviQI4W8Lrs
uZIMHcfddCmuXyOhN3lTvLLqJpAYKJcDUIbcl7Ol4X1fVo/lCcQlJ+GynAhliIWVi7RklOK4IPvZ
VFybDeKolAaqv5G1ebdz5gYmrsicMfy0KBcpuFelXiIVucqcdFjzWH+ON1KG36tcLulcnDiREV+b
uSLB+r4i/GvAByZwZl14Ip26tqF7bgFRFqsD2IEGAk//ZkVBtMY/1uRqHlCytrr4qnfpsO+lyLYI
JdgJn9wNCeoq5b3I/JzaZVLwED9AlzMEEUkcbnpDiFe1FOY51XvFpUEFZtSE5RmZ54U7g4LYf03q
c8dHA4RBAv4FHDQbZLJ1jY1MayHhnvUpF8QhgikvFz1DE7X4oFM5wC06oa9+JmBhFED4CIdKAnF9
PMfdbkHoc+NLEygmfwwrafmK5zLGJiSRk+GOWrJvhjTGxEDomxT8Gz2Pr9I6YWxFuwtWdsOvjqVV
fvuogyDcTUlOoMOWSwcvvfK/1/M9yrNUHRL8EWuqeRamiB/T9gFkBrwquLDkY2rKzqU1CobmM9AT
eK9NRkRR7GZ28FBmXKkUpMcnMqFg1z1z7qqt/8W3+I70w2qwtcBzjF5xjpG/LmX0gZi6hAG8qhto
vHb7kKL7/LDIqfnWkLpipYMFsP0qR+MOlXXax9YXSOyGstmTt3EgBzpkly2ulaj0tPF3nOGft3fp
9CVUQ3tg4paa12AcIg42zEUU0QHio3LuwzSiHWGKOsr0TYVIV2pPvvasYZbuMNzwlHnYfIPVb69D
ZJC411HTVLiyqBhV9hV4LmXQ2rpjsDwjhlBS6f8CGVOvtkxp0Dq2AiVBRnIhW+ugW6HXH3lgGoER
qPYLyrO87UiQFmfkn7vkkHzt/wdS6z4p8qzeduGsLbIgZ7OJ+pe4J4++ucHu/0SoAo4Bf+NWhHzC
7MybC+lzJBYrPLgIG2QSWPZ5Abajmi0OzCEynWGPbgWvv6HZjOKwOLgHMKpR5hbTrrUO+xenPLCX
WN5+0W7lu1NM53ThKW3fmhd01fQSq3OSh1cL058Zr9d+qFBxcYeYn46CFQ+xLZwPZhnMqGVRUKx3
Bd75deMCQ8ZzPSmkNwcZtnC3l3ER9tTo0bexmn7nDQ17kCfhV+Ud5p5yiLSmKR/ap0Oc4lPW2clI
b2s28LkpzwhlcC9tSgSOV3ruERT2bqlHX8rtPpw5c4STrn634XIo4zYxOUPPsyP+JFKYpcSgxuLr
esWPOCh6eha6yRaGtvrsdCXg2zHIhdbZsxuHSOzBMTZtD99M7jP9YanyNT0KNxiVNy/hIIlXWKfd
OWlVPgGUg7mO05FCjHrtdlud2oKhXksJjyb+wm3xvY4fClfqYaJjDEPvqCAriMJh9/COa31akOaG
2f2l6i4XODgRi9Sz0yTtffYbKNE5v7Li583MHOEXAu68Ujb4BOjRouNg/9+k8UHs3ChPNRggOc2y
wELW1KYeVPCYcRauMlcf1otlrzZGPXyg5tkCBhDhIe7sqdDhbkLcsnoSijMpgReu3x2mpjXM7SuW
kW3WIodJnWp3XRQucFGimM7doWn/gBtz1yZNt3tn224BfH92fdqgitcABsQlTsOdXz3cSX9sU3Zn
R56AZE7gyMHktwBFFAp8ILxZeb7/AwHFD+ibINoDAo2AvAnTVNuphWg22YwmOPw3yotjOadOk7HB
vtHjkzaQPjrW+7VFVc0yU7dxaesJyX/ATL7lERNrCYoni3No59WpX6AW9eNaUmZ72S3PmaoccxPl
VDngSG5Dy0qAdj0A7LCIyBj2s2SghaUV6Q0AUVFTcYhWyU5x1XTIWykloKmmUOYNJ0NSvvJ78Y+h
KU4iiFj1e0EYdh6+Pv4zlZEC2eSM0CW7Skf24+J9ccHd0ReMCn5Gd1X9PChDqLlshxud16QWsPm3
Z/+Qk3ms5zsqGHs7XINaiirbJHssfVeciXazZYF6hyTWloAMcjUxyraVC5D4GhEEbYpoWaibzKsT
nzmeJg+sGNSpd6/Oz0ic+JfIw4AxcyMQpySvSchZ7H6u/ME98tIbO9h5GwstNWr28fXHK78eeqRM
xHErOeOJnDT4y5r8uZ+ME45/e69y+fgoeg/2ALknbYjrYY6Ed9qWwDEEUYwqo28rK4ueR+RwCNHB
ZP5AWw45UhvjX0fNQf8eMbnv84y8YIiAT/RzMExUrebBHLklmyvoEWTSPrNqJJnJejCrzun/qim0
hz79K2gtEFxJ/xPPX0Yb17SzxVHKmPWXSOq+M6o0IZ0d5cqHnQ1787Htk+uMCBNlfmEXf5c5XRJJ
BEcmzoSleTh2nCBpAizoP21/0yN/HlK4/MC9/2cFG10LdE6iKRn20hqgRb84hRWXq1AEPl0RhobS
GuottsTpsuHgQ9/g8cOUHEOByCOkOJ27E+B2Ttc4X/bKs2EEaikfoVeay15EOYSMvXIwn9qdEPZ+
3qMKBzHLCCk4fg9Q6XTijv0Zzxeu/5WK4jwHOeHDyXOsG0na8GVDkgViINq/sZ6y5uis4pVg7GuW
LjwGiZxsVjZ/oDqFRzGTws0dtl9foE67LXKfBQH6bgkcoeG2EB/GsnRgYBDhK607Xa3TVKvlK9ow
cMw4kjtPRFILL3AltkpMUer6tu9qY2V4MdLAgWdvr0uzqHbYAMFQRyPin8ECt+FmRyuPSi6GW5v1
Hf9syr3QiFObFPkKkoWsvtq0Ijg/4/foV0qFAWt3t4dqsGDOG/ca3JlAWNFfk3FhrCS/XQfN+9He
pFWMG6PcuMkV/92JsRzj+jKGnBhUqrl5seUgAVPE9SO0sv7r8kHrcS8Z1c+6FdZkzsBdS+y5ByO+
VnzkfKMhHz1L6D0FjBUQUWUCZndUsxYa/O3ggXe3whnCsLWmwEjrRaGjlQ71fhFP3LiZTtGm9zz7
b/4IsdfPgitBHdOeo+hPEehG8AyPoDc8/+n4KBa1/FjyNbZrfCPIaSCA5GO0pOp/uTXxoCMJ2yfF
LMUFOjESFoG+nnLwSqheh+SRL4QQ84GqOiEhKQvjey4Y3ZAmMg89dIRNCKLKrjBZ9uL/0P1rwpld
DrE/8KsYrxH605No5r5OKRWBVdAaVeiCt+VFOT3FhLcsyOu1CWKxre5i+1EVp8S+ZAhfXGjYnNki
DuOBxibdlIEsfC6IaB2v5yiulhbPUdrsI6bqr9QYxE9dGNUQv0qTSMyIYJ0NWPSrWOZlnwcAtacN
NcPgPGr6OuOTSl0lkMtKPENucBztMvdOZq92pCV90oAT/Qq63MwwI8iLBc96E0aTJoT0JcwPVPBG
gBwPYJtYu1AFuNsAz+AM3WrBM+U904HqyXL4Lwl46p2GFiAVGrlKQIHoGqOBUFzu7taL+seueqQF
5r0Myr8b2BRE40b33bvYySLaEuFsBIlT7clcSCneC7k/68iM8a34U9Iwq2Iauue1I3u691wdlb1e
BF4H6jtUM3icdrNg5+62ZfxxSNgKH0+mPjtYwdZhi/ZQC3nPO6jm3YtxH19GhUP9YvoNucVhtrie
v+CUM/wjgS461/9hi4pdyCFEhX/HkbaeRXXJM6+ArtDXZQX2ZopUkikLfxdo4ns4DR58jjrks2Lj
6SS1K8KibuggpVzh3dU3Wy6bZ0M/7jLhrlW4YwAVyxBai1gFZLmneIEkdJDGA/2Aj5ElwD6Nx+vc
3KcpVP+KvGo892j9508+TF/gnQSQ3OWGt/DDAUpzK4ihh2P5w6gCrMrHjbT7hDvJbYjEda89EbuP
2tS85KFtQcS+GEgoYtG5DgtH40yZ6B/ColJdIxpt2MXGgvimGWrIXRTTGTA4VCVei49ZRQ4W3F7+
R+Tf46r8v6tEQcDhhvEfClIe5M/YKe/HlJNZAEOjetExNVAxOCxfIvQu2ai431rN5ebNPGGBsY3Z
/I4TZ8qkkzDRe1rhx6Oe7h7n0QUbrrBVoTDxxvJxwQFtzvNn7fOF5NBAVoXWbO6WKR4P0Hh70jUH
VcmQOK15VO/MDMRsDmo64MltvCto8fsw8kDoa1UjRE4NcDewkGZ8LfbBANQTuSAqHOnqLu3QeyVI
ioInMojkjXah3ut+3pLK6FtsLnFsLuGD4+y2O3dUJQq9CZdfAgiZSVo7T50jGahCsxfqPIYT+jli
Xi06ow04BPaUOjlZGYbNnMWzkLwtejwzM6QdG3REIuBRH5vdpuK5MnK7HxOdfntqU6Mbfaz9j4fG
bEC+03XdZjUM6q6gDT+1FtYsLUWxI4xVKBrnlJhUVoa0lTaFCPnEq0QNoBJy0v1k3FEm3HbfNk/g
FYN/B/QrcpoT65KngAj+FC28gnraRbHO1HGOKY8xlpry3zAixwoT+fi7T61W3lCkdSOiIe+zqGvu
J5i470gOSE0JNaRCVPnV0GmBN1pPdtN6MOOG1xdTHLnIP5RmR01QnxcWWRCu7h+gb4ATEA37da3X
/cXcY9yIQtN0QkDKKfdDcgI2Jj811UtZMa1qU0g1yJszetnyY0eGmM0qdH0RhQySDxjgbMHxMJso
1QurpOiv6ugUe1HJNsvZkWvDvSDh4GefHfpIoc65jgE0an/xAvBHF6QXqPIeMMX75ImdB54aXsyO
/aqVnXsn26YOBoOA0BkZtFAMigfxwigs7OwnhKsDEWAPNI4wDFpGlTsmQXwlnet1xwdHbcBl8ZA5
AjmREjjNfdLI/dFqCr1SRmec+anbtkKyXuRbyAHIQMRMdS5s8qPkjSZh1oLsoEB4QD8QfyHuujjx
C7pCahsMoOiw/S6axBUn7T/X/GE3P0LSQOyXSOGSvA6JjhC3nW974cHvegZic5pF5OLqRReek+ix
8o+FKRPH8fOqB9s2rBkxhHVnwkkH7Q2e5qDJw8+Z7sNQ9rx5QvoNJD1LgYC7jRSs5PA7u3YkEi+F
76cATzxbfyS6ddV9vnfy8M40dnk64CWh9gcflbVRcpw+s4TQtNJP2umJZ37gCBXBZ53hB6EhIm/U
J51ImoIkBn1SUJD0XPzB9MaMX66H/Tg89+zh+NKP/KPzS7rE78nQ4b8K1gpC8mzlCdxtXwAcQ23F
vthpfzCNmVBxL9CpjretzjscqEYrPQjzFX9KYAcXqu40a4IuLC9+bnblCTAJ+nLKbjq1R3mwxQj7
THGZGcAZv+qLE3wjM/MrZr2H3l0G2GwTztpj+7Nng1QJuL/dzKS8P/6BTJQGDmD8IjYuDfY8XKYj
BZMmFR84eUWMSFRYZT0X48S3uEFg8eXGAdAawLWE/Xe5F9njhLg1N4APQXEzISmTCKD5ezPY+Ok5
sDqrEmFR83UD3eGaGQcdCi09ahbr2X8Fm7l4/FBzdWlktmwtwCFIMqW8O98hhde7kX5eN8QYFIwr
U5MaJMDXuYteipVez3xTgWQ6biEnFgYHAuhKNG4P2ZV5zguU+MuJnjTinFsoWY7zWC/hJXcKeyYd
u1eDWdr/Kjcb4WTY5NIxEF7rJJWZTuMHGEvxKRTy9En9VzPX8rNgMJZZp37K7bEbd7gtZyAZVIbS
VoQwr16+SbMLA1xt2rTbXnnC/bB5DFy5S35EdeEPDkqmvWun59SOyfNlUIgR2ioI0xuF8zSkK+5h
AAybLnJ/5V7OfdcpRpcyI/6sNVqkEfexBqPzTVL1uf5d3llMQsi/F2uHGDwMD5fdEWYfFRtBvj9V
gZfen7bmkmEoN8ykmZC/PkpsszZkvB9RzrpVbWpnXXVkF1atPrtSI9vQTFFg4abV7mstT+HHmVd4
BJPa8r/VR8EZO9bJCiyQYdkZqrrFtK1dvL9/0JnT1wnTIW2KTuJ9rHpg+52PzarAvh3GFsp09/f3
CkrR7YcmXlxJ0EfBfLPG0Utdzba5QVKn1I95xkeITIHsWzO/vwZLs2uh1ULUAp93FVmO1dGhylgG
kRTE0+zS6k0u9Ezyxc79FR4axNs9rxD/qQqKgRythjuGB/qAZ47H8OJy2JIXLBcQEfCW0X4sTF+C
oatpvxECxBSmrWuEHePFfxSIO25dLv55KfrebPD7oMA2orXbvh/XSJVVYzBrlS4xrZu2qZUMCCrM
HZgO1Jo42toks4fuvQ/zEDTY3D6n3jQzoevunV83Wn2GXwVLgB7GNRFDeBfGUP3gIrEc8TuyUMAU
xo19UurL4buP71ZuIP7RRybdyQJNq+OqAeUQCiijG3APCgx6LxpzhPb2DbwyjUD6+bLycOfofoYu
1D7B4CrE0F39YoJBKFNsIyROsQhC7crQ2bwCU8a+WL9o1cn3lBeShXoaRZ4UiybAk/acPP+5PCqf
n6J3I2ans94+6xdBKCx+t/9RAPvC0hysQmwG99QdTmfaL4o9/phmsGPFJED0JG8kaFO1zaxbw5ZO
XnyIW3DxipnZgVDdyHhKqSa1w0cMvBMfaD27ZN+XrXv6dmw6+AYuKhADYBfepbPv7aO8CFYO+OeF
1WYTfk4c8gx7PomTBH4ZHXIik5mbIZj55uaZ/3FK//4oca0oq8R59Wf6SJHuXY68Bkh0jWUIOoAV
DjRUJOXBaE0fAKoYcYTwXFqwK2HKb9I4ni28eq4JcyI9Lor/ZvHzpVIR/wz1KG8fB4JrS8Z6X/ro
yFBYOYGfTvaNC35gw+qZ3MWbyzmRSeahGSF3vmOL5zqTT+YpO7T8Xf7tyHmfJV9yQvOQd3EGY3px
jwAdGYwg6t0P8AfC81TjwP+UvgTHrUX2LKq1IxgRfAPCkUgaSB6y1Nr91Vt0cQp6DHIdJ5tl7p98
NX3M3ilEjx67943S2IR6pRAIy/0lMWQAWCtzIWSnoYIWJCI2PbcxL4dREg8HlQqKeaWtGsi/1Zzt
GeQSqs9NfTHezxHDveHC+PUGarqGY/bKJiTUvjtUlLKqXbPHCPrj7RrJJI9SonGd1lAYWqg/m31R
3ObmTFVZg0MRBZ5MFoj1LXieCEayds9sI0uONsWVFS5fcFzix6YSq3bBj/nQU1eQtlxvVn5sVmo4
8lqpKIhTx16PSaPF6OKGiGT96yt9mBFJOaBPhUo24NorUnLujksYtX2rLe54dcSg8Z3QMtD08udT
9FBhXXSdPdNbEpbET48KUbUNCbjg8sn6bxazkzrVxCalGNf1OR6Nl12qD55LxZ/wQ9CA61qnwW7h
dtHhDzlTNm/oXvLjsKtaIoMqwQelzW1ormCkSo88jSSeOTpMPoA0gnrz08U1nTiD86h0+s5rNH5P
9B27pHsHb/gLunSMLVxAHDrmEk7b6oCKu8PPaZJqQJuwpGJ4iN16QtcQ+EqD4CVvco3ag0duuSvO
esHE4assJQ2PGrL82n7S5bW1CXX7CvzRtG5H58Bj6cy9AISYQfh/U4wpjf2Vaxju1ekSZH2IPxNd
3lTfcvJ7iq/P1UXpkI+V7pDl59bRiKCrh4PFafBrRu/zenBVOSlXmfzwuboe5Cl++xoZGl6pEYoN
piZWfhmyYWHUiB6kMSeQMyK0WanLXzM3JK8bpsQCyqzZ+aMYUOiFj621Ac0Y0GzOTBmZO7BOj5i/
5AuLiXq/fdX4uFm+znta86JY2jf1TZVgUwpmmfPh4U3t1aIETzDpFIHjFC+Gr20yenVhW2OtAdXe
DxLp85gLC4MzDUDnYgrwxByumbcGGlpgYk/RQ5YGNap8OKRfZRjr9B8B9929iW7i3/GXEokONPlL
RWA4x7DrERZh4yy2zOEn59j+YBDdNvltYx4ueDQ64Ld5eC9gP0y9RQj/7hywSmVW+x+ByjHcT1oQ
0T5ZmnZt34xSR8pJfHybG7alMlYnAJh5oH07PdBBX3GeR8nZybJcvEIP39ARtX9HVMzY9KmhkB3S
dhHpq7nJ3VAJsv6tKVtPYSpNrznrSwvySSl3m85qmlpGvs3Bm46r0oNX8RWOEqSVCqKcBpMbpn8W
FZ9XNIwt9FwpXmVsu5c3tTU6FgSkBvuJqY5E16fRplwLMBRLEeFGpCqPMoJNrwPW/gmbyqmWodgk
vjoMt7kAWm9QUolelFkRYR+ggt9WEDCEiH76HEfeasphFHZSaWMZo1FRvgMH694pw1dBgz4Fy+26
UoaC6QVAmcOI/AuRm3siWVn8FITRi0ka3BUyX5Hu7LEoNd7CggV7lonh8GKE82JhzHGbiR+GATKP
s882f/MWR7CJJ2o+QF1L96k7DmvTgn5gpLty4cL+auZ4kjdQV7eI2llah3nvXXibXUg0vfKkJY2B
kEJ/V5iIROyJgPk9txZNjj07xcAs0u9cKlt5aBIIRxZ8j3r5YFant1h6TUZMZ58IJkTr7hGonyWU
gb77mRPpBysqiC0np1uiAcqO7oYazBjQ7ut6rlAqfV5k258mY70YOjvwFms8zgZX/aqCIt2nzXuC
bSDyCyIg4hWQabhXz/7oHWyDrQBwl+qtDQ6nqWRc5SJCyJMmwpVj0rk4cLp2e9XgyEEQMRnU0Kfd
wXoVoX5MstECiSZlQX/EshexFfoDVGwSyIkZv2tkQPCJvJrXOeCcpo0zDTu72UpFc/0SjUwJbX+0
uyCoFe97x2cK/dev6vkJXtxebxSUpCiMXa99ED7rqy/8weDf/gcO5GryG/PeYV9oovyTG3CRG1HY
1W6aElpMUzZSL+SjiDo/J7NQWdo35TQMd67Ac9iT8olJksLEbnmpT9H4Jm54ll6grCa+/nmvl3YT
S5sGLaYzJ/oGRZeKKtBa1svNX/whpCUsiGsnPMXtEXa3hXjMsiu00V2YWWRE8Gum4vBuvAyD29oA
jnoqEMUnGDC5taRjN9FEOYhdPrDPGLxIdeC/Bs1YYdJ29+aYS8RNalwaqmxNogJgPjOJ3XbuA8hK
zs+iMIT3VWj9y5s9zK5shdQtnu/glwoXwTmfMQcu8y/DbRu8acYcaZY/1e7kctRg1skYMMdFqJPw
zQhyC7oLTvdqQm5nXCEaQSHn+R0oMdu2bbAkuTUg7J4NEdoNSWavJfA3MT8XK3gYUuVAF0/b7bXv
TT13B4MeRsohI6qqZ+R1qfd++TEgvMCxP8PIvOnBr+l8z09Viky0hIhryW5KDUuHRXRRtSD8Dj5A
f7mdFpjLN5ndYSyK6Ul9OTjXrxpSMsIRek/4OkFWeCC5Hsmt0exZ622eHGLzybnz+Hds9owc50sF
boXZKhQ1+AF8iGYe+0zQztF9nllVO8+IUfMi+/w644TjWuI5A4lvUDMIaonRWoy5lYhEVdzjvPre
jgpgGdDovbmtVjJQiFsfL/JLT17Zjm/mgxKs1R9S1n/jD4IHb0VEGbH/jTkWGtGdgFruzduEEhuo
4V6AswO/+QsbR+h+Uw+ohLdpIAAlPDSBFmbYAPy5fdQwK+2o/rqzRhCETJUApt3Uk0iorC+ZeECC
ZApCjBbHsS16+ah/h/kG8cignuT+3uu6X4XeKsLol2VpY02wA5xTV2EirX1Z/Rn6ZJLjqp2kObvY
Rmv2JnmEjxF0KqUJ5kFLgj1uzHT4DOr/jstGF4OWg4kuCaupfoGN5BtcxYx8cXRKiobxbq8LzhGZ
R+Ik2/CbeESlriDJP0cgDi5lz4LHSEiRgWIdzhkBCBtnTgHP8nRDgrhsHcHG7iKPTvsSke4GD86W
0ZFLI6mkl1z+bd4OdTHz83Tgr7cOhX0hAqlRcxDFFdAxkrmoY3L8bPkSYH0ua8eZiMvublITWbzA
y0l9RKWnFsIgL1+k3rPAQNOgwV+IJHgQizqkY5eantgEpTj9byW0uqiuZwRAe4BM7FacK4S05m+O
UMreF8SHLI9aL7MHETmtme0Z92aKzU0GbRldcF9fwPxUMY8vlcBwEuanaRHKztsw+hn92tAxj9SQ
WMnV7N/NhyFHKIm+KSYigYI85Y2j8E20vfM47tJfKobFKUhU8OgEQDZNhDcBGU2mFBhMyQn5TzIp
9yTAOxy132bK3vahLeTGe3elrHgmYYyVE57LBUd0pAJQPA4E/6ZNaEjojwU6ezJZGHosr5q2dhJw
9CrCy70kMARzThz59ikFr9hX9Xvdl+4ci0wNr32dtmwhTV3/RF50n3hoLTSKw2KENTx0PtJTyczr
OQ6ST8XPJLncVsNOW1nsU0ZTBinQJuQFgXvEDGdyV61He/obLUyFAHKvIlhxIie3J9wh3aZ/3+TI
MPWRd6AXIGUJWj5JTi4Ihe/qiCQio2dY4Zh2mzv7Nmd73wts+RVFPyLp8ozOjaKTXEB6kbI7s2p5
xHFM2bAL2EQoCYqWt2vLBviXYN6y1JZph3vz7Ox3sFRTBu0uquUf7/EKa8wDM4zfpFrLdPb6kMir
u3DD7tjmnyg/dCxid40A9dHQidH4hynl9KawotHfTvr5zm8dQ7lUTCYhA/C6S/HOv0JzbSGuEyCF
16wVNbu4T26iEI+W+h1mHFL/ooaIjqXC30ijHIDwUY1Mt5ltjjXtQJusgc37fi3aVgWq2K/JB+GU
5CXJsBAo+zaMko127Zxs5/QLmU8q8xERVV1GTohtpyXTtII6ZUipYnNhjOVcJ5XmCXyg7lW/R9un
n3pWq/D4e3AxlzOxC09M4XITiY4VudhFeK8CUFf/gCZ12Ah4pe66p1ySxLSk/8eA+pp6lVI9C4qm
8OgVk4I2jYBktikPDrQU06V8GXOFxGzJWTJG1Y3tv9VvjF/c2z1j9jVPW91Z4VG0MST/nnQVlf+Q
5I9qapzJA35Kgkv07LIY9VgVuQEFjisxoZ09HneHOnUJcx4bH+4FDy9XSi52CdfqNMu9q5KnKnQG
YqenAe37yE50uPBFEyHra3J1QDMYWITi67Q6K5kHeos4IrsAbqpTanv9nKgyF/9hgLRhyZUs+91I
yD9maiGAaAO5Fpg3x+F2w64AaHUS23hiq9QF+gsoyE5yfivdnW6fLVdd+4r6InXzbIOUInHEEoVi
YcxTgCDtNf99cBIz8xKOiLgMe8XidDK2uzCVDF9NPKtW6Q21sXAMiRbh42M4o0djvP7V+TMvasMC
hf1LcsC0JuJdzsEUVVk6VnTAxWtnxCCQsZsonCmTBGOEfFIXZoaXGBZ99OU33r/6zESzd+33sw6D
sr+IQm9BXOFNKKJZ1kpUDNBmdJwHH7LL8gh2XZueWg3h43gCzbRJzMHx2MTkc+o4VhzwODo0CrkI
9W2gecK7rEftrgQQBDw+7sLg8QHSWBgVIKTozPwO8V0USc+h/jpf4FjM59Nvd5hONWM9vYQLHOj5
pJMtjgRu7kORfPJwDewSwVQkZxumzerrPvqGYm/ZABcfL6svnM26f6B8hTlmVS81hLDV1Wk/zLZf
I9xF304U76J04UiO3RLZac50vH5MlFk4PNHQByHOmrxy5Qwzdm6NB/iuAyHAxX7rMD9ZMVH62jGi
6LW3LXBrlBlLAYGaMEdFW8ik3HhWe5M0S0AkwSqxUtS89ITsojXa2xLVLvHX5nAfIjr5MGCHEiEh
Y4+Cpu9dVbTOpIe4bOIh3qfL61tS9cx+/bQgLKRuHk1ZY94dpAkuS9by0RZW7jkuX8hXJSqQ5/Su
CtRDuGLv6+MiPpIXUWsNMA7zNnrZomeHBrc3Ynj7WTlQX/Z9KTibiMbMlWfEDB/Vy4CswyUrV76Q
U0T5tRCyzlBVjHR4y3OlOpTq0gAkrHR45ow1M4N3PuT1ZeEPrIaCefPSVQgOaavuiJh9d23t5dLp
VheNAL3MeSiVuIxarR4huDk2Kcv3Hhtd1eRhTYAXiL6dKsMpnPZL/2CPjYSHFjSb9FSBUexi43TE
h1Nl1j9EAEPm5BSY/PvXiED5rF757g1psEFd8Y5aBnpMPV/5MYPHPVyUlbXEhk4fIl5pimRJGPbB
t1NKKOZfKpFYL6+Zl/JSZo++ewH/gRU6lRcp9ta603R9I3vJua5bw8BXoM1s+DauSXi5mOStbyPP
TQuVviTI2OtBvmNSesQORBB63YYI21JrcKE3u/zDl+go9bE5cXkRndxpcxsNkcKAxLGftvgCb8LZ
AmzMSydqJbN6Jsmk6Aqqd22ANd7HO/nLkAb6xMLPyuOUykSYAwEXHVeJQd+fZRRrZbABDYyBmqhY
zfJg6aztcJKbY2eH145gcAcTY2Atixc0KzYJbx45YlHytgvBwedID6rcvTC8opeQWGm/u62v6ET0
nuttaCcQ3pg0uRUVNufZQw68+582aFmvwSP3g8oFdcEtuGfiWKmacAvF3Nb8XdDsBZcqIWwY7iDY
3daIssVb9M25Po2k8hkTPJ24rW4dnsdbCbwmllptm5tG2VsYupFlvOhITxZGJX7cIH2zrlkQozpl
3bdrdOtXHybDOxA80soxlW/IW8X9dOXgSCKqUkRYsNrF5dNWAjpxc3K+T+Syk3OtXpqiUn2q341c
v1tu/y+BlD36dl2Szrx/yKpdh3+R7+P4+vZRHoxR5cujKyleWKP/A+UNOaQZ4QMeHgD9HolkRaoX
eb3/FAnwW1dZQXz0QaJOHp8bLcx5qE0rJ5z6OTsA71gNOjq9vcZ5yx9XBRUB3syBUTbJQnrMGyik
8vi6m7Tr9qPybejsf+wEMvrQoSfyD7whO86BeO7weft6YUOLSQucRd3QS4vgEgnrh0lWYF0FHSAH
jx/B2soAqVuHRhbTZtxa1nyoFOHdHURQl0ZX7Qti4skLBnQefQaaA9V0xQ9M7ib7gAInn4c5yhxX
WHO9+6H9BqCKvJEyjBxOxN2Sfx4sSI7wt7z64MkNdacdnVYhM0COFyoPLLHnneFQmLwSHIZ+eDSG
CYx6BJoTuRjuVa8K8NcNfcL50MVCcX80aZJ8Btk0nmihm8U5UKXtjRXlKbcPjqHTaw4GZeNvjy+I
XrSh7vhVo1bhyVeU7wkydZyP8oh1/uxv8OOJ5uVhWTy9N9zWFRB+C6rsUhg2jgRFBcZ5OulkV1V4
HAReh3nFt8vxqtt+0k+1iwSTCNiRNOv5BKvBXLffDpen/ojnMAkkKwL43x038cj604amzU9SYiqW
qTkdxUgYSm/YU901AeHTd19Z8hQhZkSd/bTMJaS7TQzQh2m+gXPdfJXnL+QqvWrNGZWd4+zRPEiq
lyPzn8aqjOGLYv16CRh8OB8zW1g8fkvkvVmhsPlhND3UWf800A8UQ6VEfeOd94c1veLMdpsfcI7I
mxtbBMfSRoKNHrHBsDYqfPjnaPptPu9WZD81tlqpwtXkt1FeVTtc4IyWbF8lUWVLVXJFV8FmRwZF
tGF+1dCG3K1SN6aXSOyeeOSmbEaUO80q+W/NrcPFzi7FMKjx8lSgKNUTmt/pjPQK5txNxSaEysl/
p1SPRmvg8ULTwcdHDToKx+bwcLr7D7tBtIg8LTAtLuRdfdsXtClFJLsoOWL9+RuTtU8BKOdGWjwM
/0bxr+8EIb4Zf2MXICVfbFQAm7PmXbCH78KP/pwOGqvtWvUyGYLeHbwHPMS5iY+9viAjeCkg8YRG
Rhm3l/0Gpk3dtPW+TpIZdfZ1kEG3uPti27qRtldjSkD2ow3qqf+MIXQ73pTTAmhE8gTnpzGKGvFm
JacFcO17amBf3Nqp7b4uZjuIEIgV1OOb72LBoDjvWwdDPCOZbI4Cm/fbeWd4i80XlsTTYjmt45Wn
nNO9K3/Geru+xWOw2vETkuYDxmOkYRNL5+AaZUTnTSw96b0SWq1hKY4FS5tZPPo9sAahjB7kKr0c
qbD718sTZnOlC31EV/qdM4XLlbgetk6chU1aUHgvmNhraFfXVQv4jedkiD3lyJ7LvVXnlfgjv2KB
Z266vxRW1OBZ6nalkswSLyNbllbDPHlrlh+R0ABOeXsTp5VY07wcQdcwk1+7x2faqM9gaf7QxTQo
KeVmTqBChFoz2x6JrCGghRq/2L8uZm90PhAp/FO26hDBNii41Y8HiLpXoiSUdnxRue6SjF7vl/pC
HB1y+k7vOTcqenFx7I6NeGSnDacam3SQRBLyEnRWmTENHcuF/VpTxWM0aiEJbEm938/hNqJbEGys
E9k9vYtYj67rJX4zfwHFjmiyZyt9Fpz1SH89wP8VP1RmxtDdXkJ7FipOZ8PuPd416NjXuc9C1RTD
gQ1DtKGkaV2abHkAMyfprSw432gpIDpVyieGuGknKyC1t9RCzQPSOJQQEdv60IzYiax/Xg7o0WxQ
UJ8OyDN99yhqZkRC7OP+F5H5Bh//lkGfTV4OGXXjNBKIWLmtRYDa7hKtcSZV3tNc8d/7mHGcV68B
DuYiBDxc2TjxmFbL1ktIJtWDi8Kdsq0pPbng5H3PvlVzM/ukRdd/ket5KKtfVjm3exW/UEJVIGVo
qaOxKxK9Z+9sBddAJ2PNcWgFPnRnRaKwwMo+e6MPR9ZYJPLQtZ0RkJ3AuUIIOUq0jsDrzkwRk4Jc
k7W46xRs3k1radMGSRpvj0T2PLb4pw41UFtpLYcnwoRSC/FmOkx89eL3FkMdpfV+eIu72hSaq0Bs
5L4nybnGYcqVgixWvzcSrCDWh4pkOkD59qrwbd0A2Lu0HMsKIgHRZgCDv6NfI0nP2+R7XZmauckk
LMYeqgIHiyWSBIKIzTeGYfAQj3ktfUMc3P9guqpn4fsD8zQND7J8qxjZ+kDZBH/28GT7QYw5Sstl
+Zgd8iamh3TYGVTyCLc8vyBqlckCHOrC3Q2DTrTaehrF6RcXfZaXUaVBviJgK3CtYZqWmtT5LuqD
1wfpEGDy4fF6KRgFe3EsSkXvf20r6QdZ0018LPT18J6jKYBnM/FvNTqkbqDO+LDuLN7tYn1pYUq1
cUZIpO4HeOTZZYdjaADrcp6HpBFIEySKx+v8qbILQHksQG0mQb1oghRgJcagzYBL+d0EGX4tBX/O
b1coKfLYkvuv4po10cXlqVoL+pGEQsB9lGs95OGpbaEVDMO++gQFm35gytBojMcPX+hnzRV8MWaj
mO4S9sxAW9x7xmellXx42DnUL2dkO9KPIN3qCTHoRMCJnATMETDYq/g08pHjcOERFUnhdvhKmLqz
1vTw+e5IZJ+OPYzUELTB4wUIbYj111+rY12uT83UTq9Lq7PHDrR8rxRMepc/uqPRmLF7DSE0ZlUY
mhJnhNb1Br9kgbDboDSy6UQRTlZ9itvRdbzZLdNfwsnHSFR9QdJvp9thJD4a6UIlVcstaSgLqqNQ
SPlWoKs5iFQdlsQOOcnbhqsQh+tLEgtDgCM9e7q6oZaPVnWxKI0kEBiBInzz+MeT1LcffEdSN7a3
qgnN7mfe3U93B1y+RJTCda9Tj/WRG1XzQYmvALbMhadjp4lNc/qx9LIO62+0eqf9O22QXd89OIDI
Z76Hu0ahEkuD/LmBfwJxOKZ6CthTHIqKDB+yCLk1q+dIvuXJ2gLwMGOhWSLEKgSEBXMIsCYtBZvU
utEaJU+4hq60r8V/3ymwAGwS8J/nsnZqlPYXCY3nF6XntW21JeXcOiR7y358S7qk+VISKclff684
ZfiwBrBlIyvk1FDNcXQy15gw6CRaaYK6M2Oy0LIWnZ9Qx+/8i/4CxRbSncyk7cQAikxAHUuLK5EK
Z/SC5Ap2Q24fH7bXgNGeWeMF/TdvLf5eeJwGc1TVI6Y4avnJT3SNVHz920S9wDl5ZSNO6o3tr+cN
FUxnTdHxCopfkagoa1qRlyPOqNThBt/cv50Nxfc6m7nNK51tALTS9WAykP+tQ7PLoOu+Wecok/Pn
c4I5/BB9jISIJv95dn4zA/54zRGNro7qVxVYzcHdFDQAwyNEJNFTZxoHip9Km6iZti8Pxxgnn2fY
p4nfccbZxbfThbF2/vsxJ43vj3VdT3wxTr9Nk/7LiCOnJv6WgBBXNZzz0yCnTQDm4Y34UVc5uc4H
okpO5TkVYg0L3RG2ZzH6JhUW/8NxvVe94PgHCOpncrDITZyAyQOySEDC4yqfBDGVCG91m+MuWXpu
/3n5VBkqkQaFkV7F3lwgR/QGs3iKCVmiyf4aZpsW5edJWCc0zqSrtcl4iyuo1puLr0SafIxLtK91
dh2HsQKpzHUEdwHOLfqnMaHeQ4lnxgjwazwBZx11BrId6CKuIpAN4fU98s1lRF+JpX0M4BEwx3kv
tyWCuTxXn/5DDI0Fem+b/OUFfYkqUMVsf67IuMRoQ7Jy3LlPS9dofRR3XIkFp0JSoB1oxZSsLCLg
qzr+yxYCmZtaaW4SiC+dEVggnoqEQ7cUxZZuu2hz0Xuibo0bWrCbgDObjJowJcTaxBdMkO6pteFG
4yoJbveAyrf4JkctE9k7HIlV+F8lKs8tnkGkFrrbm24IOTfczQoOs8jnuQxetvowh1Rq94LSeIKd
0z5vnWgvQsfRLydfb9v4Dhp17pAcslu/NraxevE9+zqWJY0V8998Pvu/TSZ1mxsGJSYQFwyaCvuY
a7RsAIi8WYQ/Oo1Am/dqsF2fZrnYWQdOHMbTc94xjXhUWQaJTh0+otsxTEl05HQIQfto+osRdz6S
84G90EXQgm73dhI7DGsteL0MJbDenSF7DX/r9DG8VVnOxObKiozYwel/WXtwQqFD6tfYxaewkhQT
KZi8/39o9FH3CeVCBar8lLZ2eeg0FY/Bz/NPSZ3hqJavuxMYDB1Ez90RphPvMqfqqCx9Y96kGtOX
OYp2eZPOlfP0A/oGROGvSjLAUW3lzA4VblMOMUFA2bBxacDR74NyGN/eXEcwYw0eapJwYegoI/tv
VnjJGGzFcSkHvkTD50xaOG/oZF3Tl2CFsBR8NCYqV/xes/rpeb5FxOZAGyOfIFcmzaIYqpWbEBVB
3je7m5hc99GHao1IqvmNbHDqACnXp/NambRHWzME+K6Kz1LCPN2HMWOEQEiQXV/tBf074qlBvSFm
BJ4KMgpww+yYNU/AdteGL3JfuHnZFhxmmYnurjo9tgwkkfmV1eHED9kVVxq51QqrLIL/V/q8TGu5
0UmDM1qy6oattu3h1iBXmCLN6ZSgPwTHZRt9jEQM182RKXgozKIpQWebe2jRobpgMQgZsrLagNkZ
HaAoanp2eLnXhyur40Y21M0Ria8VmBpwxi6BzItD0NPfJAoJzFyX/GgS2gc1/ZHe2o1UZoPz1Hpn
acaLdmnbjsX/EKtjp0yw6r/Lo4i+io9vr1j6fy4IfIoWymg4/F0bLRnDH4T2KjQcAmmOgJhNCS1W
OrqfJeKftqXM2Ro5rnLOafZ/QItBJNaHsVUiSyfUkrVjkZh1esYr0EJdqyJ1b3noEt1h3zJ6frVY
347Nx8zXsANAQtivDxTneM971VcKk9pk6YxQBEkNfoqzI5KsmSud1uo8unUgc+MpZq0e5GMOS++w
aXCGdlHgqF6BVUo7sDQpitfjz7aoDOSKCnkCRh8s0c3vHQEonmQDMfUpDi+6sK2+L1MQCOZWr0/H
KR9yFTuW81OTVBjfRPW3joceOB/UD6nyTNXUfXz81DfK74EQ/WXmeiCzh5tyRy9LTPiYtMMKGG/g
SQlBLaD5295ytrd983BhvXT0CmIA49nwLS1AD1Veh6EPe95QP0Y0OwwybqsWQgBqRZA0lJx+N9VI
lXBnbiEqROKdP6J2M++nl+3Y46j1hH0B+yb86Fz6TFXoEyLU7KhlunpafJGgypVowefaHRy8J+Vh
PglaYtj6x5BfR9XQ5nMhqcfehFxeyqvdWYvINJP/lZeAqQgLBEq4TN/6/5eF6Y7+LfZ1KdtXdU3Z
Vt1X+YiRDNhevoDV059gKiDK0xWRyKJtkCj7t0vjsCQfCd61XT3n+IQ79AkkiFy6he3KcJeP1+Tz
VR5/9JO49uIxmDzP0aARBXLl71cqkhYb5Pe+uYS1TdRbWjk6sNOII3tbdvpKZLyRPo5IuvOPUdpV
AD1Icdzurm5hCWcyadVwfFU82aEcurYdPB9V2VS1HKHbwsyBy1vOBwUWUCy6XorYVoobEAhq+15O
OBTIiFkrgQeZbADBPmQ/USF7XKDGschIJo5dnzPkVgHxF57WeKrD2+dFLmntq67lZ6J9GuE1jjqJ
t13HgOBBsVBUHAluh62Jg8nMxtHN6iywnLqN7rnpQ6Jspsk6IQ32VHPo/nfGMY37zeOgseRPEixX
zHnFShnRZxR7n1FI8zTR4sb0HFgt4Yn3h10cZCda2kEpsB8kp+FZUYFtCUWhpV1Tlui7x7lOJvnY
nLOIViMH8YSna+fT2Nn+F8k5GiDwSiQ9OnyXIttt75h8YarGbRS+PMQMoY6PL7meLAGz1ozYw6fV
mOaoe5tugQBpDSMs+9X8SVH666F/v/tE4Vr4Mj/D/Rkv+5kO/IDyEpKVhhFTUCtWpMZwgAwXNvvj
l9TsKi2+h/TmXUg1uhzgBGyN3TO2PXKACJGJlKTHdzdO4hmV6EnQO4i00ibOPUqomUYmdVML2M37
pZCx6DVoVvOR8owx/XkB5w2kzhjRcGUWha75aZx2FKAkjbkjdZ1UdIg3FuXrJt8Pex1SKq33TISj
E1uv4JpOb3i1dTrZXYjMev9istYJOr1uSXlXPbsdVZSIDpKgnBigZTub9lff//VoqCqXhJ8GkSR/
fQOy6y+L6Ep4c9RaVbdsoeDr7GAcdQK3gJ8K4Gc4f3aaEQlBJz5SweMyceoB5ru4nY1HHDYSJQ+S
KzGzx3QKb0mdqW0MPizppviYSNo+OpbpzbSfSrci1KpzMtf2kSQNeG/w5uvvyobFqiZXPNKWGE9F
VtuWhtoQ6zvN/7qG8RIgD9AORzils3jegMa6Uon3VwphHOVpvzAAwJPEqJA2ibnsY2tnH0bMk7pG
diwyTM3XlSSb33FIYTIgJs4kKOHEs8XlDFsM2hPPYKgzlAP+xEvKxKCl4GyB/bh5NK7Al5Xz3o/n
H194leKEnCtr30rXjxiw6YVQlgdySxo55XnMhNqgv/Os78PqzACRfuuGJDvar0WDiqZgytzY0x95
eFkhYCSu7Pf/85Cf7eOG8gJ6r8AZ19CTfPInhg2DzkjBK3Q4L3D+OvQ7i8x3iSBXqtmjr3YCxj9d
PgH46inm/x1q5yn75lWMAW6+gExcE+Wezq0FFMxiUesr7hSrg4BbcOsVif4W+hNTiqikNmGMInyN
6UcbpU79kgbkKzKJmbu731JyxfPvr2uKqOy4XQCVMJLjLVA0Pff4mv86Eyv2EULjJ87WkcQEFQG+
cIJ1NkyHZO1L/S4lj7bxO5GTlSdmhyog0baoRclYHh01iGlqVT5NxDdhqgafY8h9AGD/bNVT9so5
GPUzfXo87ORpECPXUG5TZhC/9NkgB/mQPdipygwXp7eyeDje4IS2BPpDbBnmRHS9Uk9ZCf+jgvq4
finckiNCJcYNxMJI89pC/lxB96TagcG86HrSUmp1KbM7yJZSuDwMeWNVCG4JqSs8w5B3/56v0yeM
AQ9c857e26iUutstGSmEMVO1aV2I4gdN+LwWfwfcr+Gu67Na4IDxGZpgYhtB84B+mDjy9d8Fv8H2
G3vrLfQQdx+UdVf79B3HVXap1lk6tRfUM5TKDkGZXmaTuUC1arrUqCTZrBtWE+ul5F4SsuadpG75
PvEiazwohN6AQBRIqyiLOtthQG6wcRzH6XoeQL6A1OLwsbpwgKpELKvawdfiNl0AWiOAEsyft+BK
5UmWGKXC0cteOV3ODV7vfkPygeYg4iiwA6qLTpqeQiwBqBREfq6l2o4mp3mczU43sSZHMmlsFlXn
Tr6C1v8AgAm+I7ycjxHlcTr5XvZES4knDUaNPxPqD61a+rspqyF76ZCUPEk9dcdv/FXbFeU6qcI0
IFi0PRfDhfRKvQonWkzmOeMlb+e4hgqVehWfZytb+zxLshQhL+DWMY5O7qUrzSVMsGTaXQdSH3ZO
/TDMAvx4jw5hbrSMgo85jKqypfmcum5HSuAtCE+2dSwUyg3961is7T5+QOb784ZERBLQH0712sJw
gmbajkpkGiL9bfWSZCFAhj35iy0VcE2Dz472nQIX2tYXLo1qh6l6EKmTbAfND1fCkUku3GPkPDyp
KpLJUQwjrTbZPAquYRcfH6RoCdOFhXjq0pBbF7fCXg5Rm7XZmys9klPbS09MPkkkKAjeG390wa5P
6YxlYv0ij8IX0g+2sNA7uZQoKYqa3L2L4XdNtObYoiaUg82M3pmfIuk/4u6+V+UPdf3asmJBr7Sm
K1i+DIAkTwAMyAAFKuz8+edvge+Sp/J7TlsQMowopEmjrZ+++qQrT8V35x++auSoirC26ZGQiFn5
cLT5OdQ02HNRCaheolD2fku90B6W4pFgVZTORVaBDfEDs5phAb43O7vTguQnblLhobRqZb7aCTEi
VeOn6aRtxPmUrKsBdIwUtGQMkppQsbufNNNnFFP/rhrd3w7Koem83g9MPVWpcxsO/bFnEDU6HCPx
SVLB+aa+zAG0bf3fnlvkBiZ4KDY+eoyprWMsqPGZpKq19kmL8yqedR4exTMvEDMZbuKSGL0tIYR0
wbaJM3hSOakD00WjZs0CJSnhLZ5mokLfH11yh7DapaEXA0fzvukkpmeIu+5fn9/w9FXNuwyo/HEh
xZ05CdGZrcDRU0CDVC3EPhg9YrzcNeFUNre5USLXV6xSS4nreTn0HTxqS9o28O1JsixbxWbXSipA
zE1NP+q2Ui8BHd9rmBHAHah5tsFqtDV5virfWpGtJauCJVqTiUp+UgYqSx6heUzfwATTbYBcYQEb
Kf1rr7ZsExNm9uuYqHAHAGGvCw/Uyb8A/DZ0/qNXpj4ezOKobH32jF1RdNs7Xslz8PCFT9rDj62l
Dt7fZiojYiZ8tkS5dbaJ5Oy4ZdE58X18GL/EpnuPvnxLfAbPCYNWjD55xMyTnEghsAggX9TSKgyN
BiyjoHfQvX1KhIUeXFqckaBjKzckTY5UB/HUmue+BgaUV43QdvPQOCmOoilzEr0utRKu9MbZClT5
YvVH69B3ESXV3C4MHX1qzD1dqDvMXkXNRBEQ0dzDUrZFdGSIfcfeFg/1VHwdj8ZfzFaWUWNG4d/2
Ur5KFXXWMsLXiM6BZCaa44AxtF7CJi60k29S/yI1pQM/CKTRQHXIHJ1a7lzc5o+b19OnaXlSATxj
c2nwC+r7lDW26nK/mEuDEd2fW+btkwVUY52dbtb2rFIEUxrQdsy6PSGyXVE72C7K1QKPxJwEL5g6
gVTPNGLYvwSjlgZ/HS9P2vovwVFO5OO9Y267amxsrehmlUrDlljB0t40RJww/xxlY77IRXRdU3sw
3JtoGbZCCXot0y9glf8xqVk4dU7u7ahfJ2WI4ftyhQJCVm/ecIHnLPJA9fc78T0gZIyGfShNX7UL
qo3knOoLGJ+wFvMP5qk0POoYxZtmf4LF5yoLv8Bpmf8Yaf5GKmIP5S0Ycag13se64X52OfK8oydN
Qxs9+sHtrgYByc4/C71536DsOaQ7HQhbbBrUN7sbDACDvnpiVgOu6pOVRThRNekfRxelMPJdRfkh
wEF3IkP1npTA6XEIXcFo9iTE7bXkfpxV1FRRm7OMvsxvqMkpueJp4k4hbK2X4vxgp1T7l2yk3KZJ
fVkcpKu5BImK3rLfU7o1mdRNNFR98zN9pHImaDjHhzALFfyo1sRGpJ0VXvzGRITsKwCI+ObK+jP0
F/QXO1VpGpCOq+46indHvewdl14fGWFJjl3U7Ma0X7SO1vitrEV4S+yGtY2sOHPnVcXDogw0uG7V
mORP/3m8T2Ge4DxecsILpRG/Bkx0mECHi7M/JVfISv5HrPt72sbH5QLINdCL4H6UqOiCMdyUX6gj
7SQR21Hr2eQMLIzwPi1UIvungGvRoIzr0c0J62uypLgjPdJK8xrxTZlpBr0WTwtuBjbw15TLQWwv
XDHLlqnG1BZvENExO0twbpuDy5bPIhxe39slKw+2NS/VrbeYnnnG4OVHXCdQIYX02e6HOHbX8sc5
um15LlDtNOeRvdwDsOoLdLo9u8lbABZ7MTorStrTYrMouCRw00j87oWtrEVPZ5XZpjhXeweBRmqb
D0kLdVfGPV257cojUklV0wMTyI6ZymkZH5oC2PdHJdQPZHcmmEdM/Qs2PX51zT8fJ0ZlA0k8F9xU
Es603vqWSsJac1OHDAiSu7MuKroUK9BRlvvO17csyJuJhSEIAF2SEETtR/pOtvLBpMGVOb1oNDhS
3f+taM2YARGsH7ih2SqJxJBEQjR+Vvwa63y9FZ5BkafQXVOpowRisPmkOXRZcxaHYKu3Qa/4KvgY
oENADGb3y7qU2VpeVtlZozB+099/EAGZn0OQXIgXmOgzN2SzDBxQ7o6VXrh7S1d3CVky1S16H1+t
zoyVHAQuNIQuDyzBOKxpAuBSalIuqbl/u6toWVWKYa7Gjbs5O5TI3ilD470TfmVqz/l3OfxmPnGH
UV6aOPQJ7jgGYYML4PgjiaIVHbsFRdi4OTgQySf3Z3WARpIGFojJZaxMzCPnO3xCs8v8ohcewO/H
Ww5EEMJmVal2+TSLuK6Z4hd03lmAw4VNxvgLlRFTWW/mDP/1acAwAeVBTsmKX32qWrORtqehy7Ar
3nP9VeblLV4cO3cvZx72/lS86ZybFdAfaAIUfAs3iqWkHANFfzDghurH6LIxvMeTNoQBe577WCKX
05Z07WSqDFK4YUZFT/Pw+tfv2fYWNe7ouDbyhrQfHaS+/OeUpilnNBx6wN/XH+MEalesO/eo3Mzu
iqhpRb/gY4GxhVSXzumruPp//c9EFaRtCRrLFCkHNdNIQpIl1/v4jLKZN61rF6GchyDv5H0sQ+Hw
qBto2JjC676Y+Idzuc2Qko5M3TAVqZNkzDt2xuOwROtfhW0gKUu4TMP7uKBk4waWdsH4pHY3EsTn
rz1ksAq+q8NhAR0Ky084ehO/aKFaTvVzItJmhBCx07hmjPWHVe+QnaCSdWgBLouyL6W19QaCi/oB
pQ0KXnSUAYMSfdAYc2La5poFKEeG377B+aJkGKKi5JclLCf6aPblLHMYp/LZB2y6zx3pbeQOFvua
hEsPsA6D3Go6jGiuYcHMZuFoWSGh9h3Oi9+Jq5Q+tiEC4UE0CDR+PZzyvKth8YJJgBuTpbycA2f9
NojN2SEhN7RT/WKTjFSqkZmizqVsRFTAua9VWzQL4Ay88qBo349rbH4xnEZJAKbZ6zUK5AaHS8Ik
/1oGRAh575KpnaLNcgIMJBlxSW+Ff8ozemjhv8eU/K2AyHdM1oHQCTepdof6O7TTazWEEqqDHg5h
WX8od0kqUr7fEwGDHHvJYMKVpP9LUKkBoETwWbRx+tEFEgGPVSjN9lNi6BuswTVJduRg7YKiivm/
Olkv6nL9ebO+UnX5uqWudItyXyq1qbJRW2qAduEd+F+qvRqeRHFyWYogs5o1YR+llMbtxKYfBEeC
hVl38Lofgb0PacO0xRNckBS0FrTmUIbVqH5b6gM15yFVYV+/LfozbLbnN4bviBBaTVAsVU+LeKJ+
jqDt/FVND51e8T+KqhDS0sxEcVd+SbEIBbhBCzs3tuOAdCr3sHM0lapiSwQ3TbGDsL/nqRm7NtS6
uqSoH9aAHH8FSAO3Mur8GeD2Wk+ihva7KMR+YoMcmHuxtvOOHNS/uBJSU08n2+bwWr8gkceBhD/V
glNI8bbueqCeFMJ6dySnv8mge0iyeqmvZadEvK5hEnoUzs2a+mSYvT92nm3XHl6kIb1JZyQadC7h
DafcXkIuJSCng43vmin7HdcXmCp98w7DvUg6L1rv9NST/k0z+Ula6JOy7G5mtAfqASN0JEsIVh/I
lwBOFdqRTIV1L23OGyl0Rtzry9Q2SiRjIpiKBPXDdCOyEU9mcNVI7TJMzWfH/K9GizPDvYJh599H
Z+e9+Ngzno+uo5V2aD6R1ZN/Kol4qfoJWtdO71GbD1g6vOpRHOB0t7NylWK6RFWcDmpKUclv2bY4
9abu8wybxDR49kxVeBymoA136PE9rewnUwxRnMXxkxtgdQh1Px1gBtMsGotj+LexPzgl0QrP6+fr
ozbhfEMCAFZsKVarxDyjuGYvUDJXDiI0xYss2M026aazD2H/FSmD6g7nYq0OyN9roXwHD8nqd/ac
N36MKsnSJe1waAY8meQqDjmrsfqD3h5IWlgMwuwkcJZZbMbQ4Ds7Sz1ftIN8JsGxFOXtUUG95FYZ
GucKJgDW8ogd6Yapk+cnUQnTEfW60+T/OxjFyP7wp9mWdWSVWnzR/QR9cT3YG64ex3BULxBLNN/T
4JiAuU6o/3f2R2cIxCaOtpfPFUZFHlA7Tzj4n8OarMi+iS6nYIJ2LIkkQmZY5626BUC0T1vEnq4O
u3YbyXhg741wdVWkTBlCU0SMJaC0+cDOoL+i5vReTUr9i/B5ffLHrtrUyM2XeV3XPzNefb69+Zm9
UsAlbRb7bezqOKIvJOH8QD8mIPRwG4A8LffkdZu2vLKyRKoq3HezCdlQYJx6CZJFQyg64cudcJL/
60ycLj6rh2TMygbzz9T1X3UYrnrHsvm90TjdOgJ46JxVs8oqx5UM4hDgdySlfCrBarw7jqeYO/22
daLnH/B0Omkz+PFhJtNJLj/hjaAsGRFhcRN9v8GMNz4nxb7PgWlzUs14XANm0WzNq+m3wejHsQ+Y
aTSzy3MuTSIcGsZ+lGq/QPusxxGlMxHc2eluifc4sYITcra6RIrVITLhrN8TDxN1LLOUPD0zQfQB
gLyIgPTBcnJYV98WPFnz0L1+kArm/fXKZkcV68IAPiOwvuhF3rSFbWBWwdXr4RhfakoEVv6Uuh+s
0CZxE9fftkXyuzn1Y+iVeFdpRpD7dpATFHMSVbNMYM9m/aeq0ZthecZWUKi36Puv5exRT0nvg1e4
U5vyHDEwVYFcioSADdv3/KbljDHzcw8T8qshZsQzoaRyqZeuT7Q8kLvcMZVnejs7Nf5M4BL4P5HV
ab4uKm2kellYdghPXuGo6RM+rouHmV8qAg+XNvRKZjC9RxWVpodqkHK6WrKlWN4OtGwrDO5sjnc6
7YOjWpKqAsY2XmvtUJ+PM6XRiU8fcaarxWmpZraDfTjaUnLUJjL514RV073SlLFZiYOVCmB1DgUM
b2V12cgAuXQE0oOiNd27xMDqvwktZBc0yORR6zFWD53cjXxyt0pSj9ox0yD73AfKwhA+IyqwzsF8
tYd83g8INO1honXWCBEX89qKukGByqskWKEdUT7Sgfvav3ftHwofvAL8Ueax7jin9lECsJKXtdDW
Yezxn/+N+M5fHpNd6lvZVYja3+rFlxlf1H58OvkOL2ArTEhFtSxMT5BQ4GuBIzNZcsZEaMmK+e7I
MQ0xk7i6w6TL4AOISQ61H8LLUlhSDV39hxPsPXwzWYJRlXEi4a6xRd0qDlC2vp3EfPJxpM7eg1vN
bHE7cSwbw34JgvK81sQ4x4OPis71RrVcZ5IEX5UnCaGpZdZWWSO+PKZp+5lk/Sd008Ak9LKy9gOi
aYdK9XtNXIfYtP28sRiYhJzGYJJT2rpPR6BFX7LXwI1cBvJtUlYMa+wRWnEe8ZvLc17SJeKpK4vR
syZqFJdPolUVQVqSF/qYzFCk7DHE6b4HJL8yvYo1FYkDWjNeYoeuScJA5qsGeeun884AJg1k5krC
xXcd9mdlLmlAC7Ld/MpEknVdwF8A5xaI+XiaXFJN9Ue/cZdWHjdMNuSRxRE9TC5a4ncAsoM+dklM
PCssXHC2GjOAI1oMvbEKqrksfRNLCezZ4IeFH2faDqwBGSav465RldTAM5a4HzE6Q4jj0giE8uPm
mygQgcTzA+B6kwf4MMDKjSOidst9z8BqQqbdGuMOscE68IMroLekDgQ4GRP/Zp2aRIS/qy9KsYhj
sAAAXzr8DehX9NXCRxF1cyUKgMcXfLGfqc/rrqzbxyeljbZnBWpFB/vFTBnhbRN2BaVIlCBMIl8S
uVye4GxcWH/W6hHawYzOLYF1C4OC8+F6s6H8kVNClmohQa2ykafnwZRc/pi0FKyZh//lhMunnFgE
bDTIxPtQz8/ABG8idkJpz3NUTB7DykrJpeA5+QZwD7JVbHMbh/GUfE2xDoby+HFOCTg6cCS4Bdgs
rbwwgTZgrh5CnPqTBrXPMIwybL22rQG3UkuvcC9W9mPuyLKdfFpoPAPChT5dxTHOMdJeBkLlttXB
tjMhHMS3cfRZfijItxGV5+c5ZajSJAW3aM+cCCD1Vi664+geVhlRoJL/uPA9mtdr75kKW7y+3any
RORjGEJ82Q5uXYoV5D8QaSZPz+BGTwHdiIvnCRjNea6VK4JPRQA1oFAbZGLWjHq4mKJOvqeTIa+O
SFEKxjTcI2518Ln6ZGVjxjUD5r9mRhTXOcxp/RsrsIi58q57fU9yXOj/8e1HbVAHJ+YA1xfA1t9b
enVJL1hRsDFuCcUo7rLZntGShhTm9VB6KAGtrUR+mS9/XQnZLTfMYPkPhdowJ5awdGjjeKhpA5HU
evXlO4hwZI08FLQR2VpuazYlt3Nib/TmNow8milHz4rNlt/IuQyCjWkfa8rqDvpKeThHd6xLTFXN
5dzbQA5sf6kL8D4BNk0pgfqQ1BA+gFQe7lXawNNxfsO4UaUds2wlJage1RGMSwbuad8KcYUojVdi
DuwEmf6Wg5sEMWZJt54cf+Egd+Skrpo4MD4kI8p0f7IKGc6J0JmeX/6yy3creV8vOhh03ZiT7e1c
LGI4ux5WLLHYqDV0xcEGEf2dMD4AKxtcHQiUBvrtuPhMS8UsC0MP9k7T5NAPto98BngBAqCv1m2o
c04h1HCOmJoet3gLBSHfTnlDzUtwQ49TMPd/jx8ybk4kWgCG8ay2zB/qY8NyfB1EKPHR+GBsfKxJ
r//LvRuxm786a9iRQOrLSRpWUEMa/b2WabwzqawYkmeHXGqLp2BqaxzPWmXBokcT7PFg8KspcHCD
R1PL+Nuyk3v8HTDvjjfZ5Ds1pmnXz6zghNh0MJ8NCRrZ2Zaw9IQVQoh7X2uI93fOrtZsg7coA5Tx
LgdJqv/tQV/eb3wlg1yGvfRqYnP6NLNfKvfttDF8UF/o3Yc1e+brsaH/8nEu/eiUf0Qv7LJTGXf+
pLcuGdNLq2lETxKd+RYRPv8pGdpJs3jAfHfJLLs3F1Lv823rKdu/upETudoE7PtYndpmIICfKtsE
H4+a7uGv5SVhaJ7tvKY0tfOUwNZv+pXaHU7Sma0oer43t0byz1Zk5bnEC03FayPY802C0lsDR3/E
DNDVPU3TElvjxukK2PRkS9l4B64RscODhQLfug5Pd0z712AeCKmki0QQmGXgUNUANwLBPQUz5n1c
u7lbt4ltoYhrteW2yR46/nDOxyIMZAM4vyB4GpOYk9WczS5baPbULnZT/bgLPqkqqdC8fj+430Na
hAyapaGxMEa/aOOWguex2zJDOEJ1WccWn8QNU3B9d35E2NDpTdYC+xM33gsmihVj5zYMwD+9bBRi
XhX6AwxWnArIXfAnPfM23WEwiLm6C/gXx9c3i+nQ73jWlfLHntoNGBw4GgEi+l3JI2D4VuuWQFJW
kwZp+o7zy9To21R8md16UyUy7R3+EtP6JJ4cM8//f6zIIZZpxASyHeTZkFgaSzDInVf/csnlXczU
egi97LxBF23dGjhgqkdknQUfUQ8tGT9CY7zUSAycxoa4WgNbIgvY/JYKemtymghUeHVivYPPOgIu
zbsutKu8+v0NRbE9ZMsA+4iaYzYv5t3IPDT5SJUhSqwYz0gKLnGiPMQvYOERp0NZ2KTTwqSwVI7K
G0ASkzssNM+qJgflVvykrIKBhf4la6kA1r5ShfA3qEYA/gPt8GY+ycJ5qHajBDX6afgypY4x/7j/
JhBw76Leh6A8SS7LBGR1mp+9m/fU3FhKMlOUcTATgSsk2nCJBYOhBLoP0T3VEhiJKrzdFH7egucZ
Imz2BA+xmhItqxbHiE8YmhnFDPa8h1d1z8iAje17wsvhaDcMh0aJEeD3harOOt/a4qfLGvTRnir9
XKsqwO/39w3mC13JrQ4JPyx2C8ksBqvkiikpsjGx6ZOmEPooa1Ps2yH6SwY+ZDfXU9LcAixZ/1UR
fzHGK+yFAkBMofjqX2VJaiZN/3AeWSI+FA6HSa4YgAzRi5RMXsPXmezvzfXJA9/uTNp04QLHCPbz
ae+x3IU91iQPQzbRLgzD1Wx4iwDDDZtoFzBvhV4cWHDaEhjb7fE4+6XtdJRnUp9fayg8Tr3HZSlp
kFWT51IZIb00hEASSpdQd1MGO6pFMdtNbmFlAHUCgi9mHF6iK8jWXSbNh56TeisjvOiumIwvdYRP
aDwwBnKnRxk1ECIDlYy8w6fQDC4syNcdmwmrIYG7k9BMaw/NNIz+9Ofn4ry8KFyLHP0NGsWw4NTC
wXaNwLenShPnOJorm62R0EGcpB7xae2smCubd18Kbzs+hyXiFzYLFS9flxsYlvPv/2IU01lUVCmt
IbWfxZVZ64Vw+/7sb7v+eUQP7rZNncFP2G73ewLMonpi982cxUjdV63vfiH3LYSG9hJL545SLGVP
IYRBmfUW4mKrsNNel7ZqGyjcRmGrZCsRoJfIlJX9lmc9x6Fx43Hii6NfiCMxtHP7wchOpPLArvR5
dK3J14JJxKdM09RiTsGNpJtZPsz3NiFMxeW3n385pwqDQGirOyOeAR+kg/TobSlQe4fLfzR2D79o
c9hdJFbF0TRGaPtjno/ouWFiLqmp6cmzwJ4j+7y1D800UScs9JRipFRuoNmFIFPXkYCJh/SwPmy9
dSA1GynbeXtcF8/NsTVPag/hj5mqBQEY17/UYBpvlOpjkR2t9aqFbi9G+Yw9tUWppwdE/yGbiWBZ
E2yKxaNYNzZiER6VZJnrLp35ImTNopeE259V41mRK9gr96+oGk7G1cf2HhSA1V8TXw0F7q8I0AQw
ECrC2b6dPrxr/yN3UmQbn3W0FzpwwnRwMq0We6jgBu+RFgHoJiWN9y3v487xuGNG53hJ5+/VE40w
88OOElxg4cBoxgZLRzVTx6dAwC6P7GPdyNCuDA4JvzFlMguUEPAuZl4jXXfjrjiY8KpiWW+KcBuq
E9/vL7co28tCKIC9dOe1s9M43YTv96TtIvqu1FNQ5IXFoIqYPMvZJIWtfZMD2B48AwF20kSLSfKd
VCMkIGD0jeb7EyO87SjuA2NluLW3rS0U+3ejQg8PKXOjVPmeRQf/rJTM36tWAz6iQF+tcfiDl4di
YZkZ/q/HXIbuQCfkfJc5OpTjJFME7xEvOWyBJCy89KLPxJKGP+gnUAc2aYNiTszUHeFkVIJK0t+M
PkxBNqxeM8pRbE2NUrQKe1i799nEEnWLnSZc1ItUnDhhPUbHqtvbDiQkPmF4/8DHm+bQPqzC4xb+
cTXm6bdD42MoAZi4gCTM6atItBHWkLDqXxoudQjaLhMtlj2Z9/Ak7Oowu/wAJ2i3S/8M4Z0WdIuB
aXjGFBZmyC6NtfidrUhwMjmvnMh46JiSBB8CU/49b7DoWIyfzThVIB5p6E7mPB35mikoYzoWzu+v
zUqD97/5VDgxebdQ83jBMbOm31u6hSTo7qJIt8EGGjs+/EaeTUFuyLaHODtbPiIshAqZwOaWSFdz
mjaD+UVpjs2/QzqlCeOnevzxWknhBtGw/iYZQbjc5g85x2DQu6U8townPfL9Fm4ywU38W6ApAv3T
e3h4nGbvB0FcxeX8tRtWBNPUVtnXaYp6RbKVROtNBAAnbaECsNlmhWXDFMXs0AHhwFVF2ZLz/njy
nTE7K5MQOZY8GZqGVnFMFm8gXnfejHF+HnB+RqVx4ZCE+S6pB1ji9JmDD0tQtcNz0CkFGu0BP+Eo
hEix+hBGk0HUP4UOXij//+/RGBbE6CKdUbBFyh5Z77OWUXNsQwS29oUuA3ZppAdAMw9RNj3McXqy
MnRV8qsRotvw+n9VIHvnB6FfCLqwR0O6835eXmHPGEbnZhEoVl8Tm7Bp395zUte4qOpaKirsMdsQ
b926tqFCxHHcTQUXZMVMk/gRCVXWu0OYApERRoZRpdx6iwgYRAStRR41QAS+gVyrRS60gTg0XRn9
o9vadugvK727lHt287J18kQCvtjObxQOpA9HvTThYvrtWp9u2NPlXtoos3dcpz8SOmz5XgLH4Tvv
ADrsCJmp/an/mZmzJ+WcLDRi9nu7BcB6LxYKs74i705idJwoOFMk1uAP3qarydpQ1jrKAZmKGai+
yhW4Tv9qFTBKKjfzrsL8i4RAqDPnQ39BTrMX+eB7q9n5P9aicf1eUU8kK4qpPLJrhSTKWRxMci+K
OzO1G8jws8qabjDi3ALjApY+0DPU235+Ch5hUsNb/P6kIWow4IoDhyapaJdxtEvXbY6KFpVUwhhd
wu/YwEXJetf4IK1cJlZRMl18zeRq6B6HOCrGbxIjiC18+4pvskQm6oP+vR9qcsQ+SwIm2Bj930zK
kdqAo6LPCrHv1CG4aKrEnxJWZuK5CHazoPYFAXit0V6sn9hUQiPcPy9xuAAYzBi+40ymLBurJR42
aHzsZMUGid71rCi3JWOHCzOMNGVZzeuCpWt95Z6XF7HveviLh0qGoRJ88JP7hw+ey8KVeUW0/kbi
nJzLCAunP4YvpSX5yYijo7pNF/KvGytMlgCBUH+EcPvE+zTuDshb8nq5QBMo2ue2llgULyexMbeL
qLPcO51dQ+h1tUu7CdEygkl4pYuDSzafQ5y7rrvryvSoHmrrajZSkLrmbEkH/iRnbwFQEKJqtUO4
DJz/KJyxnbVC1h0eKmgL0tmfL3cXOFdLTK9uM+BdLM1PlRYPdfdw3r3xdgs264yp1vlXCa8D+RVV
Xlt2rZqVgcNFqj5G4+RUh3NPbcB43/H9Gr1GTAXu1NdLMZfbfbxWGsMT5DqBblx2IQBZmoLe4550
8I/mPuq53PaVbFQXfK1DSkWM0fr+1PbL5M4qM3NqWoSk08kd0TUhx3cyB7AyQMkO94rUT+Nv4vC1
oCb0Rv031UgoOqQYjuYelqboT3IsQJ7/h+6zd/r5920f396S3y1Vt0b0KTinO/gTBLLvKCo4g/mi
XdGF3RHhppR0jf9CI6cPZcCpeETYvLrM/XQ/jvKjQeVkFbh4PBETGKRhMpXgWv8Zv3AxlYTiLS8J
t42uOlj33H0r81CCoMtj32Cfk7xoNZo7OsW79yxuMQYgYn2EgAcpqypCk/zWhg9oT9mrQftDrZDf
oLoEkg1vedyu8GiElzyYQHCJzZo37wSC9Y2vsulm2fX3Jh+6yGhNCgp03TtJ7V09LLZSA+WJ9GIR
++mL5hQ1iBqs/nAMc5rvOZBXa2Des9nH9+of+HEn8osy3iNrMFSvPBRxWRH8RUo4cx13mEKSIcLR
1CNuSSNa2aDP6Di1+dtF/RZF7j5SLOjyfCaQp3uhoCKu7eNXTRhbf/F1Q95SBtkiNeMwckN6Ft9N
8ZfizBwv5D+N5UjZycGyVXyhgp8ZLp0nm8n5Fwmodf11BalmBHIRQO9q2zHCPeIn1PVVebwFyDhj
DLlITGkBuwz2bam5XFY/Ce/o1KVV+aoZnXBSPpmRxHG+NrNoKWpNyiDiYun4/vmMxRiYZQKADhdr
e3GGLLMr0ZDctg46JoAqhYz9ysIGi5HbEyvAvdDFpJdCsTLaGF/Hv2y121d3C6o3i59O2DqEJ/rJ
afpzL42dVyeBW8nm3ksOlsK0L9Axx3+OXZ2BdvDC3PWQOdjpdEeIppTW5mr3wz+FSfKirvy6iqUy
G4TIKFNjAG/7T3Wn+AYDwV15Sf65/Npw1Zvi+5IqyX3E/IX7ibQQfjR0MRZsKmah+aeabXEoH+yv
pz/X21tqqEP6YnA3oIECHLTXWJPX5ufGKCBvIYgzqxlql6UPPrNp3Kuy5s/4R0MLf9Xcuh4djXgk
XP5qlgyBFejEbCuIvjLzBgSSiJbJtKEuUCg0Pg5tE+UCE79trh/CccY2CTrCwBW4sduWCa55NyRP
SsikmTUp3rt1V8FutYLRJLItnc8MyHa3jHh8KbQfU6PlK9YMk9aIX0FHb4/QftOGX9LEQOszc0+P
q3mPeAcRw79XQGkNnhELIZVAS/7Ubp7yHaMajMOKAshUA2L2HXtO59IMu8PVCv+6myq5fcbqQFps
xHHtmxotE4T5QOs6f7jhiIAA9d3Qtjl3KjKYeJJxvC7ywOWggHxFZZPf77IL1Wts5YZmDH4sXWZA
nSx0DjQMz6h6bVnpBgE6+iKDlWxBCy9LJmov1YyoTx/tzsKlI5X4m/3oj27RVi6qMbfBLN7sYTDi
yfnaAYErYa4tmQd+XglKGusdf6XH6a9PM2LVewyV1V1fge5FxC1ESQhU6L+h7ACA700HHt/E/dvI
yCuUJ8NYDkWkHHD9XpAww1UlG7Ugt5tkZHQI/CfsgSAkv50QXCzkkAyjvbeuMXFJLMDOR6xPl7SD
r++ssGVTXFVUtrg+RDWx8RbWMnKaGjl74zlC8lT7n5orGTzDvyLuOz5tuR9Uf/6iYZ38QHgW7Tfa
IuDGex31vGAsPWa4dR5zBrObq3xn/e3dcDJ9dIyD0a+okHWScx/97MYImg2w10T5SNIve1jJF1eI
OFKxYk71IbGmXOXi19hnVlS3FWDPowO71X2/qK2w9Ods3dXjftmDnfYaoi6hJwLBGfnMXRU3w6T7
SEnjMCZZTAELWgDescKdVaBpbJRKxqT+k4UiuhQzDAu3ZuS+JKQIoFGBBV2IrGab7u+8kwhDyExg
/ipci81jcYRoROpzpzgzvTKJGmDvqg9HmJZTkMNe3vlxV7PKyQUlOkIKObBCWAM7t+JY62A9932U
Yb9cwrsQWLXQNDNqXRDtF0oXfaWtjh8ihhPNc4s6o6zQoxHNeHn+S/SPmY8TqziQ45pE7hr4Xm44
qu3R0sYIVKfmeqZ5FHicCQPuAdYJGyj18QBEgLZTk29qafBOJrJL/0FobUSbIe9FLQPH4qoU4aOu
Cvm6w/LcUSJZP4Pg8WRZPH88PxJs9ZfjriNeDXlWKSD38Ck7ZAsnVWqttN8H5glHRoNJIdAlUm9m
vB+tXyl2ZHILvFHS0Abyk1erf1gZykcayL4xYCuCXz8zEmjcLR3SBUKMOf/HZxABNE6izXYBk/WD
sHJkEUYbT4N1hQizp98RvrcYG6orvvAT/ZcFsrgrBEwSqcNJVHnqgbl8HW736xoHLNpXNR31axEO
RUdp2b9XV1mVsJJg8Dc+ZKyDndFPwRP2JsqxH/xFZ6GTXG6dAqAuiF70x7uwJZzZx8EtGgK1D8zp
7/kEUqci8CaWD5mEOIaKpxxJ+iKSFIT+gBKptYCCGpV9Df5gQDcyilo5qt+RBjpxbWTa7q5X+DAY
0vC9r0yRaXyO8sw6p1HusezqWvI86/80Pl4Q7RaMKeLrg+4/XDn6A8hvmyL/Ax3mUjpstNqLOf/Y
+4hLtk4cTouTg5spZS8HB192jyrfC0BQhRw5/kESyXQo2zLTWz1YKDroVZDagN8adIzuGf2pRR3d
cPzC1MV5hXpfjM1PJhu9V2EEdweov8i8qeVIxxRjuATsxVdaXQ2JOY8m2pPSgtf59bJlvaDIz31U
YBbZrTDF0Gefs6hW3qdUmdC/JiSZLk/TyeXQ2yFZ4BOcC0Jr/ELiqnazaAzzMiWxypqnJiw3KpjP
glX9vdcZMEBbMJdmoCK9RnPVTZd5oYUKwPxj/my4gB0nLcqN/EKblQfzr1hg9mgsc7dmZzgM7D8k
OlzBjCqn7pg5++5+/lRq1zj94TtWEVOxMJFJo/JTKhP6oqkIGMcGH0vk5nMJBkSjAWldPw+ws202
eVEFIr34YINAHPPAKKjNrAIsVYgDjNd/SWcbDtniNf3FLYgnDPU/xWK06Rt9sye0qOo/KT0joYxR
2k7uoBCtTYiPq/uIqNvvQqWK22AJJnACeS1aXKW+/bypUZWmvu/eot3pQyICurE7yc40K2rfSOH7
mqZC54Lwc8/2xruHtdcuHDtiMyQzMkN/kOg3PfRxs1n6TR/dpQ82HMMpgjOM1Gn62BR2dWQZciSk
fB8IY8LwMUO1ua1AqxyL9jcwgf55Llzlin/cNwhDIYhOE4JKac9EOrsDHNYy9GcNF6vthpOixNkg
Wp9ZCO6+cqTqmNpRuOZEIs02K//NxH3r9PfjVuGESG4b3QwjV162RZew6c+f8Hor2Ss5naNHxqpc
CSW1kPPXcTLgzUpQYbX/cZXNfc/Q3NHblnhT03PUo6kZCyGyxsf/O6n7vm19kT6/Vej0F6o4tBA0
Ia7prO4fnwpM070CYkXCZqQX08ILIiEwqlQjSQX5H5OJrI1Z0b8l3MR5QuUW2v2wRpzjVtInzHcD
ZDVZHIB57X7CL2lbZDakGN32x5DWL7ndWRPpT20/BJJA++D5nnS+tBGR5XtUQntGJuh7Dcn0BmFi
0sGhflDQlnvPosABkXhElix6y1KnhXG0q8KLDwEePx2al5d8w6o+bUhJb8jLSjGQu+LsVGxjoeZu
3vw0tfIT1od3LiFxqxKqFxPURn21qbyo9CbvCNWKfs8yTMJGErrtD52nACzg7P038oj1WiKURRDs
36t6D+4266Oj0qd1Ve0Pj0M7rY1iJryk0Gs2/LeZEt9Qe9IcL7nNpV9ns0vil7tzEg1YtuQApFzj
eWQoHXTMiBidtInj1q2CRfpbSSlSfNLTS5XfpU65xKdf/4aGHtvjWREmCgmQwFSmwBqd4AkoVxmF
ZNsJ6CsfbBUrOStduwckYWJGsaFIkkqfE/X2KBSxUg8qyN99CKrJfhUF/UuGzCSTitNi7922Yp7o
Upwrnr5gh9WRK0sok0qp8EAfpWwt+zrkds12M5d0K19Wmvpk5V0wwF6Jl4r9EwzIMKCAXn357Xyd
FUg6WElyevIzEaQ65jTYmhx2BQar2fPYbK+tepN51kAOy+EG+zV52KP2v0w8b4/DzTzw3wUHlSbj
7NnG6PwFDWTIaQzbUrRP+pH2ZDMobE72YLTxMXWSBfnLqrhl4Zx7vHo+z2JnG9TME1dCB0voKNTR
kFrX6iTpVd+9iOoXpxKiN8DXUYskXATv+EKiCadq07SiE5j538TBQCXVDQN2Ren+Z7fm3Sp9z5CO
Ljza4Kl2Op/tMYmd2dU6Wgu0ai6syaAGtz+bkGWERmdq492sk1dHIo10vKR+lKP/p1J7hQOx7wCp
5pgmFmX7/tdJYvF/tQpMLuvldKjvjvPILtZwLoBWkYCqPjlXW1TcLNcocRswEtD2CNR1Yv0MOK3l
Z7nkrLqylK8/oSdzKpIhVO2OAl+57U5dTdg/uWNVcLgJyEpyyZOw54bH7bhpjpmSbevm6k6pngQr
98LotpJItNGvXyx+RMTA4GQtze4d+AVkLG3wgEhzYCHKrg0kCai9QccBTxgl4PCbfcbo+Q4zXjWk
oMcg/DjO8cqeM3offz7unpH4AqYX/4nvJk6GFH+5Iy8Q/xm6B4sPGpns7cW2p9G6a0ejiaqmAdAk
m15XCn2baRzq+xaLn3oGVQ06WNmX8Q3jgVsv07B7TuLBJAjAqySdupnRTOU2QxYRvKgzhfB1WAxQ
sYkHs0eM7JHXZvYxGrmHsIywH0Co8Q8s+6ia/e3VSP9JmaBO3ZvG2AtMLO4zUAHtSFy35HuzyXKa
EajuEDwL10N8B/Nz0PXHwelBXsacz02ZusuaOq6CLrJPbi7m1ZeCFdLKgNJlF26z5VVQvYLUfIoT
6jKWZFv1QlwiVCVlwDT2cn3dco3jXaElO3WWwlIBqEuMglWdzbLM/eSqA+P2n1lcHodGcxuSIKDp
qEpLNjR1q3yfO9zTryAN8hDrnS9fjrHg18zJZv0DqqUFHfzYF6m1CptkmhE2ZtMB4pJLt6pwnFPM
CIZZBy+R98M0FwKwlqyliG0ErM71fSsb0elWjMM/PwCOKuD+L4Jv82JZIKJj9B+xRlPHuquIdZL6
vpwTTnmIVyzRvfKHNblAsbBr8OO+b3OuLmDWPVg4zv9vJZiZSbbKHI4BtaPeKd0IzPd4Ripf/Hyx
I4ONmiWsIKVjnkN78XWOYswFn65wnt7pMr7Sx9OqYD5UhORZLZcAQfUJ4C+tnqAdoMDXJXrJ0969
m/IUN0gcSw45Lf/MF3lavdp3Yv41W5op8YkejBueZmgXEGkcOp2O0fblCMf2ssvfsSy2uW7+11g0
nYDOJflV8aVGqbp4sQSAeEky6aV6R0EixUK+eUq2EhX+27WgRF1k5VI1zf4KjQXZ5kAoJzL0y72l
14a7pUh1ij9a4czPNkso8nTGvyddKglDYGIsSRzKumkoVIucuo7/GrXAc8YdRev6FN+LS8woDSqa
r4tmpeBJ4jVn81eBe4uBdatRi3Tp8NYKrL2Ijo8kNHqYihtWA/rXhq1UTiqRH2nP5CXgWT4gCwud
8O7XL/+Ta0axZYH/Q8D2Rx8JSXUqlTYixCV2jTRgDeax+MxW5uhYfIg+m7utvpwjCHo+EK5Zu0MT
ebPXL87QuRBLfcf5eNYnjmdd1MsQnDYBT45nBWD8gUeO+iRb6MoTp3b85zTVr2iACfrxIgqiZaCB
Kdlv4Tx1MV3JCiNKom9WY8m1fkd6EIW3CSzD4RMpgZz0PN4n6P74kLASIUGuZ2ZkH3EEPUYX6tug
v3TaKUl9xamiLTRuV+1QxlYNGmnXEwi8ZXarUzzEAwcAeheh+vYtd7iEzlnWVJGQAI8S6WkYs45E
6js0wEA6sd/v1/msSBa+cYyj+IJkAFnArQFxi65Lmfk3080U8WH6GHCpc7hb3pu6QV74Y+ssWqNv
fzG9RM5o4Dpf3q7UYDQ9rD3nd0Uvji4GcmAcW7FPhw6u+y1KWcXokQkWyDL2Zkd+xs+pt5G504tC
aRcCiBGYEbxJYnyPpMWkbdgXe3BdKZLpmHOAQ+p5+wNziAZkNHlx4gvTRQfSj8e7SBSTnwKPJqMA
fX9JBlhD9dNYR2Homu43ITBa9608hBOBkdLoc83PfQDrL1SCX6smZodzgrcYmGG3889I/pG1mzJs
zuP/e4iAd/Y5inrdl11VDarDC/jfLbkgUZz+qIHMhEvdoys278ydRc0mv8OWk7l5VNImFEaNvKgw
AxDyYL9zRFVhsWCqq01q9X1nLjmqGsskrqZm2H1AdB+bMMVJgC8VYOFgoTCmri90YezN9B+wh+bA
ExhY4x+JPDJ9GLnuw2ItX7xrvfkstVCaEhK5QSVmuTvDDIUJo5Tm0VTPPQx+nZrSiyezncHUgtgY
s48I0xmpnqeYiha4RmPWWhEd6W4Cr/UDAYAH6nKbbT5Iuv7eLvzL5QjdMulDBbQ5w2DUzW1q97sC
K+rQqU25yA1n0aA+ZbFpN9hOBfoh8+O/v6G4Apn32jt6UuAOF56OoZJmDeDD22DAPaoBvm6vmXjV
4C6ry8MPqVerYg7AMN5R/CgxviaqxSjN53Y0hx/csLcfuUcadK/5jnzUUhcD9mwG83SL9uSfFwiB
mgVX3hKNM9dnTByu8fhFB1/nNW8JpFN2f8wHpV+TCAF69DAQcqQo896OmGkpTa5lahLBWj+YhgkV
uLHKOsVAltES9LnnHZ6EBkaWF/vzEK5P/fCMwEmEmwu2a2F3pAgBidhGGf41dYDKJwRiBH0TEkIT
bdylx0lcaGuaMUSrizB5dHJ+zubHiYA/WuekZdrXxh3ijgSjXXs3H4lk6U/gPIga0oiQ4jpTqnT6
LtqWK+IcZHTC4a6iAmxf8sz46iY2J0Me+hPrHIKvfqTg8Dh+DCd0rzzVVJPswQod0uP/c75K3FOI
OOmcDDw+qMKulqHQgv59eajQ80jJQFKYqOYIISzV0dHDpWEIEfdPPnr3Udt2JpP6Dsp2hRCp3MOr
lBmsFextWaWedgQl4fF7zWWU1kW8kgAxUdHq8+6UVbYjdUx0q+MkB/Uv698bnEWJEZ2W5U8Q2yU1
OCX1BmUWJzeb7ismI3fg6nZw4f/djxkB07Q8TmCyHwTvFoY0RTvvG7nw47g9FsDXNjQprh9GMLda
543wjHwpLK2GmdZ8sbh6K248guIZVVK6ZN++IfzmSOCxWRkPRA6Y5+RWc1C09C5J8llZnE+hCE+q
Tx7ErYpMYNN4GLUcDFHrdnAJyvzxyc2507Tv4/xHnZQObiKqkLfBoQ/0KK/hgf7Kt2sBZvEWSwxm
YbHbq/6RtnTnvhHYhVhmMMvqSKMa8mVAmOWGSzk04wMQaFv6s3VuuiWJH3CposVwOyLV75xvNfcY
kixnz0PtnsYidJZ4DUnJuZ8CgFXKQIIInVndAnETxZJY+LILXQR84cQsRJF6/3zGBYI6pEd2MNwn
v0hCrEPuB61oTa63PsM9KMQIs82M79u9ifayWJQw7BiFLLGH7gfM6S3PmRT3P99pRFfYzx2fdkVk
N7kfNgx/1vyIIeVkU0Y9dHCSxhWQfp+9T2OLBflPXORKBFoT1W+AU8YQ0p7QicDu+qZLUisRSzM9
+Sba9cMad4iJh1EdcH8d+EDEqWR61v2mb4Ohs+7ZdJrrmc8YsCzWvTN/8DQ2+qO+2k7qjClKlo86
j+ZhCOCmE8Aczo17nYLdMsX4b0ZRFncZtcglsHz0lc1NdBz5OYLBPkfupL6qpKJGrGr+3Hq1y9Cg
lGyBfeqN7Gwjp2MZ1wxpcP0N3FNz/dpawAcyBW+8DRinACE0E0NgHSw7hoFL8w248XJZTV7sB3au
v+cx4xQGeeF9RUola0BXyaNgx2CVl6KnB4iAYrIx7zDTVmb+iFKykf8dOyju5u2421uF/YFzBIcF
/q0lMZ1M1HbQQn0r4OeGw3WLggABkAXfGS/olNvESz8X6FHw0rSV/sMaKnKmXhiK9gpMMeVAZVPJ
zjvqmS4u0JfyO7JncYAzF0N45daLJCqKTAz1KqweOgF7oH7tU2jG1Rb1/PNAIwp08/vABQuNI5DG
pAMSvDC8qOqIxA0jnfEScJpCLfyRbGQMMxbnp9f7M/59YqVjJvR6xO98nVBn7TQURKYAvdR8lwL0
ewpkPBi/8gdVSscDTx5x9sT5aZrPshj5kSElAkAX8ySh8iamuKZZ+hLmyll76nYOWkJ8HbEaZUTT
WlDp2/gCIMTnTUYoasmMBB4xm3QtayWadd2tBW96DmUxSDMmOtWm4kmRilZ/dYRVuojQBWq7QubY
e9pZNy/YUbzY9eJZt5PDPX30v9VEuHG24IGy+lBSupCm2APW4D2kNq19AYN1CWgMOFdY7SEbEaAE
Td+HzKEx1eTuWhQ6cdHOQbX7w1Pg7wXr0IIwMTG5TX2vyWp//QIHhbB1eh84OhmZVM6FvH4KTlvn
78rsQH1mDaZQoykXitssr14rGi9CiCoL77DoIMwIeGCwO5XDtPgsYo8OwVLtnpEidPcyORGyjshb
qzk+EiL7wVs6Pz/FAeWgkzsLwtiikRz+SrgellsgnphCCeBjojLWfP6yOvXYQ6un1OW4eHrxgBta
5c8WpbHQFFmCmqRXoc4lCWlN+N+jbguTsVjR1FlJTtLZZiHzYAe9SQZzWntHLwLSRRonxcAQQUww
jZdGtqZfOXCQs4sW5exStNUYVERsZjeRUO4ujXc9Vks5lXkmq47AbenUIDYLGVhRz38d7+c++j+I
nUolLWoeoZu/8JWtWVmeqgCDDIEnRui+FnxN8BrLZ27ra2+bV7T0aIFKm/lebVTaXzy4Ieeh64Ic
xBTeBLZ4h4MbQpNbBjoZZx8+O4gnWqQErpNjMRbtwX0NUuViPRPNctzV+dmC9ej1cEunoVME2hJz
XvpEhcCFAepThhhaZiUHUYldDsWFGkpbzFthV/iFfnByFbgsFYaJCNzHOgMzweIsZgS5hoGBWWhG
JbOQBY2y0lvJZjybup0IbRyRKC5feBStAxrD+qJ6eL6zOk/616Fm5FFV3rm/dJpa0Oy+v9qhC7pz
JLA9qg/1UWNSamBXFDYuK1Si16kThWrLK1HdC6al3EZq7ibRq2Mp4o+PSo5pag8AwWK3uF7vyCzj
wfogObFA+C+buCdqfj7FYKwXuWAZ2NFbtJa88EQ82ACpeH2F46IcoaFWJpIjXxMP/+pSpNXJGTzQ
+uCBmpXD02/2OIWfK0nNW5HL1U4Bu0ghDXxNU41uGkYJDOYBMrshOAUBsEFeNGYD9ZZk7UG//kHx
sUEJimD3fTZf1j3sy/D8zT8MuNZWBXSv2E9NB/fgwavhZnb8NMbuv//biAP1ZJcNk6jXTHjf2ymg
nJMHnc5JxPaBVG2bU22BYUkMh4gF0ZGfOXVyb9VrAKg89nsc9r+elSy+CtNmbhQCyuC+1p2Hd7Y+
aZ4asPeEPMEvQFzYrdQ0mZlVhggePjIm+y+H2MPBshFY10u2yg6XtyITtMexqSAF578h4yYVw8SC
hN+RZx/9rn6CLJWJpzEKxPhFkKN4/bVIjVsNBxfwSaqVQs0y77wMIPRDCx5kwH7CZZH+QQ74PkVR
8NkAEe0UnCxX7I58zvpeY91nT9VtDIuY7+FcmlgOLzrVG7aP5l23vPWq995ZvYN3Nbla4IPtxhVl
MvhZQfIBHq7hwHZw23c7H92HQDXjqSze4pT8XCrjW4y3SI1FExCdAObpyE9CJXDnFMwoGULvyv8x
OWLO5CK68B54S8wQtWZIPI7gQw+/3BJ5YJ5YRb5cPp5iXY7r3fDK2okEt/ivsNH6PKfMpQV11bN+
kn2IuddZMIYzN7ijdVt1gCC86XM6T8j46OsfWTn+jvRn5/wRxHtLCbDZiIzFwFIuTa2No19VOxQd
AbswHYTQXs7c19sYEVmUPGH01Z3DzNKvK680nt5tdCnE8ZNyOc4H5wFkTz6j1oqHlb45tAMcrLWT
jPvWbpRpMf04f5NyKzt//c+E//b8D/Ac4I03n3OiMGWfF9qwpNtjtxy3NJ+vzYeBRAQNxwDignVt
kmHftf06wW+WnVWcIb6oINc94ObGion7wwNHgxmc7wucow+vEGTA1wlhFJfUQsXg6mwWsmvLhzau
HrxcbGJyky/4aV5usPRosdrEdkPP5auehWCtZYSOg60syQfz+dZhtVTZHPlb0c9Y2Mp71P9X7vj9
rvOfeFnR4X0u8fuqYxKrmTGQL4C/Of89WNQjSP35kpAmQzRxy+JGGqQaNwxES8Mx0dcq+lidgAOL
yXGtWE+IV7FaFSAVNIIJtlfnrm6f9C1zkK6BER3a7yWHF7D9ej0SiH7oK22VDMRRGx+IrDyCmUDz
AoJGsRlXd9lcOEIxV3SZaSPMq9o/pofEP13y8WD4aEE66EeBQ2sxJN7w9qA2PlztxJ+neQlAZZ80
FaLiKFc0VpFv0W3Sd1la+7UvCk/HOlSLy8HUtqBslmY1dhvmqhjkPFkZycYSN/+8NYDyFk49TWND
Wq9Ig6MgVMEwzRJnLaURAR5I3fpS49VYn5IcqN9PFKx0nXyu3US9q6ya6Rvmy8CJHb4WAhhFX7Av
cWBA/eRlboE2XLoj+N7DquFvYmLGnSHLOSuTQnInArXjliVaR5LBFoFdov2ybtu/5BKfZYqxsH4e
Zu5+CFfZyPIh/fXNqABSSxSCNVFDYdgPs56SmwyULPGRTsxuXcnxjr3fK6yBsMd5EtYYqJ+s3fJG
Bakt/59hVy/IBAHn3fk71IxZKKM8CGKtYNKkIsG7OFV1a9HXMM7R2Fhn3XE4RhMuRZ2uWSM7Ld7K
4gYHdOB881Y0V0vbePrk5m3UCT55dlC4EYUHmC901bYKd2iYlADZxUN9Pwd+vL6A/hmyqCInbVbd
6qi3aG+CxJazWdCuubb/F+Wwi+DR9CfFgHfHNjMXfzJTf5Cnde38pRKmHaCnMld8bLKmtlFmAYmO
G8NOiCZZw1upmfvLpDSHediiuJ71ZuzZFNh3sbfEjWrruP2FNRANJYhHCOMI/UCWA32UkMvmTNcX
nP2mQsVJrwly880bnIBLdS7eDwi0vhF6sI9WJ/bAQOSm3gZTE2QHAu9E9mJgmbKBmAtk51e1WzHc
zwRM21CMiY5u2zSxt24nQy3CUd9xOVpw2/je3Q0FF3Gag7FdBEDzrmN5GmIBJQw3L2X36SkyvKHM
Wnc61TLmtajR0Non9cD0dWYpDUfblSlOTV3NEO19WLFuL7U4tlIuKN94NHmk6BhlrCvsy4EGZVla
15bx8hi666SPqlqfjto50rT1LEYgJCFcyQzdSGHfGxbHuBSgVeL1LbtD/DMsjIRYBwsWoIDPu7GU
L0L4wD11AN3RunrVrBU+3+Bz46nUmX4zVWFHKhMKxExLAXH217L0O+0cD3ZwkyfwmK1IQO6g8mM2
pwf3Jm3Ly5KQwQ0ef3MQSNfUCionBvYNf5IwR72cdXehC7XD1KrAaPSKH3Qw/qXAve7aJ0amEwFU
q63J2kebLj+8hhXLzkmB9Ks/cIEbAiUK62aALItMGL9HRhv1PVExcJTDRlMbhYsr5ht//wcjuqFf
8fWeK6dorTnYv8JT7oQRNLdk5qEqd7vBVbJ+uZOYi9G3OF44IQMeTblxxgeAK0o6MjqofMEKELp9
u7Z5n3GIbbjkgIveCSOgvaN0fMSrZnfGUr5sFoky4WyxNiBtrtE4ezJp5S2LL7HddeWU2C0bDY3i
a4abaCqMWMptqPRYlMBOyxEgr40TLpPKUO9Wwa+pK8s1NEzkyKnYqk+gx5gYzS6X3BqmnLoD4KgQ
9En19VsL18ZcVGsUobWTDS6tGMXH6Aj4T0tBlyEq3M+s1qlAwCVmtPplEKOYPSTnLv9oTOHBmvx8
BN9tyuSmd4FP41qizdm46Mk1AujGrp7Bf2u4Xo6Qj1SftL3P9iroVC45MAJg6nFdLU2/0y/MXviT
lOfWPtBf8jphRVNEExiNZKgLYKwvfG7UKbfBxvu3ki3wiqSWzaBbpZQMmnJcrxWj/XaTaM6W8Kt4
D3R9v1gJph5gJcQ+w9f06/OdwMUFk6t9mFF8SG+p5pW4Qx8oDU4drAAF/K8OP7+dEhw5zf0HKTJl
WbFq8zBq607O5hOFdUJtlzy3a6Z6kBANglRpXdO/5OMVWELsdFUz0R2wOx/jejOYVkmHbKV+qG1+
a+AacjSGnGXrrHDlumwPT+ZpJLgAbZOVFVF2g8lVU6RTb5UDJSdpZ1cjhWzpLYfylYFXhgLRtrww
VDOl2EIafZ8Noz4UEAfFAgL33BaNXvDUONeq+9pI5ORkd13yCm17fzg2YbsJliatl5/L2/tKmYvk
Q1Wv5YMfiGSf6lTBfkfu9BviLS0o6ncaf7eAkz8FTRm/8jC01rgpxJgWoKCKUIMqmekbDDxFeycU
EjGEX4eDPcbbEdJY9MiUA8LJISz2W1lUubOCPxit6mtyORbMBPgpkZXwU7a7i2EwcCzHRTSu/3k8
q1w8dpxZ4GjNDJlBAisK2DDe4PV/ycs1AzhwkTlAYQl+SC/1qdAubO/SGcw4+ctEk3wXNLXLBXQB
tfTR0/zghRH+P3fv57hDmXFB+8+hyTIcoZmfalk2ruPVQ/BBn5l7NrRZmbTQteeGXsHKDloB4r1B
ycTWhLgmUpwQJ63dSuUgXnCTVS5CVxQ4h2WQKw9D5wIDeDYVWc0XzqDpkyv4swbypULSN6NGOvfZ
UPQub8+EqDfFzOdcsTvIlnYs6sgRW9NGXA345Jva5zQOpc7wiMtbpwgJNVrvGSDGBGgpa+4QOLjW
nvgJH8CDmBUgOwicKfyWwuKiGgsCvo463hBi0MlKmJ7MESjozUM3vNyHPnoKViygXiywVIobSwIB
sTZMnCrsVo47EfIIDQFS+6EV/NivhXx5zbeO1JSgvTwmYiC5p7ItW2yLzeDBi2qEXH7V2P5DaZ5J
RrY1WkNLam7i09XPp94nucBMsb/nTeGTLAAbLz1MC3+7cP1NDZvuM2KIUGS00O2iPVfOUQtKYUtr
Ecsz8/RP9v+xyTfLtM0KiKLasGrOlt67XLFhF3xxyHB04J7OTJqi5tveU2Ny/7ObcKt6BTDpwZJs
ribpZC46+ksXU5mxmv8CyMzrYbC9lf1usCeXQbWjmKlIKkhwozx1CdLJHeQ6k10prA8GE9aA/Is8
B52VxzW3S/av+GiF/a7eS7CJ5JhaVc1qBk0tVBAZP3ERHgn1PXbHvynP+jAjT+zJBKnmxYtjXmhP
DezUmNhARN6x2wFeP40A7p32LgrvBWNdVHcgju/OPjV3gES+EDGgWlWC9K3UeqGLZTCgF4zq4sc/
Pgx3PCsT+LVK4yQ8LuHMueyqJ3GyuoY2IP8P/PuPBHgyxqBrTpTfjcg5mT8HzcinZSv5Y1N/5laD
FyAJ3jyiEnsr5XwDP4jLkAXEA3PBHQabyNNNcjT/6ia6eCUj7Zo7xLfuJRd73FBcJO38U1gn0Ofo
NO+qXYsW1jWGuso1EsiSgCWDJDlUgeL/9VbDA0mcUwOwXYS+uZUg7DPHtaRxNDXUPloGML3mbvbn
ERkjrOAXbdaxflZhN1/E+OMAHwb0TiZ7D9YSJrRfwCaVMmvmvsu6gLzOa/JIkUNNag+2DeaXgBkQ
YXMqgjJ2gqYNGtohSJwrx8mJwhT8gOBnhOzY7CIlEShCnoNB0qfvGZdGXb/wt7sddJS8GwMgz06B
Ebm3FGNCSJkVdxeDa9GzwkWoMslFzmoQ/uBTxMT9s+bep6cwM+a4xgypxH9Ww7W5Bnc0Vn+/MlIK
VOAsl8Kl/l3IDr510NwKXD2AJwqZLOmSDQrDcOiVzkDMCKeGXbz7JUpD/uZi/CEZAMW+N1HqokPC
K8yFYjSqcMa0bTjnAYaP/0jXZA+NxUAWLJJ7gHk7nXFuXsHS7rDHEOVQfkVVcih/AxjzKvsiVZkD
s6js91QRcF0GGEYrLO2vOJQRa7Es+rPA7A20HI3iIVCD0Cb6BWueFjmOhN8xnLs7ILFTBVRfskj4
F0DXGneWTonTPd1t/ilyIlHbbi6Lp/g/O6cK1iNBao1lSSugUBvq2dczM1AF5m7HcAhjQ4RgB+mA
+msD6fA78ph2OG3PIvZYsp2qGwRJIHlWAm5+QSs7HgUuLRo2cZxR0Dx+rUjMcNrudEhSWmnF0ap0
iVZJED03kErPNqKUL2HVPzQzOp1NulvqicC0hU0g8PjAO6kikfv3DkyyV4FN/WDhBlZCFn664oBw
1PAMreecJ0bBLJ7MB/FMIpdPszp/A3j6jZbxJ2IUAmHrVR4N9XDAqWs/d64JEhML0xILzkbUd1Zc
+eMuQ8JSssxic8N1sRs2pEXwtZNmBvDkol3OvtTecCCGHHmbjE0CM7C25+M/QaxcbkxQJVERrrfv
n6y4dUGfF7D2aNSFh9iAn175XWTNNJKG+rDphagY2BC54RSPHNrHqkIoLUP7KKcSjeEz4tR1PGcI
qoRkJPc/iD2K1MkNiHl+nOZJ9CU46xYyYHoX6MUrpvQOjNHTyDQIEfXR5grpo5N7y7ayjLKz8aM9
6ssjumjFF744tgenoH+cFGo/41gCrhF5MkabTiDPjDTvS5s7Hjoq+eouGtR4hnjZ9zzJ27+j4ZUk
U6EGHong3LPQ/sr33zkQlaeMs6wy9uXxbwSrpZM/uOW13FdkEsnKp7j+nli6q7QD4cI90/5eD+Cf
eojLaUrXZY2O4ZsdBsykMumEv7+wdndpzDVrWWM4rN/B0W3D53iLbopLA/xTQt5+hl2i3K1bbtY2
uKTGA0Y/v4wLc19yBgh3wJFrdbgVZaIosGKFfkMF9dLHBZEB6aVPlsFzAAhOvfJAl1vLoeEcrd0w
iOL+/vBz63z4VzgCkB+bIXfTQTpP48sBRQwR+GBmB4W6KlP3vQgG+JlxMc7cHzvsvWnGbqjJiXYX
v5mOXbMxpHbNaeegqeIoJCKs0xGFetVQmP3miO9LPQRWVbBwksIK8T2sju6BpC0rPMq+I92oXleo
HAXDBoGONC/IBi+z6tY1MU5T/P5BtBj6+lYH8Xv9e0g8+zcRQ0Trp17TvW7dQmAl/IhuF6E8+5K4
GLz9yib3WY5YfFX5n+imc6AKpNJaAYiPY2KeT0/SW/n8Iu8NYSRG52fYF4jkA3/xjMtPYSjo0uhp
07vD6CHF+rxUb4UlH7pwIw5zRTiBTxCoGRkpQrdsDZDBLWmzNCB/JO6yDKx6oXeIXaCs2qTUn5d+
BXMm2X5Eg1aa/J/iHACuVLo9e/8RyxZKsiSkn1z0tlLeys4wtGxOfK72Pk9/tTAJLHU+2SUslNh8
JSd0kioxFL2Qxf3YKxRF5AinjgwW4Ya3ILL4LjNt45ezpvxDW4JPKNcSbvNbEm1HZErQC+BWvEaF
WgoDSVD8asHdYWjfQdi34R51/BgmbrT4djwE9mbMr61PuyARN//0E7B3ccHob0ohVLNcbEo+ZksJ
t8FNbVnV2gBh03mIHxHA44rPaXlPrNK6cRIJUGhB2VZKp/obXC12tF+1K8w6EHGPio33ByANNlDx
ALGObg5LeLq5SoS2x4dBkkzqsEeLt8M5aLhzQzaMA/VUufjEuBBIKLKH3dIJNeDSykfilPlzw8Ey
ULZjCzpzhHwaibtN79Rrwj0S14B3veMHMbdctm+u7nuCJ+DCJbb6QeSZPUSQfRTwtpTk0KDRF42p
D29buUUN0K41BBYi3VdG/JlhkqaOFUpfnhsZsmz3H+j5IuqxZhq7dfMLnGN3rFRierLIkO9f5y0O
k/crdgVRss9a+vt46EZ39ebGnCX9KL2z7rwICO62a0fvPgHpBN6YThtBZ/vBzhD4e+1IEjCSRlhy
9BOZ8TN8bcUGyxbD+Kh0x/IRmy6F2RHfXtfuU96BxbstbkiuFeCMExBc0yetOnObAShWqY9Io4C9
p6MCwe/zvFEfFOneqcgOFRAkPQFHNE8eMsb9YFXj15Q+05b1b64jItWWiItulhsHDuz+pHJCj0Tt
IaG8A79Y0v01ZBqcUmAwZPScsuYY45dHZZ5YA9xkHksdFuFSIKdOP3/eY5lel7XRlxoOkaK0+IeZ
wmCu9AUg4XonBn4A67zNogm85hhcJCko27TTUqQ8CCNQVZRnOGxYlDCUiJp0rlR3MYG0fGd4NErI
ghmq6LlGo+cSiQyq4W2E6/8VnWqcdcwCq2HCbqEbKaKQGgOndt9eP3gSnnkHw3+vgBiNAr8KuWbq
jsi6aXD1DRbXgLQ0t1bf+z5CS7vUAI4fR4K6QR81qzdyMptJtSeD6xBpV8RoeAZ7aLjl3C+W3uPt
jR3Zwv9F6smnUi7HUDWsAoQWpzpSKS0xDeUoyO2GlHU4HIjvtjJEEedWlMPhGID1n8yJ1NRyUbq4
pVXjk3z7K/Tb/pryllBCrTmPl9J2E96//yKmqelNMj6Z3DSxXNSQ1NLbqj4s5Lcv2bHgwg0oi5M8
EfMWGLQZICbknMsFBklFDi5PrxV2eY/9e3+qXC22AXjd68JpyMxOH7Bcq+z8YtCWuuFD0uehstQp
30sgYTz3GgCOdCKj2cuqJ/qCTXeaJdnOn32FUorUfw5lDiG0FsyiMLkFqgcOuAunMk+S5z/c5rid
MzNc9fm7CYznUpp3nhKLB7WciR0Kf1RoWKQqVgXQ5W51t/frkgZ6Gi78htkSl7ikCX0HAQXMLYos
UzZI7w8B5HipruoURmc8z2OGQa175urleenCRK8kRyGbbdlvKmUYtvAPC3Y+Opl3/VrmJDvaZlsu
OrA4Kb9c11JR4LzQ1cXv89Xaa6TUUYkpo/muMFjhCPIUfGMI85ihG9KAMIdSuRn+2UmD00gFz6mz
qyjAMyzy/tPGFpP55SEKPd5RX0hbRxGk5Jy3W8G1rhyO+Q3yMmNV9/H7fuh54VNbi1uKXS+UmAT9
+H5zKOYmmjPWGeX8J02NWpPOAm/MtPRO7ZNJQsLtt1/aU6/DUUlfQtkdgt6yGQErbgTHrOzOtZ2D
IKytbB+WOENP0BOK9TM+sw0GZ+IttfE8NCY8EZcw4QTh8AiYiwfr3indCCKfl8Jr3RFmsTnfTpdk
9uUN0GPyFnctTkZn33uaUZ2/SGD4Cm3Px/7QEbrav7GEN9DWsewkUcgn4WWGcDtHITQjL6DvS3iJ
2fW/uC8s5BxUmk+GfDq5VBgdRhiNCo4IaUbP8NMOjoV+bfMOkDnVwzmZNOaxB78JNQwiQBgikVmR
ENSpLYL+Rak8nFkS5tXnckjKSmGGjCMEpQED9Ir/yaSki6vk5idAvdWTs+6tGjkWJHYBEMwOqMw+
wRNSWm+1kmisTijBufCnWZ4nBHq7smBljKN2SxFSRzxY62Tl7pVEbcdqkYqHdaCvxJZkIYo+F54z
M4mjyFbOdKE8k/GSaiPdw4qIIEcHTknWBEbr6WTLe7roUbkyRxaJqrR3wYl1BKgdeIjV3qvHNbto
eJPqrHaQvtqIrOpKPRwy//jsweAAvVlyQAuXOsfEFMbey+oHVHjG12447FmodvOAAJMsLV+yBHJq
7ijZXYiSDSXkiLMpOjaZfTTWNVgBxwVEeatLp4s0CmaWBQZjO4s++wI2GcyC/D7vLHqP/3/3r0nJ
ttGwp73OJlbNnQTxCKjnl/gIQclLgYJCdeWXcoFfCDEO+ASMhPfYzg/qYi0dz+o/HmGFfmKNgME6
R3WEqukQOo3PN1fvTuKllm/BKAC5lbFJXFpSLqtOPB4PuR5ROfKGNpecTXqFJ5r631AO0cfjHt2M
SPbIg+0MRTimqaZufzWJTDORAX3NSbrLgHO7SVwynE2U7dQS0V3hvuCyWa441SYZaGLYCksB8hal
FaQnJf1qGSKWwcsvuTE918kP7V0J6VMKF05h2EUnsgUGORYB5hZM+YWQ4tApoEUt4JIx/OhqDgCF
j+UhoIfa0v6uzR2TsaCEMPIKdqlwIJpX12YVEoVt45iI1uWUY4EIpCO8qgc0TXdvOxInG13zUEFb
lYQ5oIK76iTOE90pMY0ojn/jNee+5Zl04yKcEFgNaO7VnrITIP1K7nz3VFs7tREkc6KBG3t0mGuk
MUiy7+EGQSUhTkQ6cPVXZmyKrIkc+uyp9dNsAJuVbrbqu5oRuThk7Tw+/yK2BLUXA/Of+amsP7Vl
AqaqwJWQuiLz3R+WRfQlR/lZx6bvP7KnOJRWu1uZJ405l+Vs0NGbt8AIC704y55Al3AhpYD1OeCn
fyAKWUkYbGal1o5RQz1i8t43KH0D6KhsNBKl6535J13sl7oPYDlW+e6ZMZsq8W6xWW/1ik+0WpMe
wBPN/bAes/SnW/BwYJr6IqAY+drtdeJG1fTB1LH4N/fBn/oAWfvyAM1BdGmH/WDb6SC4SjX+Xh3x
ZVtiqh6kHrN/dA0Z12tMDo6wZi+X2oWtUTWYzeFrkofoSruPBtZ0vLuG8DEBVLV7L8BJx1Wk6n1M
rQbjTK50L4SH9aUNSzd5TMojxy7P4L4Wsshp5IvG+1yyF3ec131Ke5wNi2kYqZ5cRR0jabg4MQNa
m/qM7pFk8LrP4+ycgti3sy2eA+rt+n5HrcvcFjdw6rpUWBq9LmaIcfP49mdJZ47GUeKjTKf04apL
LHfX3zYCom6FHOKHstJjnxSRwJQQWWyw7Y+akQXEeCqy7IPw5s28kQrC4JnCq6sAFXpNeSHNO4Oc
jPHSLOJyliLH7ZUbswIY8KDt4bzQRzTlWyBALjdNfDm/yoPOAijoB7PzrZN+dRmMxykoPfn4H1F4
Iybdhoidx8WAsdKXhIET1iioYjace9+YY5yOrtqbojWsNAtOCD7i5X1GpAXFWmNjCDUGblpTYL05
utuHc+YvmnGL/Z5gzLk6ktJUW1CHKXi82L3P07ylIOMR5zjPCsrILGIb4Sw3Z5aiEk2YlICKzIFr
FnjnB8xuKSDOkcVkn7WO9iU8RAlNkxXscdzVyMNLSOhCyA3G/MPlvxhWDwUrmG6M+Ya1EOQBHd+T
LCfgpmIP/UsgGWE3B/C7g/3L9vh78pXG9WU+yyos8uwP1b6O2oDpm+Snn1nsk2C1fbdCiDYeOmmM
5CPvk6Qi8fuwpffaPnq/UoY41TcrrZO7A0SeCE3fjpQ/h0eS6VB4icoYk/7x2WpEwyeyEeWSu749
nD8/TPZxmIBLnviEgB7pTfdAQFygnxmwY9vJDdPhaSkNoHmUKFkmInKGuy/yGllAGN1lvFuzq6e8
JyZ7ATdgQQ95ElIGbvB37g4mIjI5+VpBUD8GYZnyIwCrFfOFrZB/uvECkDzJbnfcsEPpeVPV29xm
PUZE8r12ja5OSqxEIo8L1sj9kp2g4eHDhgC0WRv5kD/La2WFzLjG0YXHDUTenJciDQfvUlvbzv+g
4bmTryVrknN8iMQnkNh0BAPOmSb6ncspfljEdoWSWpSGW2QKHSeBPPxQgIYKHaahlh5KujK6UCns
irTVXSBLbruRDOv+G3jd/gy25NUwoLi0REeY8IpY3VwCur3fQCqv07Ns8PYRMQZmdXVM5w/stjnK
uwK72TZ1ns5GHNWDL4AY08oyRAl1uJZxi4pv7DuBnseru/paiOpyBy0jejnMlvFSKm+9l8fbQmSb
MRyClaC0KobjVb2dIIHIdkyEvJq1875sl9lfwhSeNzaOZPhaxwNj0Jw6kBdlEZJFycCeRIeTVi8D
hZytevzJxSshVUc+GfilAc4YwUD6DPG154Ok6321bBNiy+/CUcl36EtifpCJh53mdgpZ3iRJzzDf
sz8aAMO6cuKQMLEWgu1EgvagUEszirShV6TlXZe+x6/3tY9HG69Ux3F1NUYP22hdgmtK0mF+GlDe
u70St1jLYwVfsYmhmBwTDzUJp9teoPE883hkRNb654TA7biXgMnx2wVVQnMEqLELGDMjsVkevrRY
Lfwp/gUoV1ImTyN0kVfjOATY4HeBkrV+jK22/3Qwomxtjo7C11QDK1Q6yD6/nxy2mJ8WH3K/qo91
z0DFi5FhksDiQIMFSbWcR2V3u8QpLqSTzEUGmjj0r+azdzBIAM2v/OMPeDuZiRiMoMlFsBCHjsdm
NQko4D/7ZbKdLIitBffTN54tO4z1vBRP/KghBnmJXUgoNbO5io+4/yx0mozG5WRXQnIwzJ/MWy4a
cSpL2g1PJ1fkWPmqmKT7BkHaBHpJESDtbbKOrh00FKBNgiFqnBq76NguDrFgBtYUODNc9Qo/lb3I
+b+6xKJ1P6x49C9ENZk8y21tv5BP0Ivfh7ySbfKnnCjWoi1W+2P3DOAQrErOmy4PLH3N6ovIZpyf
7BiCnh1Bhos1+MXbSgYC/pbz4QCI4gZemVb2X7WzSG9j0BNvLZAdGPEcnkL8tYAoDriGrkbiCB1z
6GE3ndfdUdEPA81vWRmhAKA+oTUNiekNS1xfKVKtC7mUXUPbh2hKnAfMpgJYSSTJme7BPbrjpX/m
wu++Zl2Av+dqntVxQr6adWedAuG6FszecmRlt2+QTK7prEuit55JkprFaJOO8s2JPfZzb+u0dtoW
hS7JSeK+y2jP7b3+FkbBK2bw7b/DqmNCpsplFkgN0Zg4UvRrX/A59pK7nTlWM3c7PkdxZPYybXdK
pF6QLGZv7P/SkYvM2AX3A+Nk/TtOHFFaFiu6Pvja+Ph/+8y4h94RDsBosYtcmzk+Erx3/XFka6Ft
Pc7BSv92t/anRJR4Igq9nO4TRsbjcXYIEwZ8FpME5791NcmGu5oxOraLDhOQ9i/pgEeyodOR60Rg
/T13sGZ1nxe68S0jhBsCyRJqUlifgJlOslYWImQjrJ0sCSuLlresw35FvSay7zMSESPwpgb9+fzV
ypIS2EsiJZai8YtiLsIJAVucr/xrZqU8He0DJcYSEv2IvdmesGxWXW+XfbenRAlM8w/q8/UR/AnG
2RYMyAhP5/00oAxAMCuvU4eFdkMn8BtoAwoXE3V6LkEhfjMZrzoUm1WZhHzaYDVpqbjNLSrikClW
M+lI2tViSPGBARF9PeZs0gC5NXmBWRjToqp/baexATV44iZ0NRMRG2ulWBgx8WeYSWDat6diEw3r
jwQ86Dt2pAiozub8UjhwlNemSJTE/K58iBq3nE/HEyQM46EwcbEr4vNYWV/m0/0Yq52CT9RGvcup
lSPasdHt9fFCaQMg2PmK+yTZ22+XrbTnXN0reWyIW8WYVakJA93VXnmqp+3JBXZGe95dMU38NPdn
P8p2eyGUlHVZNLavXniXScXiqvu4R8La/dY+9kNkGmsVrJ1p86TzwGjh0sXaI5/xT2npa30WLZMF
6W+m3Tsff4Q3fpkxhF/mE1cPh5eBPcemuhTzEweflalvBhW3qNJn88eNCkJYl3oFUamEiYt11R8J
Igl2ap/TbVBB2oH3qqP14XcPsogmZ16wiL5jvBk3gdWPjtj3uWLs/LQJq25VATzsQ4fhjp+E8Z35
255v3CjAIkEcsrs9NNZxFS/6UVqXoK6+4qm9v81V3WmTnqO1Jn3mbv+tO3wFD4N7auqfweJZLiqP
/LWP0gSqXtglakp/Vjq9NUBGcnj0d9q58oi622WvZhJJHcIKG5MrEtnCE/PWVShzSeSeJG8Ka6IU
di4hXnz6TkvOhJfQCPpBj7ZijHdkOXMfSvyJZ1U2F9+PU8IRxqZX2EbomzL9UebNYH87DD3HAj/M
raOv53rCCNBi21v6rtSjk0S4+P2xIgWOPxV6F4tUo/Lr7AJ+hmNxXD+8MDj4npgwNIfztAozPc5s
Kj7DTwkOk+LNEyYFuy6GFag/nZGc02+j8//RlJ511nBIy3qffRMuJ4ZX/VGeGmgY3h6V5oh1vzF3
gesr7eKleYKbAoKpKK7czIQc40k6fQ+yt+YB7qxKMC7GadobqzgDq3z9EUg4Qms1IWbCNyMCzYkZ
PkJDLO35fqufpz1TgK+wRwf1gt0c4ispYg50T6Up8h2cZlBgZLI2x74TfoJbAdnQdcTQ9o95ipNf
X+ycsjUesnogrJBj12Y+SHtulCF/RXbFle70EgGX4SI53SJo6dwuN90Tx3gb7/gnYEg4+yCv5lhA
szWGzcqlAPWL8wzwJHRBbusXun28HpUSD02vqwRUD1H3TcHbu4PskfuVgTB2nYjrqOzqFcBiciir
b5owvkUZSYkWgYHFLQeyMxBA0KT5foGQGG39zYs4JuwRa9o2j3WVoTHTJi0r0ty/6eGRzoabzXoL
M17b8IvaSX0UwgZbQBL+q/9nwqoFEQ8LMmFIKYreSKacKef7SZtvz4a6zUDflYFWvjua1uSK2foA
oW0De3WRh/37vS78+vsDpEcw267jnUr/JNjgJ0f8au6WeZpa5h6/los3TlqGzRdZq9ZJuKd67Plb
LXKYpwxcJAkSfngm4z90mTIt0pWoLvClB2vnBK3gsxdeGyHmnI9kLselwmIUnXqfXGh+UCNFpNaS
kUHlwRLcGn2ngOqdSDW/py2uGfDX5GAsuRIYZHCb+0wg1sbA2/jHAvS//MUc/iU4W1K7S/wwpIoG
HtMGLP7FIJp6sVy7P/zUqegIUHtpL0CjuUZ261vqvtM8fg9CMFqeVlVuNed2avEYjJ2vTM79g9Mp
eWf01Iu+rLq3EB78RaBAvaFxC2J5R0NErHsVYc6D9qtaoEfYLJjFM4MWlM9xo+4sMBmo3zqBJvM/
kIbosn5+bMxhhOrEeSsmNVuzMs7mpk//fA1GaY2bKzrJJXxpR6kxfrp6CiM+vXpPjw2DbLaWxWaA
SspSx6Zzq7pudyo4ijWpXFPuB+fi+fwIoIUVU4doCryoGHTiyIIdmQy/QmEdAnliasNgpj4jxiSm
v5ELzYu2wlMpxmXSgNsoDwtQBR5Se5Gl6ohS5mi4NjO3iv9a+TLyGZ9XQJLxLGxeW5YSn0rC1beY
FCoIabUpmGba2dRdZKZADVA9bqau8hzgsudRjvAse4G3GMvjdHlXvi7jD0Fvhc4VUZJiLSiYmj/l
AthjWv/yp9QhBXgbim/JY7PDL+Whpsj3kfyJpzXXasoRjk5XDRXxA20ql6vc4m8nj+DgJOYPLDRZ
BGCi/Jm3DJuJUBxJl1yPtFDdzDKiPJgtsegCDNhHtv1pnYuD025zxlKHs094l7/3lcuHFTEikRXg
9SUbXwJWleSRWYrU2kvbHSIF91JJCYegnjBrbcTszYWZGundifR6h/KeZoOAQSFVL7LHh+csk6Ky
AE3FtjkOLh8GoGtJv58MsmIlYcYLKDF35f7eT9X3YBMOMa/urheHM9Gbggkse2tgPwzBnU4iOzqO
JcsFc9eRVRQ4JK5pSHWXZgFNKYhXjNRubB8hXbpw5D5cBlmM/ItjCWmnj8lkFIgGdFkxweaREsTk
5PobeBw/OdUCA3MICN2QKcju3Sh1DE6j4LsvjIJSaqBkV/NgUkQJQzyB6n2JDLqN/8wuCyRyf3wS
0iVmFSh6E5/L86xunJ1sz9AjHBhhnQBrLjH1RbV7WUe/298oxWF7xTyykXmu93A0ovNDeTqTwNDH
fOssIttkU7w1GUwB8VA7T5EmENd+idwt+MrK5wE8qTAzd5ksFewO3jcZ61PJLbspn/O/OKkYNA/s
6Crc75k2/z9HzJNvh7yi+5QvzH53NvaayPmTwYyqg7xKoAuxANcbreUI3As2T0NKX7Bgy0HNjjKR
8pxBtz7ws0Zxq1RgJNUFI7PJWT5U7ppV34hzpkW1L+9flMiSediEjlbIwWOAI1uCCawfruRvXZZ/
73zrAgzeFOFJ+r1vWoCQGFbhMdQVp45AhYpDif4TSCJVEm2v4P+nFG3u2Wm5Vu3xUBj2D1jmKsHb
aHf1iSJtPweA8QBM6MWCflVoFa6iOHTQLfonNgEMqr1ncXUr/zwP4QmhXGUuwSBUYiyxIZhEtGcC
uEPZdJVT+pRNUWuv8Bq7VmFWH/B4l/DqZkRMcGqUhHKJrdhHueI23TnOS0ONE7b1kOlwUJ4GpFXy
NTGa73kaZVuU7frFOqRPYkNoqSSFRF1u56DlPYmVSumNPCpPvfIfMJV56L35im381okh2tksF8VT
IgPLGA9YxRXaCnmRtiZZ/gRMfny19ZNAVbLiAhEiS0D354K3+cl03DTJB05XioY4pMU37hNH2rXX
8XfNHrRtktXVbVDkDdY4gZ2AT3+//r8mLs8fDKckiOvb9Zz8g75//BvnZkoFzxOqoZsy2RoFhT4r
qjQoq/+AUnf/ps0CHG7T7JyE0lg3gb2sb4wWrwv7VP4V1fVafdiKcUQocAXC/qrns7yvxYLS9Qx6
IVvWiEtwGMFIiR4pwRi7pNQdYBKlqt1V6B5fXN1VHB+HHOqby+agUAvE01Yk1iGnqpySG7gUTm0p
MFdlRxsTT7Hly2BnMWxqTy7ORLQxfFP8ZAMu6hM34lG17xZclRqDuX4pR/cXiH7GKWV+k4+2Ijur
hmvlukqwlmTkZBKXrn+KoUWS8W1ZJaxbhiJmfxJEGVgn/LMh08DB4D9ijvySRjVa+Yz7RsMWL6ig
7zu3jjNFrrsYPIPW3iA9kzp9TiCxjCz1Tsqor+6qOlM+PmSsxEERlXbmKABPJDdi7Ei7KT+SeR5f
GPobvDWaB60CLVwbksb04985FzuwhkDkBRvPtb2wRsl6Km9SQ+W0yndpKHBlY1OpG2D4mfToqsJG
1vvEYDCjgiK1F1jza/9Pu3f8GFK6avQty2kHuhJlyKm6ezVLaosdequ/bUKVZd5vBEUcOMjO2qPR
k6HWM30pcXEWQC4HLQlVFTKdSY1CmZhmDm+g/bo5dutoTrzrgKKXLrFV62+qgfBRbQtgtBQqAo/5
UL3uur2kL4/GAvzVNspL/95D8qHsS8sHO+lvEJifkZlytQUfQOpIr8I7t6rs4NHRKhHv2RUSyXXj
yx8Iw9orrhokgRcl6MIENigEZBBIcExb56avmlKaSykjxTFE0jofOypzxDZaZTtfmGKdgcjdeaHL
3Edg4hu27dGRnExcPiZEJQvuDlB5c+rFwJpeDh1l4RY88otexwLjbl1Nse3E0dWV+eIiDHPvn6NX
ofqdUvOCN2pbb9jxV+TLKWHRVywLjvWN66uftYPLkrfnW+Fs+yKlBxrh5d6OOWO7oEdaHa+IQtBk
BV7uUl07AlkHAu4+Rs6LVz95gU/1dujYwX20wrPZxSNObxf+zefXbnF27d7xfJgurh5xL8tdTNrZ
nmVlFIssCO0ExTiALvr37Eo5D9GzrBQOB2Gp9YKmpNCdkhSf3B73dJgMLTT7twYv1yqUZwg2yxoe
L5pOk3hkxlp1SehEiQHcB8xcDn6tm7XuTtQUFYRYA8B/gMT/r4JgANBSRuhCfCRsueyAfeNFZJIx
+hUIfV5w+3cwdvQjEl5NphrNaYzzoaZTETUUHwlx0VrOltin0B++j8s02Ul3OUO2rpUYi44fnzo9
BzgLgirpLGV+nk1HDinIzdFbz65vWSU/Y+qB3RYXFqg/CG/Hof+/n9X+FF2kd2bEVwpyObkkdLVz
JBUGKrwPKwvJvpQ7VzqCCPSYnnCWULCGmFrbcQRT9W6EdFQppqd9M91Jj4MAoU31UKp3KVGO42o2
dzlL/b5tFLbaJ1ync5lOwSwgPDBIpGRCBq3Rkon5YdZMxNF5cMtRbPdj2bXwddpnIBVaibk2U454
/z59GftBfs5AAy6CS8G7/fe/KxHoBgyJH+/o47t2tHr6Fs6EHBJe/270eLzTo+gWl5prBP8grecX
1ptNHvr9HFOkPEUDIMroflJ48GP+kYR4QlpTT2ecj5KWwY8Uarwouf5D3YQ/tEWZobuI/cdMUiN1
GJBGjuSX5XykJwzKumYKFPncG24/23jj3STWCIHhG17pxze4FEXNmLbfolB4lxysX5zbi8MZGOl+
pwz/uZj9Xe0y0kFzMBaw2zAsR4IvaIQY987P14NhF3RzFviSnyOhQBADG+4Pot1/fIU8YnGmr1M8
4Udm4ARYb6KUnTNol0rYc5V6teLgQF/4nLPNGphNUHfsO50pbdsyijwhCr/1Jdmo/xJJynXkc16D
Dl0c2jNVOSprpHSGNwv0dgeN3yhtvUgLKmIRJPxTV7TLMXnD1S57JKMCDx0zURYewGQvnJpGuXrP
YI+t1w+EwJopNw1fo/71f0N6c4Bfg6Cj512MfUBlRzk7iVEb2i+Jjum1G0PQIpXExbk5c1/tJg1D
uUvSS5Rk/HCIgffnw2aQgUIuqP4JXkIWT1xHBhm9HImSxqsa52BFXk/oIJs/sx3TU2xc5RAcNBhV
DtQmX7OOgl7T9uOhNzzzvGkX4Jj03nWduhSPtxC8Xa0IfBLLMH2UKNGHNIBL3nTtSgib0LEHuYRj
vJ+R+0jVjHKDvUAETQRyU7UQSswfI3EAJPHeuHGiamgeUB4HO/fOv2CsFlJ36dlfYZKcgbZ/PygM
+yRbXRiOYgWvQfLM7J+4598bRtowXdGNNjrUYv0+UTGpLDUiYlIrvPPjFCF5trebkCyxX4crWCLe
q4YMTvfi/N2/EF4/Suadg2z76rCou7q4lZelnSvJExaRscAgLkMe26qJy6M7VVw1WFI4eFUwFMUO
OVgd2I+K3ALdMy7LESP2SA/MZbjTeVvUkPIK98odkXWU8+axCpm2SwTTGta6j/5u6CbXjisoi8g2
P0FhIeGnScNw8GNSiXXDc6kashH+DwvSQRUs/gLBRdm4ARwhKP6SoSkSG8yBFFkwpqJevruqi64M
9YUjdPdGf8DZ65wclL8x1EmF5T8AMuBnq+ne4sZcs9AVjtpaoBOOY8mMYf7LrbD+uKYLtRKrFoEK
t09/Egg8BhUvVZC286lVd6mdSywr3ETLJDC/tIDIeycMc4A/KfZB1yuAjkj3VdZqan3tRJl4GjTA
4+TXJXzkrExBP0RLVl/CsqJtNQzi17lTGe+bNR5IGiYYtgxbPKeOR3F98BA4kX/g+9mqJCNg6fpb
e7TSB+mgeoR9yKuoHOvg4+KeBb9a51TyIgrbRGOyGqRy8yuBzhVFICjLgLRMBE5wIq2w5OFhO6Bw
XfeoAV8dssn2+XYan8iH+w9x0T9GWFoApS3G9JXhwqvysNGOcwM+/oquNKAuk00tX3IyHFsNhQFe
G1OSBkYRHbCWMwWN2MB39lNi4Xt8v3mCItz8mbTL/AiO1s7y1p14er986hLQGZl95fhrvuQBbxnS
7ot+44E5RXGbya5p6Ls9Y58QjQma/Xd1/l/BxEQ1DOEc6XjbXrSJIUaUMYQhVDCjvOakMEX3jFsT
OlepKxUA2eoPN/JAFXz6SpglgqXfnxVKujtymrYDiHZ0P857lTNp6ohTq30u6kAZzl6UV+jEy+gk
Rc7wNeBhQwPMM6oHKVVNqSk8jxSaWuuVkOx4saJq/yWYbj87RV3a3fAjUJJchXG7E29vhIdLeWWv
ADBkgix9uFrDtE783JCnn6ZKJ91IvR+zxk69wCcX8mgAjr6ifLPAma9ncWa3NX+UP+96QHOLiMaw
fsF6KV1A3BcrC+yD8/3ZVNKv6aV8pqCDp5tafa9ocnOSgs8MypiMgFwEHBvUc3J0u7F12Su78qR9
CKxW6YddMjqkFQCThSgncuFWBhFeSL/hWZoD4t7Nnym1EV1nbE2QqIN/iVl8oJ3ZshYVTYnVHc1w
aNNpyhGN2l4mPQdeBUI3ou5FDcVYV+TOSqMyqEw6Rza8LD+P7CKu17ZgOTApA/JujWeVSKxaHp25
JAMsaeR4wQDklz3D9nAQnw8lR7CVsmpksluig3CyTEAc9i0vZ7rySBUbTjBYJvs8xJx5Zwyor8ex
aE6kSxIFQ3RzAT0X0459YznGvpLZ0emBwLRse13HaCCb8mD+y2zq7a+3xOhi+CV5aWEn+6SNPF7A
EC1VzLlopdxUQmhRasjrx8XMuMv+Rgpj6ARA+XPYM3ih1ComA1j7agDPj57TvmwOU8+Vvhf9ZSyg
QIQjT3plROVYBSJqjjkypTHDZt1ld2I6FbSbMrpo6+Tkre6k3zus3r+z7SpaNQDXj8t/QhZmuIHi
4WSc9HxNOsKs6y/fXPplWDPlend0Ki/+I9db3CQifgmlMTRWnwOlbBPTUueuLoQsENiB6eQnUfqs
D+rZNV6LpaRqXFckxYxgk7h5T5HNtPtKk+gsdTjv1PvYqmJAF435Z0KrCQov5MU+UnG1twNaPGh0
EUnzKogtADJyIR6O3IoFQIp0wJ0TzOnYjO15g3wJjqDzULvzq8pgWZnPbbyQzTG17RfFoZzRsmUL
oK8W0leO9C2+D/u4Jojf64ihl+d6D26VXTU6lYiEEmx/lOA2vEn/M9OkXBKRd8YH2unbtmAdCU8R
j+24LJb0yPKLNoEVfJKTnXaZY9kIvgRSfnCcG8Zqq7R0kuUa2+N1+KbRSVkde16ldiHVVYbXu9yf
JC+aKNNJkFoH5LIEihn63cY2PIqPSQ8EzgxWkLjyhEsms6skg8/egJGVHde2G5c8nh69ddghaMlh
VhTj+ZByokRt/yFI8vZMjhcbQHI5Weabdp4GG2XMzw832VF1IvEaTKSQf3IcX0CK5mloUHgQUoy0
lL9Dq8R3xPhS06HHMa2HtlbM19B0TKGHeX/sSmgzRKFTl0I/tAV/Yzjtjwph8SU9dZXuiROCJKFu
pA/tzgpVYoBKdGfZSRRcGxBUlZzIEuZJ/TCpP3xlgw3uNoLbU+NFZ1Bbg7S8UDkCToYCf6QYVmoO
Br6gnVuU2QRpoVPQgxb1VZvn/W4qVq3/+pA1tVQTJZ2tuBOGIjNJIFsTHumCl9lfMtsf1t1yIs8o
uAF1WXSiA4hhwGqKx5fHnG8ot0iwY8lZiurCktd9hSfZmNO3wcIOBluFYuWCoQMDMimNYoN8MvQd
c7Wc+IGWVvU2YtXyehjeZxSzdHyXwSq0DsQMBr7D3r49xP+mrVECmQdLljhkqWo3nPQPIC2m6Mt+
fk+GamLqvHXK9HTy6CiOTzDvU0irDPpB3DdFZujyhupKTXGTGAKeUdA7aq96Daiy8bCnPwETZzo3
QC+wGvvbqx402W5QZq0oxc3zA9+bwJnRjH58ECKevams6qQm7bVx4aWvxgF2GPHHjyz0PMY5SG3x
p/RLac7mF7oAaG4jq2n3QaDJWIZ8qhmsjb7iMiIZ/x9xfkz2gKdGmLWdCQRtMzbrcDbGpAfk2Bm6
Q4pn9zPQzKct5yh6em1P+s4hSU8XD5/N5s0KnXq+FtDBNxEj1AfCcxM05+7P+Mr+QyqFkRf757wJ
0F/GUYEjjq1lQoPZ8BN+27jmf/woUVWyxUBiai7RXUa33PcAI9bXbRYQu4tC3XFcLdrUY7uSla5K
+qkm2mwsNBEA7uRakkuZDjukEFD3AcrmfEqLl6dQWZVVZM/eN95qBwtHKyx95cJGTLq7k09xeA+2
Y76HeBCW7/aCWUYPOjRD84OurPki5963uErvlQ0HCqoVFIXHVaPuKgEqD2aeu849FZ9wunaQVtff
X0XuzEF4dXqHKTfWfp61cRM40eQqU2XCWg9XhkFaE54H/PtLmPQAEUpt83pAKqH7NKFVL1XrYZIH
N5PwogtmEC+ugxUNIs4r/xLIlzTsjdQxThVgmF2yPxNwbNYo9ZcheCoU8iA/Ofw2PTH8Hw/rxtn+
FKPySdG2iTwYuze0qTrW3yapOYB6KgVecURDVObEDfIk9YvP+J1Tg6VYJHyoC3TcCVm/TgxR+SRH
OSt8PCxP1+4GKx/d123tDQcAR04lJppgVeCMpWjk3eG/EXWtJ7izY9VKmmwOlUFc0R9CY75lJ2Ie
h4OcwiR/BkY88Pn58XPjBfbjHiTxdZFN0mHBN41RsvfcRQLo+nYmxVxgnz+MivPOiIRzRCUmrN5Y
jPxzw9hOgzchb7S1ZDNSG2ytQUWeQCVjt72pgnojtfEtjxmDqlmcLgkth9i1JBsasSzCoiaImUr3
sY65XtrrzrjcIXZsrf2/KAYAB3iaXoLXCx3umvNWLXwwsunPxQXkZFusjCyl/T52OvXQoC48qZBW
HTsgmZlpoT/yRMORhV9XPkqLp3oUa8zna9May+xLUu/WC1vZE6wukFMCK9x/Lb0oEPlkMwnas5Jv
HZsTrD/b+Fk+q2XjTMcOxS75KEoeN42B7muzaAvi3F2gEGDLzLG3pvbvuu41EZLKRRwKV/MaMiVa
+lxQ36OGjsg72fyVg6WrZgiLNc8S6235junXT68RPqVbT2hjqLHLnNIEmes/s58iCqsIs2VXr5bN
I652rkpOn7RUHI8WGxvuR7yURO+9RS3ePUtJ53lZWKPU3FGCxnlHzP+a1RBaqQfF5UoaIjHpfnlK
Wx1uEIq7g7FqSiU6IQV/5H7O8qNIhTtJFgW1ocS0MVD8FtTJeC2Q3f0PXh9p4C/UGq0g1+YDCXqQ
tiacCQlEQcxkU8h1undj9tcOgbUsMyl0JOKK3U9MLM+eNk2L0CaLk1m8WpNR+awTplXhUmYEVakF
ARxJY6SoTpPOshNupptKnZ68pXQkFId3W0OoUMbEJN+dFK7PovkkO29p8VikzrjdHRE+Rp123DH8
Sc6cgH52i5ucZCBDzW9DyPktFUpN53uAf+qGAtF9iUoosU8cl7yAz5nffYdTcaVWgfFBCSsileji
q+xuvdTw3BdqtBaw8BzLodu8DP/mZrvjKcdT3i6J6EUXQV+aeJNB1MuLKe7BilyKruxJteQDGSYo
iHlhZ5fXMTBfm3rchSdMaL9vqN3rK/AvrZEHo8qvomcq6LaseGxCSq+D57c5uy+kElgKSq0lOO4t
eUnCZOuim3rx3ADpHLcbwnFJRTFxIIwQzMWKVvXc80bdj0CjgO1ARx+kNwMtIUNs7UhkYmG3GfET
I35c4EnYL7drDrETO+sDFq+FyYXriylvOQDZM1PSa3FNc3ly5yL3ZQ8P8u37xRbLywKbx5LZaF6f
rJzUgJdiuot4qLgFNGU+nmZGQyoI5q3kayZ0Gh/0iY24DURHZwFP+Cv5sv+Om/ik1O0lzMo6hK6m
Boi3PLILW5fm5dibt/QLvSESw0y8aWntm9wcB2WoQNuK7dJ1ZX1fSfBp5Pt91Av5WhvyJqM/+hYi
ZcviH1ZVm2Bchs3TPqjWVRrR69L/O/WYa1r2zC7L/C4W3/RXnFJlkQ7kzHSlVJ6nTGtcXqvbix5X
eZpLP7NP8/tjKE/fsIiBQSwAwdSfG2KxZRDlmhQ+7R0jh+iv3G/F2fuh6BmPLZ53D0GrBVUJU7pW
P+dzV73tcnEkfRqMCZSiekwAcYAUBaKFdTccEg13UCRGSAL0qnif0wO13VwzzCmwjpQUME2GWDLb
ZwrM5qyMAEdNWWkBd/lr4R9SQut013Htuf+HChCEHtlfeH67b7EuySwji4T+8MayPzz/gxUs129d
DPAfDvTTSr8TVKquWr0OCiqG9jHHlMKoQ1vFkFHtQ6HK14D/1eB+3sp6aHWbKXubHC92XOlr1qeM
v8SYdiqlMehGfRrfNdD+XGu7KYup+lANk/EF0QcofKAMHQqOBoH2ZIGCd/9o06gOuPIGbpb93Z3W
HhPszv4JeoMIWSK50IYecRTFIFijoII0vynR9ZE+DPSRoZN3JVrHgObZAy6rvmQzVOxhSpSeTW41
HyNVzt7kn10jfm3B2p9qjraJkt5o1tm/tKRxy2zdD73BtXgbz/g+vfoWmY4bAfES99h6d1b+s4Fy
x/n93vbP61AQW7T9+PuFyAlhKxEWQxVISAv1rIP3DAljepsveFfsgCAtXJ1w9XZymYiV/K0uXgMp
hy7FYIAnQyN9n0rS3pe1inmbfReTmkICsioiiiycXr9PnoR0YVJ7tnmTB9EQYYvCpcs6x1DhXLuI
mrQb+Ctgd3okDkyfnden62vMPzsxXgNThmCmvT5lIVCx4dONGWN2P/BnzUaTxYjJvwpvdS0i6oa0
DSnhc3p3EGqQAtM6indXzOagIpLrG26HLExaikWU3s6zgn6JjN2u4zxW6wk+XasNLxSYo9H8rSS1
OrMWozmnPdTY00NWGtsM5g8ioVD8rzxFcUwdF1mFziMnZ3PofvNvUDtA3Rykf5M7Gxm1dG8sFzCp
THOHM67ZuWSeVXykOO5J4HZEtIUJpjgU0Z9kF4OAVD7qj1O8ojUsjK7qHYjvzKclu6EwwTRYBr1R
j4n25M1OWqax5It3m1tmPRFbAnzlL75rAdkNICSonVw8zVSXDPScE8AGvpVuFcVIEl0/7lbvD5xP
3gmdRHKLOlE3ftKIIzOM0LOApRrk95FQ8PekyFeVMm2k0++8IYy1nRrjyLRgpwggiWEu/q6QLlJL
y49OigM32w1JoUa4byzDd9SNvfeD42Kqyt0jWK01PCY5xFzkUtoLxoimP3bOPHkWPIlHM3GKwmDr
tTWRji6Zd3Ln8bXp0Tr2BuFdDKeD00vRrZBu2tfeXWXofzuo8Z3H8ydmOQmvrVbG/m4F3G4WyfRx
XLI7Ex0iDfdLwFnL6sySf38obkDreK5bp2iiHCTWf6HjK6RqnUpZSjuWT4OWiTfQ34bQduJ1DFZC
ZY7UCj7HxBkvd0snZUCHrqCklQLsG/NM4CtIn4gixNNhl4myf+8N1b6+ngYYDP75gICpZL88InrB
trKVTsKGm5PNbXhY3Qc4gbHJRqN52sDPvCQTqhq/4jP7bQr9G8W1+qgL5ttn9g1MRSwTwPBnBsrf
qIAZYMLKV1O6UfJLGHm1Ad3THVjMsGWUdBHseLaVoWDPOu8hpIewJ8la9gTn7s8e1GcG561vidO4
r8HD+AyoNeW5j7UTAGxKBRzjkSctRboc5FXzlk8Y5MlKF5KjerGW489tELeMUz0nYvKXjX9u6WZC
7COwrOoWaX/4oipEBhqlmxtrFA/XDIhFELFgUJGrZiWFmRaL4urwWzg+eoa+p+TMHcUPevaHKXQq
AdAEToOIiVHsVqhEVx3rb1UHKx1HzEClqOSPYcr9SwQPQuYV8WB7wWb5O52TJk1ySx4NgvmUfW6+
XdqFWnBj3mEYue5m5L4SKU2SDeNxOGd0XDFe8mObU8kCt8fJ0sIGLlkPi27FhPQ2648qsVN37e2D
MaSIz5X8B6xlHrmzH+N7KkCxG9cQdpg4mGldL+5FF6Pkq8jcrx42fAhMCtP+RoXys++vg32grwMi
eHHLPigg5s8G0bDq1nQOxz77KbvlhBUx/BKLEj80NuuZ4n25QqUibnH578bQYNONjLMByKsPBpFK
ia0KKF2ixLXM6WbHDdVog9PTSAyCRdINNVNxvPiHbnlRX6laVXfuIiUnJAqUIgsfTLzRdnSyZHlx
sS+hg04qAvzBYCxjQKhMGKwSl1TgE9KYpN0D5rweHl6H260i6L4BkbKuetCspdAP2K1Y+7p2ib6l
X1tKew8iNsZPZfNPjrx0jQLODohr6wakkrPyKTTO6+TLTQSRDI7lI3lvbOTB/Uk44+DxY66v90rH
VDwbdez+H+jlLj42V+EjmO95pKiNLE0d9pNtk8/jP3Rc70jIQgQyo+f16YXe6em81gRpesMdzHoV
bEqMOpQCAL8t4V19dHWkjYgZJUAU4rpnfizy5+0N379kj2XQBB0KDi0KvgUiiPrxDyZX0+YkLb+e
xb6FdyjVecWtNbDwAo/ctx2LUumdQXRF6UK6RrScGFhIXK+bKer76+xRIXjSDBlyTGg753oOuVim
vIC+VKu8/53fVSfx0ahqV9SY/Ypl2tIBVTan0bQc0vCkijFKDJTVMznLhqkgOCaOLArel7Y9G6bk
HUvUOHWIvx2jsMoIgSx8F36wQ5Uu9rdWgyVrNTbdaiWncKPVvewJ7ZhNbRhLRxBS4egWsi+qcUED
iLR1x5xLpCosTOCT0ejydrCAoA54Ykq3bLF0WUH+stRCXnm6uLMdxSFuLr3ww9rzRfbqvHAL1zcg
vmaZNf2leWDRdSPTzjfnDrFKvUSnCKimJcS+d3kA8H1e6AG6al5DwU2tCm+VWWcL9gnxP67HwsCz
iS3euApthXGPsG44nLbwyvLmJpodPlz41FtC6IDqZwPa9IMF0ZSjSv3AqCcgTrb9TueWQ8wbuCAm
UUwiGAoMj18ibeX48ZEga0qGxEFPiEEE1xBIquf7+HH2z3pPYtq5DVsFxgxeS0XPKA++vksr29eZ
P7b/XsY0ppMR5I6ioLwcbA5nEdYw/LToGVn3p6KbJnTG5oFW8P5yp7lvW4bZQrpUsUfoBl7pjCz3
OwxLoGxqo+Mf7I6vTA4SDX2n97xTZ96NbJj7fxLi2ZQYS7tgisKFUKNf2v62nrEnruNRQEIOPGBu
/ZlUleb+x8TlG+s7MC+A5h+WWYWuLcaV0mb31L4P98eYhnvv68wkQDECJWvhJau4M8k8iKMqZxXw
hMfegylKQh5WqgclAdR3Sr+wYUfZs6VIROszwwPjgp1dgxZ3/BgtdpG4ktFBiTJ1n6DeIGz2TVbJ
5AjqMWnrHQ6/4DNWy8ObCTx5JSKZ0OCgu+M+4iZIE7ey2h3eGtuUg4iJ6R4I0DpqYtHMLLs50wpB
tw2esfmXgO9aCUiGWowQMG16i+KESrCvls95c5fetOPYyWtBdYBbyeHeEn1v+3HFGgWmhHYwSID4
ecoLVwIT9QW34Bs/4pSNYIpaEH5TlTHk861NKQovm39G9LJnr2JbDm8QXMjVevsz6Q6SxElP0FYX
J3RfeTzednJyAbpn37vDbFqyxZ9TU+VUHdMMqpsXDEtkCmMhNNgxG6vraLZiZRZgfxE2X9NKL936
Tuk0fQqiXk0R5fgjPEExHk9xLodZOMldvRiZ1XfBOvp1es2X8J2dmc42Yn5JPkYollSII8+aYiiL
ehbUlMGxmakTga40PRB1TAspy9d13eDlxo+WJoBLJ/dQ5VJ/GV/++5gsE09G1JfzGjvW4SIbVFNG
YFjwizt7xihwy5JY55EeQsl2AJA4VeLW8kxljRxBn3wUMaHu2SiDk8T8zGmgwD6ATeXljzml6fI6
KGD9aRPCe418pAd7aO7wqO7/HAu9F1o4WVlZDJ9CzFCUUUTrlJ1s+pUHkxp0dlajcvXw1EefQIOA
U5ktzP/PN9OW3bQjeJZt26JPq15J9hVBdG3l7FV078VCk9CTK+TvC1itAQocsxGsOkdeDyMNtB8P
shcpHdv96Le2ks2XH18SpPkkfeN0hTEzLesuvk2PgekslEYlvB5TxpjHnzqzx7lVkmZXwAnP+pTv
phtdH9SCMqkUaJYWLA/duRJq1XYbY31ENuCeKBhNXB+dd+IZwXzyzR7vDJiotGKRRxcq+6S9W/zp
4tJNj4G1S1BIXawJyk5cKJtiQitpvlvx28uHjlNbvO9hJfNLQdivfzhUbTo7W0cXL+0qDjyPNGPw
jdebjbPO9ZwYjAEBpsEJ4E0UgjPDBlRfgc0KiOBdriEzhzv2fs3fV04QpGk15vTdRbMZS+hVERWJ
4EMq8NGxl8nVUqhjSGKbhEVkbwmMW+sVOBEV70EwEbXZDCrXiQfz9iK4/F18y2WJuVhQQwvxnb8X
CgIdVcL0f8il+elxiIGqiRXwLbC39H97H4JdNlo11Ee0OW1uTTFZa92mpdl03sstAHU3jfFzB5gD
V6wBFwYqGHnENKzWI+wNuQz4JJZ9FGBs92TNQPOBrmRs+DnINsTaUUrWOqdpbciEx6GhDQTOn6Az
5WnrfNohcIGqVyn/qit5txUf1QwRvjv9w/xuTrd5JLkNtqB8KHk4KyGgKdmgbc5TT0/kVbvy3xiR
HlE8aQrXvg+azztvsf7UAkSoMuKRp3/3Jt41TARZQXJqcyryiuhKTY3Wn1Yg9o2MJJhQyY1CUOFk
8WeuthU5kPo5fRtBFto0UzpIZTavOhR+6rvqbubpdllr7nlqf6QQfnG1DIRC5keciyAb49k+mNmg
5FvwgoChdyVTmqhLa7kavCbeLC1TEhP/wDmPVu9/QWO/arWXcw385Ld254QB/4G0U1m4RVWbxd3G
y93EwkuVAXRdfXeKgqZfxBlNYh0J7SZsGGbknkBKPLZMAgnlFCFhxpqxmxm3G1LJlwj8A6w40DIl
VVTZSETqtkj1+UC9ZKAGOvaFIR8x04xcmZgDAWulzYBd5ScKdrXmIseSLLsm6gU4P5/ZuvNTGXq0
rW3K+NFk+XuD3OOSoVIAZeq0C2/rX98jvGpiZEarIHHmYf7nHxCYhHlisqp7siREESQUvrnrnQGB
CoRUOF0pMFyChR/IJOomSSVtmSqG2VNsYI9cz2XtVtpIrpY9pDKdrg0vJ68QlRbApK6dL1zXOTiG
sVOAFyt8JIipY4UZqrYwUa31AGjnyzT8axNbqFbGTSE+cYKtTFe0zCS1XWXbnEs7asKG/V5IQQbG
BBIvEjPBpxtmaeCtZx6IM1RKAVNDxlczenAjynU24106i1i2TMH3ANddoJDlb2DjJPFZ6KhI9n04
teCl2byJonZcRluXhWxDqo3kK/QOj57/QYm9EFQoGbgzDICVPS1f1pJR2LjQDLLa31hCUBQDR3JY
/JuWgbtO564yJoMN+jlWU8HbDT8ugM74VI7hAlGk6k+sEqOiF4pNg4blc5kR8YKKavWyVm3s8D9d
UMGvBRjDcIIoemEeAmOdpozH872AZKigDc4pnACW0bednRqfpTBX7f7iCTdpGARfa7qhaVQBZgvD
xYRh0pee5yCe80bfYaUy0gRLXFqNycMvnPiuOmK3fzpBvCRGMsUJ8afALX3Xr7iwvy4AcEoJWleG
lF88bDx/9N6/7ACA9N5o9A8rqkvSK6F5QCtkdBMNkCZshVz3/ot3EbzIY+gDK+IfOBI/qThJtcFQ
9IBvchAoDC4AjDLewLl0MsvbFxOsX3d+lze2vPDZIgx1DeHCdnGX126gFwWTJEHav/jGLXngzLDv
iIQYaPuNSms4JUSQeU4c3+p5tw7P48WJyFSB3StSf+NqlIfdN9ICiW/GlZDsouFPyd5jkuiC+Baz
nuvJvadr7XpmhWAAnH65jx6g3TFgUhQMQ69nGVJBSKUC7kWbSjxCxm81ZUBaEOjn40Splf3CuDhc
zFVkVW8JFiojBBywFHNIGyqWfSuqssnyg9pgQaP2huH/HMu9hqO80f0PVOfwZOBxaLJozHUqbegp
Rk1BxG8047vZaQRUoB8GWKmnkgxuPw4xqfRL4GQ6/tDTuWI2udHaDbUfnPxEGhN6Od9NkXrW1hcF
AngpZkXy+cKYS+xRDXKPJLFcpWqIyjngwb3f21GvcKQNogdKbOOC5+cheaQVAX1zCl7o5gOpLb2T
7bv82xy159RogLNzeSVK7BZQvpxlppyCi5kAe9kRTuMLwg79BHzSgAqWboMeojcLnbB7gr4F31FT
dcj+RttNPzmFFffY4q14PFY7U/VjubI1O7qk2pD44dbNxmIP2vQAMW0ChwRmGZs8AwPTpjjTaqIZ
1WrtzAdhs90O50BH4FyEG6s1k//HF60LWeFmIGdtqDht5XhXHVe60Fte1lUshG39jPbt6FWuQdX6
r+YcoMLDIYyFTrYG7BckVcB72WrVFKj0kO2scPMPrs8n4IC5IgFsWdgM272AP6+8BmxrdE+9LcCG
6nNfysrGsTbBqfSdhRBuue+eWASQswuj89Xb6aGKsfq2Jrp07h3nwDIXYL0l+yL6iGLXgZEJHInz
FQUh1TAbMjhAeEGpMiB3q0MMKDGHP/MybkVrZEs+S0Xrv8WDL6AA1Y7J59SubwKfFxClBdI8a5bL
hpkIoXOLP+KRujs6DjbhwVztt5IkcuKdkEuLLfr9NB7cZ4obRWr0pgjsVD0cpkPBeavtCG6KSpbA
lQL+Q6j0f9dF8dt3yHuKAecc6AqSDC2GyRQ3ou4fI+vqLfexxLwrVfKncQLhLmqWdAUzE8fR/EXJ
+Fklv7SRA0y+dh1U4QPlWBhTT3/6R7llbjUEUPgXfP8REeMkhlR16qMMiyumVZlqtw1oVJqmb/+W
99jjjWwD4U5xuhb5UoAuq2DVYXJ/It2o6fdWyMRRSfocLP3EdPj+e31L0VBA1/e/g7xDNKotcQrU
YFGNEMNdu5DlNAnUsAsuS/B34LloEONvmOVBjQWjh2G0ZWSLI520DrQxwd527BoMAzj7GGuNSNkc
CZWkvjsiF7uT5kfIT0eorbDa+fKyMD6xAKUfBLQeIAw3PQ9dj9sYWGByLTvqDkaERWsgmyfz7e/O
DMU+BWs6HR6t6+aigvsKZNlOdlu0tKUIsdNAcI/78WZEyduPlm+YrAWidjqMDCwB5d8A80cFGVWF
lcL1QCl8DGj6wSuCVkaFxxwz1DHcqM/UEpOgnsZBcnXwnJzKWI5uskv8hvTTxWPnMdIa8zLomTJ+
JMMZCyvg6+rKpy2rs+yUYrjpQqONPh/s3NID/hpPDXKPakPkvMXrYglP+2jfRvlktDbv7SrbeINb
asCSmw/9qAQlUuKa8H0huCAZ/2xtTT/o2E5PTzNMDdMdv1wqGx0vps7q/jF62HOuMEXX2VwkwC+h
2aywxmHqmbsW3lL3HusOS4gR4ffTCduuT4DmTu/KaD0teRnJBBXWny3llA0LYpRh3Ocac+kzSMYI
IfdyVHOJaIEZ7o2po6GKcRubmzKHPPE6poX7gbdlBAstcKp2K+G8HnAh+qJuGveXUFYvuzvM6kQT
+GOEIp/9KnGR+wH2JHeiAdP0JWihftgwClEn7v0IjRFY4iIyagJ00WAIIQuCvqCAMB8Bd0YWoIde
PLuJTLUM1RJeUkDhTNBSC4h/4/KttlcXMP0lZ3lRO/2DrURupOriW4X2t5n2WAE7whC5dNn6wTNY
LQkQzxtIkliD8ri2OSM3MWhsSNJU98n/d05WKeMtUuz21HBtqykTiUDtUzgIjWULfFLqYpV3sqHP
stAyaqHbJsn/kOpPkqQzCuU3IfskCVT3DNFYEI1PMjOhDdEdMAFKlk6NgTbFT046opP1QCUsTcem
AutzBRQ5m8S350hXNUwNbDZqQIoytgk3V4fQAtId2rF1yntrRv0BFf2EjGC3qWfcJPUvpgeD2YpH
GOmryqZBUfS+RaoZH3zwhnCv3+iB+aVh3kEtYpzfx6mVFVxKH/UG7Bb97gLxKrmc7hpAQhu0QUw2
NNJDbofkOP5RUlRsmjYT86iWTYt0DG7pvumc4WdQxqtEcZtHKe+QUg60qdKxxI/rL0s/iqwRR1c0
oSP+Pil9F7bRY5YQPPYHugCGc3zpXtk/silD8KCQU7Z6BsI4PKOqg4f2hPsa4C7GEKaP60+JzyDB
H8SttpSxNvAQ/TFi31sZFpfKVplq3wwDlvH4TADDfVL6KaGF90yyHSbyBl0x1SyjTg1nCVDbcVBA
P+SMS9Nr60eZzyRDTODaDgcMBCUXCerzQ0MNvWjhJUpiyv/G8Idl5RxCbJ0YioAovdiqAWbW/bQY
YnypAQCxFejjc/ceDDgX2HDZuNNDiL8eU7kL6efGzXsC7/3CghfV/WOnk4qkZNtCY/7AYsVFm7ds
5ekUKhN2hjaDAur7jGtWzle5QWhLVE2qPzaXRI7APBshOYBDRqYMXWwhr7+c2RIWtezB74jolHg3
/XFvMhWvH1If8XrTZBpFV1A5oDDbBFSgqkhvCnuZw88nLiWIuA9ghFxPh9N6DvP2y072HUXxasYe
14bmYiy4Ek9vun0zS5N//el3dj82P/jNiGTgWWG9yx4gOTl3Hx617v4eINMTWhu3yD52Jz7tdExX
ymtYXhTiY+vKmFM/pQ2Cioj9AfRLg3R7wm76Ks6ePCFVOk+Rwr2gtUnicE1HH49ULxkGAMnK3Ymz
UqusxouxXJRRTZKdUvdc2hyCl1LRx61lduQrzMyzSKrbt0jkZJuzGMaN86tLk1S7V0kIN6JvecbR
0x7H0oDr5hqwhOrzwbs4vL/6axkl54tXtZJLA/23GTvs2bpc9m8VGonRlDudUyz8L55lECgCLbtJ
faev+ekvTeYQC1iYrNy8DI5pCI4rukXLp7pwsSYn923jynYdh+bHW+aHJHrZUJpfAnK1xBBprITj
uxUCWkILIkneL3xBp/nk5b2JtvoqdnU+KDhLFpXbqYPSYiTjU7XDdHJc58Yu44zlq1zRktbQs5EE
x3+zXEgJMi7u1b1K7RALFX6kVDzXb9W+xWvxoejHKoeco+25jJzxpAWgtn+sltJaAQuzGZ5Rt2DR
K3s2hlK5S4OZn573JZNkNtMmxJJJitdbpQi1eU9oKtvKq/ST10gCzM7yN472vIWHRsHxDuWvu6rn
uvGdLEElpD1EIy0MVEs7QR1sSoEjAYViMUDcKg/HfvTn1Z5Etmui3WU6LvRlR8TnmY5Zzy9zEjWC
aTyiFAS/RSCMFyWKW2D4Q4sM0lwRAlsfqSGikqmJnolH/FqmHj59xUiHWpmOr2f64/2sHbo9FA40
fmLid2L7PUhrgXHqboCHPdi0jbwttR1bFWm1KG59Fd7bqkgcUIXuvLDWg4gvw2Vxvsn/pSjlnaEk
NQQ6JE5SDQ5VlQjGE/eOv8zzDY5now8HMpQF30h4vjdiCYQwgRSuhAK8ms1iEkhSEuH8FInSHgBS
F8zY8U1Xy92IiZixCphLrMI1Iwiu4Tf2Resf4rOMNtDIUwpDtjEPmJXBKSIl2H8IsqMFIH5T43II
HLY5se3A3J2XVelG/DmwpWuLzr7D09AFRYRGiAlnvmOPFi7yRglhKZzt32GaOJy67dSZFc7Xx/de
afjcKynps9GvulO2jZN2tfMj9rzt6ONCLwy3vYttHVYByFHCu6wQ3e3SdtHuOZWm0po6GsGAHDZe
mxhRurMq39Jr90/85jOd2K1OJTz2L+4/mE20felrbcVr2tSp27iQKJbQVCgOKH2Y+6WUW6ELQ7lh
BNSHLNNKQ47K0GfmLGAFeKCGf2j22AT/GxksIURbd3Y3TmVS2ZVmko8hVel4ErkJ1NGz5x2/Ox9d
T/3jjOufGIYgbCWZUbKVCecFGs+1HIse+vCCFNMT0bH1Orrsyxlp7HL2nEdzd+KcwgDzftnJaqlF
n6icX21sDdY5E82zjd5QYBddExMpa927VhJFp2QAr6/U5mT9tOy9xHUs3h7iXreAroFA5dOP8qF/
LVsVaWCR2GO1ddf6fQ6daiet/XApLmak40o+z1mci5j1QEhnpMMBwbu8bMEo3jMMJfaBtQ5LirMe
Nt7gDG/rBYlm6b7yO2+ON8OYDnbJtPOjmNSnR220cq5nO2TC3GlDTfZsfSr9pquhaTUJvM4xA/RL
kAr3/x+BXq7orcnkQS0h/0KRvUY+0UMTzbR2pdxwCIaPVYTqDNGsNebk7PvV4H3grELbUOwxfd0y
kIyLIjW8SouaBhBUffAUkZIttM6/H0gB4zT4NyhSeiD1Lb5dviKYBvShxPZzIH7fGT82z5aIySyX
OyHkFW02KKSfwKUNZC4HSeNRgWdWLB+38vyX8Zj9rnwkS4O7r9AAKaxHwnUy29bBQVHwgoZY6vW9
ifNNABMNiSWoKca9+4agg/1SbWL/7eXPe93gJ8bKMdqj/jXaEL5WDJFYbH0ds1AsvFkpCovYh0RK
nABnJ8734LtmQrTtLHGw260aT4p5/Gbl29oY6ySp1sTNMOv5WaKPWaBvObBMztjCzgXpTdcqdjT3
zTn5TplYDQMhIshEVu8uwKRm5r2k9vWGMkcJChohIE8+rhYx6YEIEdwnq2rH3qmPTE6EwUPIaLdZ
PDjEdZpojePgghl+QJUSgLqnQC5iKeOy56ZEWmnVRb8t1jPDKwwlhfL6ISP4w8GrjsaTcGpjyX1u
r7N1dq9VMbOnhuZl0en2Q41CTk+i5/1xEmNB9YG5Wckwtsp6Dp3EtOKk1Tx0Br7L10vh9AQrpDrF
G80dF1iqZPUWJd2lHAdg5ccfRvJhx2EToIF9HJO1o0fw6CFG4mMhS4kTqnXj8AHpp2xotoCGyCL8
ayvz9YA888w7noS70nSqR9tIYWA9QvIr9uaPaYfSA4RvFcQGFp3tAl8BMd4v3Ym9vbE95zKDU7uo
F7rr3TpP7k7oMQHnIrXZvL8TdAYMKi7Qq3SON/0jC8WoXTiJKjD6/ahKsiwZvV6i03c8QvFxXa6q
7zyybml2l6EeFslx48CiMMRW5L3RnCoS/oDeHlNtwrfYG8fnvThc/rWICciXytGunrNEiLCsPvTi
26BJbNZAu6Jm902FIg2v5ViJotW3GXnHANiZ8jzvm3yvD/Qp3L7nhYisO1DKnceg1doo2VMmfiiK
vDDGMhp2zc5TbysYgRTyRcp/z6Oufie0zpxF8N0P/Ip/jFC5p7QJA23gm6viSeMzV6FD6QDN/a2Z
IFo4CZ/DuNOwrhXLdAib4u3A13qP1SsRHShTUx+urD+ps9g/WcOIChh05z1y+obnqnF97371+pHU
HPkPGsxxdSo4xiEWGqcvfFeYkq0vGIY61lM6unAFtSzSv0ZUbmNQmKHoB+kE4NulvD8nQ2tYSUWM
Jo0cH0TdtWhFWnSfnvwwL80Ip4nTdUuqywc9Vf3UOS7qmgrigmh5FIh2k//F/e7wUgrgcsdWTN3W
4QPuKCO9SRwNLnJF/aSPdMJ9PO8xm28yJOXbehc591rGpOXqGeXyOpn6EInXZfPib5CGjs1i20Ns
JPCz3Vk23vI0wBAI8u2I8iXnHt03ZzhOq/dBTXnwPluI+0sCRRPysulpLAq9bSmjhJeal5bp0E0k
4BO/71rdDKuY1OFbIjy2OHO/c1jKQWMsFYhfWyU8qMAyTtdlwy6+JSQQnQcginPytrLk/Ie1IUP9
bJIiLS192k0T7EFK+bYI95OBfdwfOUwx6um1yZ5oKY6JiZJRUkeSCZvWV3MbyA/oo+wpROFge5CF
sRrNfI0V6ty/4ak/DXUyi1E0RB4h0bh/YaDzpTnuEKjENrjgNIYWYQRDVqBJNS8cTHSsr2LbfFm5
P19d6T7kk5fw1TBnECi5FUv1tgk25nMYhlqn5FEes1JjrplPA4gSV/xwIcfHp1q7gJRI6fdoSx2v
H+C0V49ectFDWC1I56bQvVCOsIA6N40OCrIpjIbdC4Z2YSv2FiSw76NnJNGWPoTg6LpkoiaxSXcA
110HVai0XynTd/kLwaVG1T4dF/ZQXwc5OK9r35srWtPGMt3iDlvRDvjq/blL9fU8Qr0LH0lC96hO
zhSECmKJSDWkUZQ+XeVQmA4ULAnPrRf25OpCNaYGpEFoWuHg1o6vNq1nr9RptNlNDiz9ZryTMOxZ
LfOO56GEofza/nTNdTmfqx4MGzmQjEiSZ8uDlmbE858V3VFu1bdFYErf9JzgGfDYMl3y6UjqpBRl
aJ5kgHLdEOil0UlAXQslhGEPIRVfzI8D5RI+Mg5y2hv+7km++NSoPsXjlwnmCc0yK9zyOeTs3XCC
lSmB9qjyC9YVsYxAGvAB2hDaVSEl2QGrfyJX4S+sq9/xZVc3vZ+kmDwhi03lFOmWJs1h9inhQGx7
5+VX6+i2AmCF4UO69kDlXSJ4f3vWapjeqmtaaPa7FS1xFgX91ycm2FMu+sCZCenU5uKgD4L0WnI0
NqC4Ob0talIfKMr6GoqDz/Ddv6gsFp2tjUqNI99mxzdTvV5B/Bkht7RqPmt7S9/cf9cPqARUGkE+
41yeiNDCTP4lS6mJp0LLUG/ayDyt94F+0OeIwNx/savStSAIv9YIYY0SMaHu2+VWP7h0ZMjuuaf/
dX3srX2jg2OPKQ44ulHJHBgg2LmLCij7i+7+Fa/JIi/x0egOgnSAceqr7W27Q1q+7gZfntLF2mrl
/arrKTN8fdU45/Pm5yG++8GKt4rmc3CX4kSogemWA95B2JUSLme5f6m+ZKp4qZC8dnYeEcZJMZJc
7poZgC3cvsRnwsV0kpquBRCWaYKTx+czIpC1D22mIQH6E4mC1Y86A+8sZLZk+1ZCPRzPzQNP/wxx
LFsDxo7eEN+OROWsS2x1H+8JHbwsUjvqLZF34YjiZ3WQZPyse55lVX/mpLu0//T1PAE4/gV0/DLe
Nf783EzvQZSZgxV8ZYf8EdLrSZIpmOYm/gpy+vxACYHHTY95McbgtNQLTJKSIrkVrZPRo/IGaYhP
4+eYwXGjTWN1ijgQgKZPP7k7SWIndoV7x8xM//jfUE0v2c/xW/y8jlH7DClwH01VpMr86Qy0FPd2
Gag9RDzJn9RLV8TDWTxL8gw0PdRdrn+z8pBnuW/H0fgQPHvCbChR5m6BHnyTZAAiGkq6+2H980pf
oHdUi8g5yJtKAwZ/njv0qng9Pzpnc36ruk8pAnkVu4Q4p+36W9L7sTTPEuzxIvwmbHZw8MrIVXP4
wJH3sNmkguF01qcG8K7QDt/BhgUpQSDSJXr020vcn+RrXcmSwQz+5+E8XSN8N1MLMl/bEZWN8351
UbF9YrdUnyypF1PTXKeg8r6O84aUmGzrN4SGg+UvvuaPxcWjmTFnFtxu6mRKPpoZ7b38dMVWz9jq
rYJeq+6fP76etBQvtA1fFzX5nAtQS0koCscNs0QNFWJOoK9tNj/30grOwe2ToiIhFSL3ryiWREQR
zydrepn7SoxumfGG2FRcpaot3ukkbWBgj/rA1sedXyAQvvnCJN2exy1EuCDq9Tev1UI5p4zBu13e
5u8HVU+tatQIkTOvTg7rIIPtm/lV19RwLOs7zpGX5UAJzO/tDXZS3SNK3rD33DWQOiWkX9T3d8/G
/Scfn71JSTjbgqjomlsRHihuEnIT/qwDNpYFocyetm1amDYhAgC4jKBsHAN7bdRd4MJAXSmQ6zBJ
FmCheD9ZGBxm4kjWkUx27PlpfDVWgXWL6OZDxXTOjY67FmR+5KsqvBbCKPEyLiZ5nTBUxl5KcCV5
qbIsgJFU0HlkpM8BcUwkzF1v95nYWGf8AGcU1xVcr2lz6BwoftpsazWdWcp/m6+MSMgiPYG2UKle
2ne98vSLaM8nKxToOsWejzu77uztixnpmNlMbQlTKOb8VvbCRNyMzsz4OI8BMr/J3NWOFM1KXx72
i4VQeoXs4FLElbm4TQJwX7xJuSv23fh7BkfwBuGt1NwWcjuC01vkAdgZ7J2DYO/Zr9Fkn62LVx5k
FjFmZdUmbZXxbKMQd/RgcZ/CmgiKWS/ZXAzAe3WLeAp0BWfR07IBZKFAzQXqgf2pewR9AVwUzgyL
PHR/lDmyjpRdVX/13ZQKSByI0fMaoLBAmiGe6l9lKz4BZNtnzwyPthLgCBj30qIFfRyhy2O/YKHS
GIs4RphO2Ul4UVT21UC+ZWluGJg8n7VqrbHYE+7REHAZBD22KxFlPkVrOx2epuKqb1nTWJ8AjpFs
Ryo9xOHpVVIShyomX1DYeHlq3yPUOcqITRnoSb9kEd/er5RB45fwzENE+AxFzWR96z7la5MI1s4o
bDI0z8Ad9u3OWYE9KNNK0IlYv8lotZEBC6QmSOuavuNSkk5rsIrsUhWiE32h+yhYf1rYwxveknf2
nyrHs9XR5WQWdqAm0bcDkaU15x6q330dyIbSbOKcUEQufRM06GLKAQ2UiDmuU+7KzxGOKQpRLoyG
3LC8eBTaEo/WNX/6vnlyEJxDXLCgUyTCJjzbw9R1WAHScYV6ObUGY0aGqsewUQU6KPiZ3AMofc9f
pSrAzCdnXpzhduYzNJF5cCY3q1dnIHsu2sAqnB3gnpPTxbrUDnNGja3h3z39WT74CDE+qFdG07Jz
iLpVKa8Xa9DmGYS+1pSY4S/VUbwHWr9Hce/lGX43FetqFxrLy5VgWLgNYj9ZqPPpfDrsbMZ6QSMa
wQIwDBtS89FFHmurFmxdZaCDEiHyxGW5cZq4U9ZgAJVOXwQZI6c9+nvt/gwxIbHsRICTwZrjxXRb
U3QdL7ftKslt2OB3PR+Xs2XLj1PWWY+E1V9HqIRI6seUYde2Wc5tw/rNhbPUHcxJDnooTLpyHLzg
/ogj5Q7Dm0Bag+Av4Pv7SuyDlhwlDerCwzbY63hEioRhxAucfznKEvOe9MtAasjiVUeBJNE9xDix
l4AdHhQzcUX7GwzFXf+9KFJgMRmHRCZ2ZdPHL/2IFuV0e8Z18eC90KrWUGG4jQow9+UZGvVqDfyh
Cwp3qqladMqUA6AhXUiP4unNS3aIOpZbj/duhGO4cvpCTZSLGuihGT7JJDapn7enIpC2SxJIUr3Z
HDFXs0uJENMYTjkNuNXV/116cUiLDQjrXeyS/neuDUtHZkeZvcjeCX0fj1nRQyscM163oGbF0Drz
jl94Hxz2zdy5WQhow7PFHJtOVa1zO8WERNrGlQBPRwvL15+qqH3fvEbCz0sJClVyn6IEHHkX3N25
nvUKBuQAK4R2HEVt14pqLrXbkiloRmIETt641cxANg1Krtg/WxnkM+ptIEfAznESJSY8ZEHdVEes
g1Z/RaONyFkcEdS68tu5GacMM7q0BR9JgJdRmVGM0M9CKCs0PyMLLXQt1r0mMxbdu6Z1l2zsz5Wk
uC7smTvUvV5qGI8UTYCDWxEKKxN0sjhxFRuEfMTZX1p12lEu7QMxKsWaU9l8prCT2buskoi+vLx+
TbMenm2qDKm22G3+JHeM6kjg3KI8wIcoM2yYB6YKVGJziNwezpFhU9kfM+/M4I8PwNgV8NK9V06B
fUZE/rz4nUm9vnvPDblQ4UM9gdnHcKNryIaXtASM39MvtHP+3Kj47GF7+tsYPonR2ewcfgI1LjxE
wYi4yuwLzHgYQnpVpWyq8H6vqXmrgqwRHmXsMp3/KLrg3sjw4Zf5LRJTWj3N8nZkXYfMidMfUJyV
Pyzsxmr7njMY/8BGFubmFYwUHpBbviK0Z0fp9rDe1jF8yasMttVH/cX6eEtWHeM3SyqbKBbNpcDs
xA1S0TOLdkDpoBpKNgv2sHyL4caXNumhg3ip7VAKsRg8ZLxPFRM8tz8GX+vQtqPQEgG5vTt6g82c
sPkWqZTRSiVOy2kfeevLPtkJspWlat7R17FdPYPUfMs1USD04dH6wDeRjTqRXnGNcS9hVLaPTvrL
izrbNfohq3P0hUsj4ZwSPMZdvxDwxpwuT9gi9xg2d+W2yjjnmGWsPfWIxTJrIYP5wlKdm6FL/Uij
795a/5qapIwTYJHlDmyVQEzczX5egGSCArhNnYIUHl2nTzpjcPFty+805jZDHKLa3buX3lditwfg
tqFLfNQum/g7GP8Bu+hgxOZ7L4BIcMumxZg9BQuoB3L/nzSZ82/gbett6hcMt6ZIhr2rRG1ywFwE
JwPO7eL/uwoRDZMuyxPpfISOYd/n1ThFJip9cC33XPdskYRuuo08CMSadmKr6NscQ31I3Ke+ccP3
Qs6zs0Yi9F6J+69s0Vtkyacayf+jxP0iC5aVtcpfwDkbZokE4MlykM4N3/JBCKIQEco9cAdKYk3r
CMQH+I/rXc8kEtfhLOIH7plQR4pXafNt/kS48b+Xg006nIKV2iKnhyc6PFU4yrS+K/ii/X4w1ULO
9zVb5VospUaplImMdIdQ/Ais4kacj5W+3H0YtBe1i+zc7WdyHr4XcPIyIkYC8g0Xd6xOt+AtxM6I
snKp82rBl5cL8V1PftrsEO8Sf/snKAnI+igQI5IvmLp31rbpyJzp0f2yXmtrtZlZoLOn/pZzwl6h
hWpZrYWITPuvZ5uQqq9C8sVO8kcyVpoYhAV1JquSVFtgkmRmyIgaCHBHojX6mY0DMh1heYEWiWqO
uaiu4K1/sn7h12EN2ptAqQrLVrEiZ/WYz1AGM1z7jgZ+oX79akZ5Ldp20R8QNph4Fod5Ee/7x+z0
x6UvOQ9bzN01/fPDqcM4N9qIVMAz1uBA1RXqIvUHJEmtCXYm3s/H07Hj1vW3/JBL1HNitcncMx4L
khymvsusK9PuiAyEGwobDo18GtxMnuOU4mvePGIqC6odm7dX98079TzZqOWintB8v+UEicrkccp6
zpRnho+4Ke0QNn6KadcUQyVKRmsoiZ715UgilGUFY3FQd+ku+VdInP3NHRDGO1jsr+wu8Phi4xHy
dsvQhNlDYzvhy8fadVia8Sx0WIStywJFyyNL6vJBzE1Uw5gAyk1edxSQVCCcrIJCORtkAe9s0v4g
IpyPoy73HAtalO+QlRiFKGO/BmZm57kQY72MQWWJXOcpJP60MRceHkM2VAM3heEbJ/p+uZhy8H9y
DHklpbr0SZIvRImyRfgg0rdc+BufqYZUIPT4F3c/nrggiAW5pUvWbpZgO1fuhMenRHNWcVyT8+XE
CcQ3uxNusBeCCLUtQOv3VT5KHcgi/GVr1OrrX7tH6ZSs5wwyrjWjKZG3buo88C4jDCsDJUShmqQs
H1BvfbihEpuZPOxgRdsV6qvcOU38yBuSdb9KDA+SBSAJvoEU37eCAU4GIDCUDLCHurYe2sahXis9
MAOa6xAmk6TSBZZybRL3R+ZNexwB5lqwx/Pr1EbrR/6OVoDfG8/qaiPAe2VUsGgxxkVnOGYwxb7N
PfWf2iEqyk6/4/7DHoeQPSkSYp0mRnDKAQJG+Ac7kWYDZb3HQn04ST2bg/M72LBw8k5uekiURECY
xlRzueMcwJotSkgis7kqoz8ta31CXeyLgqutO6Bj+Nlpk/o6vYnIIdGUiCAj/XKzYvWi1eQW3lyy
io++2cWD+IHc5PHJqoEnoE4W2EQ+izQmmN6y/8lvVQSXE1ft/PyxJnwxRuCnA7DExWHa/b80ZINQ
Fn9X54Azyhgrm1i1/kZXXpPHibnCiSfJgRevGs03YgBgQdJH2VdTFvjNfpK6/NwuHHhAh1h+uei8
OdTnwrqjhTyMzU1nkSGo4bUUCR/JRqrUIGUojQYRjUCpl7CoJgBcJguEMeNWkIBczc7ZfTmXgJ4b
cQkWgFiIRV2QlkUBnq/iztAHU7HvuUK+Ou/Q36jFs+6KNvGMNhQ1Ez3xHYbZGttscYlh/cbYJmHo
aupVxobJRPXzmu+93mOtpA0nlVnaHL/46dIux9AZUGut4G6R3/BRQU3xQlHr8cEJU9piTqKGRGS5
4zCwt7DnZZ5VvN7vbg1q6p+buMLQZ23TwmzSn4VDs+da+ddXnYf90TC2aOHszBSb53f7PkJSWVuk
VjKOCEaosYjgX4BzXLFiEANlqpMDoLeMlqY03akCJg5pUI1dyuFdYz3iAEN62AuZVEKXAK940sPE
Qobm02Mh8BKHsCF3AQKHKgwu5IZN2+OLjUyWODo1cLIM4dSJXpfaMtXp7TxSmQDEumGbr+tecW/c
IIR5nY2OOgIw+qPol0LFZZBssErDxM8/mVPRm3gsqNsfgutOSyVHKWGTnHrXS9oZkVQA8FaNhYKf
fN6L2R3HZndX9KCglFAw41sao4zBKs+APEUVFwyoJo+RhMCIivAlpEcmjoa+ObYJRofRIgv4aTnm
9STK3uX0OQDBRO14zxv68CuKWSmWampqMmydwxd3jjOflezommcP/INA1HBTvjldqrKtPnRVWnKA
h0PU8ji68o1hpRxN4POacUMW6XMvCfFOTfjS5M+8qdGEi81B8SwmVGzX/UF80+a/JRrVCILBPDbz
UE8kQlovXEyctTswfxf6GGo1/HEcCD7/+UWSuAKby4rmdRMY+eNNppIpT4lRTT0dh3qE+WftCU1f
yYH1oOVI+4k3UgzQrMMZrPm2BBS8Nx7iV6rrD1o6FRxl2+pJupGXejgAYJbIB7+lpzfLkQHrhZtb
+Wo8YjmZWz8zUWBPGLFLyyTNtRODFV9VDG2mLWEERvKvISFEoNofm1KdGTSVn+0CkAgeu2kLEoB6
M2W+p4zRsjpX529x/plBPC+otzA2hhWop2WuCXdtON64jKknTFUhdNGjUc/7M8jeW8lsRkHXdQ5n
5d6Us3CXp8oxGlKCvbruAVniSp0Eo8VKeuz8ZZuUemTtGG2VNesphNTtix8qmEMyArmOcYhEP+4t
j9Z7p4hIxoKzz+d+N84ie3ifybtgtWrTXkAA1CbUYW4bHL17xxzEe68EU+Qiu218dzhxp8rJR5sG
2X0lzxmo8obnTvi9ds6rr4DVu/i4UDg7RI+QsHCEpYPaHSaNSAvHDm7piIpSsSPako2Hqa1SOIAl
AeTKTh/rg440pQ2PZEB5fQ0NmK8Y0hBX/M5gYeP3uN2g7ss+GYTwPvuLxJovIPUdYmcOHhU1vfLi
2UWlZ/sQy9GZX1eLaqwaIlzH1jsEZtwbZZZAT9W9kfVNi46No3xIxocUTQZkAZ8wGgpbWLmYwg6Z
H0/H9SiByG5/yUhnQIDYAth2DMD8PQG2Bfz0k55rD6c20w1IzBC5SWcQn2Cq6L3ZuWvnRfNXbgq6
MmdaHplGi5YZ36AbVUN8rJ3Pb8aD3SZIAZe0OsQjQ1I7mf+r1ooP2G3VoiUxiJi7byh/HYtg3NC9
D1FKuGYZFL0wGUTCD5lNYSaeax2JtA9F6Zv0sy9y5WIk4OuiZmrOk/01iRyyAAAzjoWdtPf/Gzqo
jKKH6zd3fwcKYQmjrs9NoEGEfKmIAnNJxKuRCr6xEnV37poyQlQPg0H2zQ+Vlir8hVT99N/WrHj3
/VHVNOJwyCo1MlTlKcX6dXqR0mVsCBPX8a207j7IJ0Ms7mWm3ssQYCimII0UDy1g9iDnclgjT7Mp
oiZBt3Lb9Uf11eTH7m2svgZ03NRmJX/RkTEDpt3PbCIetQL+gW1h8lJ7yYxDU5S32H88c53R4Ftz
UnTDDb6AsgXSfWYxS99gLVK9tQL6+OOq9Ld36YRJVJmQAHyezf3rSWijOG0K70Qk3ypf+1MJAii9
Fu7NW4+XlMnkgM0H6fezJljF5L5qNXTUuG3f2ObLztNWP+e3AdcYuxaiBsy+aRQ9ryddfrN3c8am
N0Vq8yzSMgLuY3Rrf25HjQRSYFU1EbXppe19/z6ayVb1cA+jmtkb/lASwpVQF9fPd4r/Xt/oUA9Q
uiTtTXJDALLBzJR4/VJcJk1W6nMA9QQCqrWW0lwc/G1uB5srrKiQyHWWwSjARNPbiBOkQ06cEXTg
P+MI2n1HlZF7/Div4hfmnSCrLPRuhyssHFGpIcdAb7Ua55QmaWgbiW5Zns3VtX51pdiNzkyF7Ie3
1Y04raRB0evzj9RMR7Fz6ICYzEXrmiFBL5XUFgfbJwlQz9yqTrId1OpG5lLSN+BYXYNm0a9HP1Nq
noZFaO7XWD9yzSZV+lc8EoIAxLbfjv8xPvrIbB57AJP2NPF6GgJYLJIUlq20nIzw4O6K7MsGkqgr
sutITzuyqD7OdRc7nCQSqMU0Rk7wiS3szwRAftYYQxaU64FrB8j8NywQJVdrc0Q3OZq/AQ5BZa3k
fWZnh6ZTicRKg3/84htZTtqnlkkq4Kx0lsuPibtGrQGiEVX5enTpEosIBblxL8+nmLNiiYqp2C39
w3IsVoHNdUMqExBJOPYwRJK6ikr588CI+NxPqW3Vn2DWqsdjr+MDaqVw3HqjAstLxQHAwZWiwdn4
csw2aZjfZSGfneIdYUxsR3i+HjTLxaz7orLAbPr2lLoO/BKK86twCjpZIBhXg9IqUy07KQtQyCVh
2XtUvpaF7DY8IkpETl6gWpOpW9IlXcQsDP0OGZ+EiVzF7ZV3joeD4nm3xK2T1UWIX/4vBoZCSe6t
ULDK3cTpPcYHe6ETtGlDj+HmckKtk2bYlWGNYZSfWUc558f8NLdvfHCJb9RKwbtNjZPXTyxL2pEL
rI7bvJGluWxQeoe3TtdQnTpwWr+KQ7cecdq6sZwdbDpkZ/gfWE/LRoNN9exVSZTR0jGfaxrEckgA
StTDb50l3iHO8rDIBa2JDYpirVIwjmEQuO9hrawjnrj/ixlBS1LCEvstHsuUIfXv40g7wFXerRAs
VLAJYFmjLwRIH2Jrjysn4k3G0iZwTnTGMM+iiiC/qKQK0QCo4OeAoWN1oUObMNgTISqLZMkyUcMf
0a2d3kMUBzs1vduBSx4mDzUo0Zwm2aoGaugHmKwffawjRkm2yHiFk9BYZicfk+2eZDi/Ya3YuJsD
fZcEEGsGtGrch+TYhtecDOw5T2UcmctoQlL1h3u4/jz7RJkXpvIajYCIy1xohuAWIIQByku3yiYA
hVs9vWw2yEzJQ52YBDW6CY/UELb86qfObwhK8fIcbIMJ67P9SZ4pSoszRFX+K89lxON4eAb8PD5v
idBRJ8YRORnRiH331YGTdYYjShi9FLRNGDrBdwIxDx+gkRJSv8TIM7RhsYbjc9cmAPaX2DE0T+WX
3oWdzyRLE4Pq3+2N2AD7fRMF4HOjA1s9viqjnFw0H/cXcf2M+YJUtVm+Q+kTDt7SQkPX0uhTYKXT
5OfWBGFGO3RajYJ+P/oG6lXO6Bmp+BEF0FFo9Zgd/0tK5sdHjiO5RFtc6IzLzchhLOV24+0/+cLC
sgLYkOFjQlP7/gjxB9YWdW5RWUwZAqkVfCdPqO9CPVgiXroCbf3FwF82U9pos6c5+aC1iF5nSpyv
JJzuTmDt7bS+G3CoaI43GIxNEKi7sZ4A8n4XLKpTuvEXJIY0nVnATHAAEkPk+cEg9TvhiYr8/hS6
jrPUq6jBU1tVIydEjitlnApeyY9icL9XpaE7y9gfQNKLqdvhUixu7O5s7GZiRED5RrPSyv36+yNu
bzTXdvyPUcwqZ8bwGEgI+7isxCrdOYyrRycoFdeYv9N32/7Ska8UopmhyECxC9bYY106LQaG2Ubj
SRLROY+EFW85LRN6vlOOX/QMKSvHWIt4Iislh9HMSHz56j+QmKU/7aiX6ntUCzueWkVAUfVkXf0Z
z9SR4LNToNp6UOL052PMjgg+koKVrYiLgFbrlWC8ikQBVimySy6JU2FHI4BzQNblbqAtfr/FlWOJ
DoUct0Iho7lYByk00aKXjfMewDhxn5vc86uMVh73aA+qymnazh6tL4be/MxVxtbSWXVP05RGmbpy
5t3jxdxwIXU4nlpKXVwa5V+Za8qHJbpWmAgzOLU6LyOAdU5AkhqOkyD528reFQZha3DcAbez81N3
/gZvLpPNq3nStTUuBHPcHVPZuNU8jyG2Mso9jtPhrw/du2HbN3lc1M68tCdOXAN9/XF0mMUrzQ9d
QLnlmaaA23WBqFLOck11bZPzARHywh72bEef+3DB9LKL6jsv1tqmooAkceFN5IDtFhLrc2Ga703f
LZUkTFzHZW3f9NLBk7I0LCbkB/3vArrkESxHnM2Tev9AMeXb6fH6AZEaeuerC2FOjh0IPZTAr4ri
lJpbjGG4nNh1s0Zz9q4649+rhf9DxE0L2R+7xyJA6VwTlQWLmfMV2ssGPML0mwySgs8KeTwZ+RGK
zO84D7QO983nfVCT8WgcuOtcKvAunNAkpswJdiUIfos21irKGhXxwQEjlZ1R3kMxDETmmL+ltT7G
pi/v20owbVQcEczxPpMz9BP45m4KExA0WopaAJs3cYpbVLHC1bUsSbxRqZ+Mh8LE84OqzaWfEhVc
nVbx2euYTCAAbO65c/kjy/qC+iPwjyyw3foGP5Ij1XdCw+tdw4shW40czXJ+uO04jHuw8P/BVRH1
Y4Mox5LVNY97yagJGYa9hwoN+BRnjPtuHQo/BOlh9aJvUtrHUeIS1y6Zhyw/geSjNWSMh1huhBbS
K3PYz36HkWWPlU16ygyhCImMXWsQGisWh1zxGxPJxCT9+1aYvRFsnhla/Iub0KAPug2AuY1zoruQ
ysYsYEfeeYg10o7pJOtGYeamZJrvP+Y7ns9CF+zViKd7AitdhCtVVar6uMMtLpPjr6pY1taVu1jY
Jzs4y6VgS/f48dllcKcsQZ/XIe8PhDQ075PTOl/j2cNz9fNuWbxsLHOGUhGbZecetASoPHVbvNH7
YIbwppqNW9erAKH2YvTmUtTkhTKzcEx0oBB/Ggveu26Oxyl70zQtS3lWqEUjgH8CTjBGqoqpCZhi
orXa2AZimM6mw8AKUmt2LjLWQnaKKTHZbHebbLMvbqbRcwXL/4SKUNPmX6PHCgnzHTsdcm7Wwk5Y
82aiUJxAjCF7fsjj3gkkEhAUUYLkU17x99KBdM340nC0X0MZtBo2R9wqq1Of5kp+GMTVmCVbxgQg
zvLYin6Pxt0KRbISuuzc7Nz5IJi/XVcpvLovQouhT8Uae4aiESEm6aiE03K7vdBPBFhsdbxzT0ml
QL01/fbacfC1k4acF23sxLVgvtGO6e9yEybZjtyiYGxVG6ysgQjGD5EA7f9VrOOO/YmTkDh0l3CW
92/f1GIJ1Wu37lOAJ3ya0FUwVW8RqgfGMOs1mhsnkLdpuui9znTds+LsIdvb/662K5+eEdPxsOdR
P1UZfwotLQzkmGYHr0+dSYQD2xFwTRQhpkSwqq7P5i+bphwUUboO7Y9LnvRc7+qKPOU2Zry3L3je
o4GiCS6AK097f7N+07HiBhQBWLumGTArQCLRtAHmMQtQ7ucuWDPJKodlzFyh2kL8Df0d9mH+vxY+
C/WQkr+BGzPPHwvUmG+uW8AEyoBdd1C+k/oS0G2ovpfbedJvhZeDDmko9n9xEjUCDZqMJpgMH10i
X5sViD5+itSlxsLJxDYzzWcDPzFt8528XT8Ec4Hsot2YGYUVXnvillDFJiTVCO1GMkZvMHMWFqQ3
FGB+6NeT/ie0BsmFEbHnt6xsgRfemIK0HYdgRFMaGQ584d41cBvEgAQBrbCDkjKDNeZvlJc7GUvm
EzxPF0rtgOEQgOO/5xD5YYuqNZEImFDLpcD7HxEa8gCG/v20qHERf2uvsw/aCVhTK2Vx648wSwNV
TOQWSBaRBB86v2+rOP1p6pLLy/n9rsRVVvcZpoie+q/ju/gqmC6UBLBw2ytaRQrVzB7/n7X0lOSz
G9KH+JcuBh4/84XvuDOzQrMa0rtPJ1y317OUnDa17Ya8KZ2y44AUSlX8XjlOpXJ61oxQB/LyVMd7
87Zyc/j4KRAtlcBZRTH5ZKRqlNSVM956s6b8OOv872rmWnnpq0ErQ5iXr19wSqhj2xb21ZYel8SW
ihMUaS8mxU8JMvRbZOhspa856VfOYE1kzIOTCgONMX1JxUJgDVomMYDaDMgNJsMXKLXVbmCUwT1C
OxvRa9ESmEKx4Gqf68+/HVuSsRDP/cIWQheYYlAG2mxwWWS+hjpSGgB8SuqTH2ihJccSPI8cimcA
tb2hyfCQCq5tiqHtHPaST+i/Dypk0kh56xTcUSrAxnD0qPmeiK693eWaLzSf7NqPcNpmlZn+wWBG
deZqEE+M4jbJcm6vgpkFTfgwSDiUNqlCryOTzGy1zaGIgA3NJROdDTDLMMpqJJiweqoCqZcrzPWf
5qTp9RS2xB8gFKy5/Bl0NpRDlzFBz5oKbSUR/oq9OHn4u62cW/9ZtOJpT9sPV3k74FAVLobTaVor
2EMAX/ClSjUJh5XxAXMEjUBQopFmuS6QUhC+NIf4docCBGHbSJnzjmVoz3+ctUNXbbGux1fWoxXo
M7MtQrZnotxgZfFqyodtJ5ygvyBhqT+t9nooUfBZu1pg3F/iDYESDUmx+xWCuknCtNbR5gA5F8o6
SD4UsYsVmrjC/kacZMZs9dCIiWxBjHa5hHOG6zA1wgkze5l2VOqNeSYmacLhyKt6Boez+h55RH8d
YteVO0FHSGEyK8JKD0KkvY+b1sS1T8zWDNNusI4+JD92yzV4+NxqmoiShguShAP1KH8HhHmilf26
qSwkelaxk/qF5pC8qmRnGsZVdUm8moQBheye3raYKMcPPXhXw/bWJKd1CVYv7kakysr8CXNAOG74
IVxMETtfZ0JL+Jkf/6t+ibgvWrGKAw8Tx8I+6DPsx+8UES+M6tpFtbVdoWz/Fb7AiIF2p/xfr8KV
5JTb9V+xDGGUIVk+txQjI7Uq7/MjVa40MSdUdBxHpKLtlLYJbMpFSJFVff52DCHnpMyD6/3MGj+b
cpikj+zd2o9SMEFd8tzRa1KdEGf05PvljFWNuzYF2H8NXbt9jPyjY8nlwDBUxjiTzalktXQUeppT
QZVTdA+Mp9nf02C9q9zDjpCpL+OJHnvP793UYW7eWkR/O4LoYzwfyCQX0OGvxM1/USlIasV4QLF9
66QQcYRdupQ8SljseJlYYinpxdXGrwZwF6bo8s0+feGsAHl6bl6E+MimxSE8+NVHVwIz0hg1Wxox
RedsQpnlghscaC2j2uxSlon14J4wjCQi5VZmi71hXot3QD9n0RRhcqN+tJF/coxIcwDwr9CdOm9f
aywXqcYUkxUYIeWOrEPwnzTA1F4kRFwkZK8Uwscc1F/GMwCsQuSeIaQjIYafsiucojtv0MBUjI5A
zmrDdKtegpyT3metUgHpHo5Q1SPxHECcdiVN8bATqCQY1G7N+KOYthg8gnxPZUFFd30XBESeYsOG
xE9PVpqFnNqFrnUUz6X/6ynWHjtORyKgdG7d/4p1IrYldc0IZZDkbe+U0FiznoqVzRlXnAPyzqqw
OT50TeybKE/X6V+kGOVZtCO1t2yEQxSeVViklFdFtwhPjqNOOFioV82v59gqJjMm2b5RVgiqpOTC
s6PNSCTOjrEdc3XiewNDd2c7co7NbvuMRxfNFZMg/MLHVdH9wYELsk6dOer5sOKT058fBBWdnaGi
r58PkW1BeZ4VpwEpbDWub8uV7EJ/yAW6kNe1C8dXBW8/EGFpBKbBuHn6MZxJQ8/tdr/Ne++3MqIo
z7X1i0DqrrgM9yR3T7ib91w2K7uXNQBQD4Pw+nkbMni4rsFZrXT83i+zDOkV6sYQEfbyPSW7KvET
ZcLEX0ezr5M0jzANi+9D3cYgtXkq48RQ0F3tOD7EI3YzsYlQv0FoRHrPbDoLoTf1zHf3JbTiLDUd
5WmU2P7/Z2kk+d7TYlMf0w+3M6+SiAzcsK2pUWTc+5WVZUrAGQ60zt9Wj6lAgYgXko3f+Zd/OM+C
3y7k2w4if5nvsKp4gcYqhp6FuFBX4Q1feFfnrBe1U4oX+sONejEo+LRgxlIvFYAjpymij96ckOjH
CH4+cFwmX1seSdioLiZ/5hdQa+6Pla0OsEVlrjNuRxwD0d+rQCE/TcqPtVH6eKmUr73sYB8ZwaO0
GsyCaopvoF4ZrBgXCzF6RnhwLxlOlnD1jzxXQVpEHupFFca5xl3qZ5x5QpzudIjkdJ+30xfDky4C
fc8eg5Ebdvmey1w9oSN9azQiQN9YWDRcFvqUxj7rpUUo3wB81cIvNF9vrX/aNEoXHLKwbeFbPR5G
rFPQydkmUa6jb3fdlbqZ0T5Q6EhOZt5jSrny5RBdKWp5nuHkWsDXo6c57QbAwfK62qiyCGreG81T
igxxk7MzhnZEmD+bs0hHboDBsYtr07+LmsEA+vNnHTfAhFCQMlYUyQDCcyuU2pPL+eySUXildyPy
ymu9sFNlDKJElimiLbs7cEhGw6HdY5z97wEJE8HeY8L00DdzzoTVfBasjvrXglbOCuYnh3OxPyF2
AKPmXbBepNOhzhnmnqgifjUmHaRPDzzguOli1GQm2LwPBl6FXGw56C9QYdhtsMG4xDEgYOzhVUCR
jSXW7f5Zp8dxtWJnxiPn6PPdnvT4EozFXWsOhj3jPOvbb1VBLeemKud3/FatuSwTnR1l8OYSDAq6
TPWv8Nf3LDrRIzkJN2Z/uKvVPtjXeCdcZZLgT/5o9i+0t2U5ozlOrbbi2Fw3hwqkVjr+tvDROelJ
rX5kauaOP4XabY4t+vjMawx9a8xR2+WgRkRHrjBfvj949ROw44KlDDoxUjONmV+GvJLly18Q3R6x
lm6ACzm0mn1YFUf9b4d1S5AYUluDKgnFk21MXjnaGwF84PXRxQwtg+GlhKYAjxSoMZ6+PCn2Q3Nj
HEJBoE1NuH3LkrpuFNZO9ZC1k7ftwNOR1DrNqc1/dfvuuxl+7NCQlJD8nz6gDhq3v4oZsIomZ+nw
1UopqydEWylRo9KVJgb6Uvv+WfC64UJ0v/i7RpodJ2O5Uh9gnvmgKOVJrZdaNb/ECqbEQn4ap2YM
Xbtg1/7+m8I44zhXzpr3JrIdTsLVenLQhY6zqn7nLMJbIsCkeBBMErBzONeu8h0vo2+flXSUqETD
NR2ZY3cs1y29mRGTs3uI0vtaaSsjizqI1NZRMIgnCACO2zKW98QC/5Og9kI6ExrsOr5vrdFYYzpC
ciDiYsaZ2vG485PbWPPHetyvB6ymIaSZItUrGJmY8G9WvwesXjsKMz3LtbMted3G9jdhgen2YTb4
16r1gI2j5wBvZ/fuW3R6yiYg3E7uoTS63DeHj1sqO+kT40lMZ1yzZTrPChorllVvA8WSNBI0kYar
/kqImvaS+0fFPv/xyaM8fa2MB7EP/9bhXCiLn26b6rRW9kFYM3BnbgSrPL7WGlJBNfYdwcLyk6CR
1DozdwNlemWXVEGd3GYANfJ0gUeaX0Pd+cP2MosMffc87KzhRFBOfRs+pcLGpZla8JIyKhZX2DSd
vcBz8pagpjeSJjEReMap8YZmyuZbznHhWHFTpBuivRF74WIzNVfgKWa0kpn+C8L20B/Syh6CL6wt
WMr2k74/5IWFknj/kk6Gcc50rsCbwaHuUI5uEiFUkWhRU4JHLDZqy+Kqo/hYI6FcmsoHqwlZ3yev
uzj0mXtw5HCk9H1b40323Xr7VcFt5tCzMcBj81DEaoIlsSNjfAdzHpVJjfTB+IlxyrLNAvzhrosg
PuOcRooOHTkgrinIn6qRBndmkTk/sQi46HdrHyhvfffODyiGFKLy+l237Fdkik70cCLx5YHbEdL8
bgxk7YSAnGEa+89fbYWQ31uWhKwGrtRKuLfQSsVMZ5+w4bOl3zcs0jYOpuVLfi/o15Eu4gQD/nw7
dDnK0RnTWFBDr8CRzeKSAXvtndwQ/px0yxTBFrqrHZiSwgRLbb0StJRN8Iln32nyks1PMUdaYwIV
2OWL9C9cALgpZ09dwO8qk+yWrbgMm5wMjnh2NSJXW0QGD+Fe9H62pvqhbK2iuA9oQbY/5ZOcF2I3
tXy79kVns543ULwaXO/KQ4IsLHPBsMkni8BFWlDyttzUyllxmihta6CpVX71n+92KzZNd2YOFncs
cMoaDujN0b5iAu/YLGH97BQANfNCLS7UcbzN92f6mms3Yxzp76ORWb3+/9e/3NVmPjPfBuPhn7af
jSb4NGJ2D7P+4ep1nzJJeZjdO5HKYH+1ICHP+SuQCH1ALXIpgj4tD9GLq2wLtxONebI5lFcIR4GK
t5c9n0ZfO9yeh7NFhBpaXjPlFrnyIW/w3vAogZOGzqE0DQzp+RvSQrmrW0Q/U3keo2Wgp3hxbTYF
gbtLm41FUkg7jSoTrofqYgVrNMjTWqcsybtWeSULIs0Ddjwq9iJchWXGrVuUptmJFTlFVHKn97nQ
eFB43CnXAoN0wsarG+WEgqdHzQTmahIMh/udhD8QYGWXMqeaJIwVH2CuOG691zXcDKWa3WY5HouA
U/BvRM8WEXSQaW3CCVmtaO1fIA2CiuujsA4gPT4V4R39oI4oeM3icdDOY4c1TKmKZrfQuVyO5gXQ
rHw4oeEKt/5kFTdRE9tmD7xNWKi4Jg7ExcTeuc3+m1cW2wicte6SimAzP5rZIyohBFpAVFZE3cVP
WraTnck5fK9XREeMaJslS0sUjaKdvPUWgACfidgSgykTbOD7cYZ0HWp5X7QClAT2VgUUWc4wHqIC
T0peGYb09gZhd7fIOCeBvtHMc4LNCyRmU5WOfxV5DT7a5GAzqwRkRi39Qzc9LUtJ21KGsKFWgS/l
jCl55I8iWOm96VvX3zE0ySAUiILp4jkUWygljVYk/50XYGppz+PA546hzKmP6wfEHisosKeUX9Tv
WLRsMYexKA1MtSlOTF7ntY8mtiuHA3eY9CtHC6GOPWVQzdFILjNHKacvFBTvF+pDOsfE0O9RNigl
ixxfOjN5WttKHB66x5Qzy4k7XjhbyU598FjRDCPwYCrE+86PCIvWfJuVc9TO8yWwz+/WOaOMeXjH
tV6Ps/h4hw+2WGpX8ZOXy/26ErhdBeb07AAL1gHsMOsYtiQ7WB4KVw89/IPvTDwTSybIRUe5M2nR
sQ1gWtQPx+LQCgPW1c91NiDvFGUfr7/qB8dMYDA1WX9eNLvkT7qb01hL3oQeVhOM7AX09cEWcEPE
iZVLlayqvgVDAYK8yEusqy+4Mg72jzhrYgyKHFxhX2Ijwr7vyiP8gNF2311JTBYbioIznNwIO95V
273qgU5Q2u3ACm14B8ffJxe7prG9xZHEhbhILEZiFjEyxTchg9bbhV5blmGFDzNlcJNdTRPJCNDW
shtY6qRZSyqq7kDAGVijoet7TQXC5qk0Mi4sGTJrHj3towYjQgN2ib3fD08Kptu05PN1U9VMcdHb
idRu11EHIVE78MvebNrWlZC8idNQcxC2+K8nRLCnSwvsaTFqKzPqzTnbfZJGh9lzLXP8wLGNGYXj
QyMOIfhLN7N6X1C8IABhDt8CxnQFwTzBoQ9cvDeLJIHD5wJAjssd2+AaXE9xX6LQaiR/EwN3KCgs
FsaXBwpXc5EXGHnmUzkTsUrWYP+cZB/O5mIRGHccomaAN8UCBVvj5CxDirf1JILk1+ocebJN2BCt
IpHwFRuSi+QUtoaNY7rSa1MXquIxg/USXBVWJZqmfzqqbNWolyM/NufzLVX1sadBIHA66WFLD+Ie
jQl0wS0zj8j5qDlfdZj1m6KxNHJAZSKOWnNZiUsBqNAOLZtvNgii2p72+UeBMNAfaPDg3Lus9t83
Cg0wAfC8q1nSyQJJks9mVeqYvm/7MytSR4JwcHcLmjYK8xskz/8w0ztGeN6ivVABr5AS497ZaJM9
pKy1erxpzHPuPmz+gpultVN076kylBisMkAyq+sJ0DgtOmnVyxA28xxuQXtOFbHS/7VjepVZYUt3
zwxxbpKTPWO9rumpLUP50VvUn6cnDUg81vaTkZzXCccbpON0uPfTMyZOQqLqMBOyvigXY1B+hEOU
LoDRGm4QOdxjFDpRDEHRmzpJ8TES7gOdKjwFPX+BzSDFFGV8nasUxpOgVRqrk0NceY3YKfgjraXQ
3ovqVAwx7Vg+qzYuAGnG/3/EaG74bcNKikdWmXECToyCIaNO+BMdjq9sZAILxUrgkaLrGKr/Teqm
EB8xt+sZEZMm7vB/RijSTVA4REV4w5MhBGOj3MnqAYHlydntjUjlDJKyfd8f5JQz0tn++7pEJHEt
YwXQoG53MdCCTBuiH7rfp5bQvGZGDDr8Ez2ykCZg3RqVXDGA8TyF1o9Jxcai9lz+1faUX0GjKsU7
x1SmmBX6nir38CSdCLTpdq67hE0Rl6Cy5xxBkYdtqYibwuXxccaIpw5psPeFxEkZzlBihbUmUsAn
Jc8XNVW0YnQHUlIDj9KlktigB4hrvR0746Rwz7Wh0fnPIT3bSWML1whr5Mp9YHBBWXnA5hxe71pu
n2C9UinYQU94LhVTQFB4UMdPrm9Wm5Xvv5eoKX3UcZT+4rnBIxoAzCToy1DTigb2r5pfllw6D/jw
Mdb7k753CRTpXxn4ysXk7EK+O73ClY3b8HUvc6yMqB4Ub+M5FRFq6ND8EOwtIjTo10Gpqwd0MkJS
zo2uCcj/llX843ZiLNjy5SBxlSlyLeq+TZC+jlyP7t7Kou/mJMGC2F1aUFsjrSxaipyWi8ZSuJ3T
iHI+z3ncGY3kfxINkOUAqFIMBD34qG7MUmb0n6ZzGdYeITNqeCyG8tuc3qwSeh3UcoTFCnsHPjWd
hSQkHFMrfYy5hq6U/fbt0JifCNA054OHtFBgTKxxJ89moo32zaS+C084Fi5BXaCW84BvtPt9j/Ds
B3DosLGhOs58VELSt/Wldno8xY6IGtHXZ8c3QDibDDu/6HX2rqNSvqtwFBK4G2S3rkZebYnxl75C
KD5FAAdm7HWXNP8vrnPzodWh0sxd1vB0xLi26kinfrrHEhJdN+eurQjXDXUzAsz4fH2bWwkvk47m
MchK/c0zYzh3EGlaLO8nN/c1np20WF6/nzFfL/FFu1iM9fEt9POMI4ycIOoQCprLZfZQ0t2JRVek
CJxZFlfznyr1ouO8l8vbxfCEQzaEpVqXeodJGo9faG+fmZJ2qEvZM6EpMFEDapqo0M4CCdmV0U72
FjSerakHc4jeA06oEllvoovUFzSGbGvv9xKKung1aobR3+unOgFS5K81FRAc/HmMv1WUASW7UXdS
VTvOMSRTCXxuxXuX4l/Vjf8hgoGyIca3jnmhaPx7kiaYjAWJ5TjRhb9yLrL5JPRVtuWPKWbOCnH1
mWR8uMwmasXbvn2Ls+oKCR77cdw2E5MrnEkZ2K0Ztf9fI9FZJP1NRhl/X2aljRm9G71Ljz/+l4af
XEB8Gf/F7IQi7LLMl4r870RBEhVGWdQP4+zVP9uvlqPnJyyjE6Oh8ChLSKbZBv60Fq7tFT9I2SjE
83rg6mWFs+FXH8doXM9p+ocSdT2WsxUrUBNjkOzDtmijYPqQd1i23mKMo+Tsez99F35CGQrJVkRP
FP5VvZLztTT6V3Szs1Z8/J+5O1FeEYzvegNV+Z6iiCGt5wV/T+0pgiXYEthdYsZkeDua76ivpqsk
FUOT8o8uT1zf14AihI9E92d7V6qxghwKT0GcjioBY7OWvPqLW1pf6hfXdGDaisVOH5pMBMnNfx+s
9cLZSx6hhS/jOl7HWO2xouY4j7nsl0uVGzr2iYEs7Zcjc2iPotFJS17M6aAVg4kEFGZdUtWV+3II
P1UCPgaXArxJywAvSVSzGPTGH8x8mitNXjw3+jdVthREDscIVNIekHphwjdknpS/gmSDcpuRA/59
gxDQffMA0abHTSVBOUI547ZhocELwUhoMu487q2nUKh/HA2ZFjLbdu5C6yHydYSTQFV28jHy3p20
Lh+s8p/xDUZ+VxljEFShGhwFD9veGrcNkfSvGP7No9uMRThqJxrSbfjWvSN8aMNUZEwYnerVJrQ2
qNRb4Sbx/5GxSz450aXxdv6HV7W0vMK0hLoLnHStJ47d1m49YitRf9vUpB7BBLYyR1QpLCvKWos2
dbHPnQj0jXAGWjCm8w6o/W3eO1NVVPuCJFwwjTbZqmIE5QcZ6xk9lzOUMecxvIkmxnjjVpZDmUkt
bkZdDm7mU1H97LFqK2qZ2zBeyiRNpBEIGXihJzS3F+YvQDITm6vWbpXx1u7Hq8DuNb4G7gBaB/iQ
6Fn1yjVRAieh6+305Bpj5xJpREYKt/0srwa7upVDPqD2HHXYQtYTxKvr/n+qv7cTfwGCFfgVz/1G
iCUhUO0AjREMVLtVvkeqR1ZlnqYJXlJVAxhn1RN0H9QT2d/B63/S88816GRGWnmV7Q9Uwn0tI036
eusuf/stZ06SQdgxdys7h5IcUgB1kYA2oT0C6eajI+Oj8piB/wnDoXC4GqUxecCYO4VD1kl1fuNZ
aqeg8KEVqFOllMj20oe7yIhOeopEa3TNhdonPYUddGsGtMb7SopiV22jmjJsBtJGsid9cDPTcvZm
Ad6Mzcl0FrodNYwjiuk9lMPRu3AyMcR/5tAFkLXBpUeAMth96np7zAvsUN3Dd2P2MhfvwXNiD+/v
7nswz9bA98pwADvm2ZW2qxpGQ21gvMGNLJppv3lyRBd7WA1Q99lbdVuhzUe2HxmV/mPIKru+wIRN
fqtHEBHF1jw7yhbOD9KefHXB64dqp12DrxO+gUmJAW4gfoAXzPa0lltraXLYVwO0YrW6l3VFkWoY
CDTKniDR9LMRNW0pcdydVCkMHNcR46V3b2DFVpFHt4DDLywYe79Y16jQ1/aK4QNseGzkv1nwvew1
q0Uqna1SDOUvdpThbdfVEJ2h6BQCHJt6TTSMHusKBDnFwICNoMRD+TUroduLK4gTZGEOyYxDvtOp
jIC/lTE94vy7jKyX9surmbKBzAYvjJeP+0U5VYuNzy/FOejf99bnBCKH6e+qqGewPieJBToLaO7L
rEzTBOaL3xNfyeb5NQXpY91+ODwdcKmubcAdV6+ceIvSK7p4JMscVA4m9NeWHaZaJ9b2ZZDSpkNm
+785hBy9kQv/C3wPQIWAYW3abfp4FTksZVBuuZySrUv1NRuan3fUpjHzgeT1cMUpf9KKUBbM+GT+
RE0CAihLGX/DXt0TGPnIaTw46E3bnCg/GPjjoIsKhKsUCdp1dFl4tCJ43bg8HyspzZwXKm/ZBSuR
m8lpbHp7eSxLrHVaXaoTPyFScHUX2CRGWwjGvaH7NCQ5RwxVg1iR172q2CPy7OJ2rpq2g3coRusy
MInZU7S9gBKWR7iNF1M/PosCj/zF+ESAt9f+hTMFEkt8yrxqMbNeHWwDgDJ5KVjFLlXKgJX0IEoA
QupHUntqtlLzmg634lvcolLisGU4quiPSDFkpMQfoSkslDDXVIDcaST7W2W/2SzGQCRIZzwNo65G
JtS2/B2qqhSZPtAet/sqa/jmuWMS0Vk/cYQx6VDOlfLzmS3Iy3GVXc05mi5tKDt1p3pk3G0sfenG
sOxWKJIXnnF/K7RxJSHkUiZjcyoA2YTu5UOl5JrHwKi9Q9YuK/BYtnGgqSS84aPtNSb1Ef5N9wh3
2nAWZHfoKZVnD3FHuPfgLRaJ47w0u5cOADD68GvdurQTobepC5aR1AB12qXzkjaAMHNA2ozvdXXb
QWRsXGqG6NWN6KuVIyWGBl1iT/nH51npDRArhve6NaK7vkoD9BFWr/YFRKVb2yGpUPRpFBfeasXs
dhJ+o/xm6p2Mk48gxW7nTnvMS8Uo+HRuz/HngAfA8PbhQEAtHnPHtkLLD5Vthi7MJNpARIR/c+aE
cXg/XSLD313DX6ny5KzbBDmz437Yml3GR6U4LgSCrORBR6BmKfJeDBpbd5ct0F2lUbxsDCAIDSj2
K5JtCI5LK4HqGigrnwSTwi2Lis9ynQF51HBoBGIfQwXn4PwIjiyl5sClePXjOp8PD2YZVPOhfUmi
qpjcdrCpB8337ToZTdMBlgloyQ2+LCvKxhnwKfx/veyOZ0heS6kpYQrVPJU0drklgBaCfx2pw78o
E3oToe+IBYXWt9rUqzopUPcAO5pK9ckrnJ9Y8/P6DMMV6cojOGRaMl6wJS6zBZH8RwTVsuUjQo5y
FZNbDk8Mq5MPJXr7/bjHFiST/TL5oT3yzXgk8DTVjEpZdOEUSEggdr0Z178grHU5PmQRhU9iDB1G
bAGrzROnCBT8j3h2NRgSpAkP7MmcMGMl0DGn7F36auThXG8+3ELmFFEJjztDHRYaRyL8cXF1UJFH
4f533hRFpU9YOw9bqxjuZvkgi6khgWy4sBizCItEFkFMdMO3Ukum1f5yj365wCvqZWgx+Z5gGgxn
tpeUaEPQxCFgP1VC1wLHNnskCNANdIfi2tb58ixlmhjLiB+ASq6ExoSurfkl3/Ak8ahF9xy1WXhA
O4Mz29gEtJfL0Tv9bs8vQJxNTq5bjpyKwSZKn/9mT9YFPWZFs/UbhLeI1bf9hiMNVAm/eoKGeQeK
nDqWwN7KWO3Iw1DxcbakUSfcMNFsVotTJmbvO9rWB17E3YiVUNzjk7VPdCzAu7prbnkUiQh6oJ4f
9W56YHe03dKkZgeIz2Droup7Op4dxyHbGzLqvOHVQwgPHs/su7Z+Y4XOe7+4AQ+aQpW5XFNMNG8b
w3xuRXYjWQakhgmgo2ErZFL0pnpterA51mJuuroi+FxXbT8VpEzX4FCXb7F/MydxKRpTGmimjmSc
PoQ/OHVBj0mOxoDaz2rSh4If4zxGyux2pevuuFjfwp1yavtQieqgpaBISKe43/WoQ/E4yizH1O/p
CpWJgl1AKSeknlVZiX7oeDkjaaDmkc1T6sfzhGccynqKlo2jtC7jk2LDDbyVJeUQ1qbfRg75LNgN
ZjTtV4yemD4dNYpNxmI7tKBwjbgiNz7/X1nauiyAEWNu3pEO1k2YukbRqsh8zPQtkvtUWrcyHXcc
E0KrQSBE0FyAhltjxr5dZuf0V6P4WqLEzL8lD8R+ozY+Ipt4tt6pnUmEPjyNWfo8Ll8FbIkyrfRQ
wvLxWhcY1I+lT2Jw6BuQmTSiwIjFQEZBixzaxO8m/mEwc4Twx1HxaJgoGCOdiDqanQUNvNWdlCfX
A0zIL0UgX9U8bGT4HvRenbyAiuyHtbuWtwfof6gW2yLiq0lm0g8UvxjEQkQJJKYFN+SgwytwqScA
rVoAzZJL4b9lB3146jKAVZ4IddAWNLrInMA3K2FGMLBg6zW499jrhJVNel4BxP5V0b6zV7R4de6q
LFPLEOvfOCUF5qyodGfDb9Az3uD+SMiY+cC8ocIAQ/prHa1o+K0vGGwwMaj2ZXcJLvsNtFdSuYW/
/Jj4nrXENANE8EZOdZJDv/I8zHuOLOUhxYd/wd7ZxQg+Q+KWYZMq+q2imfs2wkJjKwtg7sQuhCnb
YPC4BGGoCsPhw5LHBeaYubOsXSQH+NG0OyuI73r1kv16++Lwgmmlaprng5zbPUhzCnW0BV0B6yvT
QWJaDfgqyAzbo8iufMEZKUUbrWfZp8tLFu96Yh+2mbmFRwd6upWZjUUT4FcxUCWH8laD8Ex1Nn4s
OJVB4BA0e3lxYHH5kSIc0Q9kL+lnp4LPkjs/xcvWTC3eUux/PlYRNaq3FvsmNYZa/NLdoL/YmHnu
ffHu+6HmqwJHH1tUjkIWwTKzoqFkXohX3/vpO/ZkUpM/mOIn3x8q1utcS0Bw10aEA6v3HHqeQ/ye
jTsIA7D5+cNbvIF5Hae/mwItokmZnzXdne9vvJQSYb7khtNaxcoNainSHhth/yIgRX6n4O6fz68U
6JKqxt5dLOFrIMFfwYZzK068xxDp8exsyoOhNGNtQ9fDti3/d1Co6AuomAIflsSSHKaGoUqLeF4s
xtziTLovooz3hhMQ27ckUmLhn6CY4OH4a9vPAj3xRWdOzM7U7labWfXLcSs8EE48I6Ky1tun78yh
G75y00mIhHFXx5lYJ6spEXy2+Z3e00clvn3kJSaD7IdLM4Va60k62tgIYrp9bluR2dbC0zmQvZG+
ZEe1mist/VMgr8lSOVygnAAAEbA0PMYPFLvIocIQYZaH5eOx+laIkIB074rqwpjJkcH6AHvNe3s1
i/nYFsRzvZym1lqaI9IgfGSdG1CoLTFYOV9yZavOawlcu/I50u/76nL7Do+BwEnfkzzqUxBPrTu3
bj0IUoIMOPtqe4MFcs67/oWqBsUl5QXUrMGR5wa/r7d42AQHzt7fCv59XuzD5PZTBgPBcZmWrQnm
hACOktl4aimF4DnRaJtXxdfsb0x2V1KWyFaglnAZ4CzMboU8wKnUZ9FdLNiDoAcD2rBUd53aR6fJ
rDcUjiDSe9U+0yT69IYtT/fCgi3ehCoEB3rHyHdpKHriFx3Q/V+5g3Qv5+auDs9FJ+1ExoBZ7IuN
uwmKxF+Lr8iPdVrM2YL4Go2qoWaMVhT66FYWEkyzOxrmL2Y9XKk1hPNfnAc4LrYhN+gKd9P/LHCN
8vqDQ/REHV/zc9JIGtZcGw6q6heGCVApb83DsjW94bmfciKefV9I1V8po/pv57SSOFkesWFckWg8
hRnHHHELXlKhbZqlmQsS6fCDwYXL3jluZPPx7kB0LQI4ZkBRI8K32ht8U6wGkIeZNFKDSTNNluUC
xG1IVwD6MJHJHWI6E33nOWqaPUxO/0zq0k/P+GJuDChorC37KSJi+qR1WsntM+TGtyG+p7UY4sNY
nWyA810d597mTJCaO8gaMvNWOBGZqBgBPy3hcAeQelNdhUOA/5Jg5axPN3ft9s128w+s4vh4xTtd
3afm+RIJxrWdKJVGDVK1JHdAr9wszRi8RiuymOIIbpmgSwrBSPsfHqtfuOegh4TvlXvRryesh16I
X5mWEgE2jmjpcid5dAvvHwqI8/Sy2Ml+cQl8el/y3VVzDCNm5YPLT+ifsCyrP1ckfHE7qzNqVN+V
gUi4Dun3PGuWGJ63Wn5xrKOz+2kw+Li8+ojl2MkzMSZzbFNI/ktXAKo1d+E4OhaPduQfXiBRivA8
LiUUxUWlv4TpIvoEWs7JgL6s/AlwLXxWa8Qug02fU2m3zWt48DJwUUm9fodvXXLWhBSfYubMRta4
j6XoRksK6OnpgbTKiTnqB1FDWQR+BMP5AzGPOXP+6OSTD/wZCrPMU/nLIznE8qnwb/V6p6ywtqK8
U/Vf+g5viRW+JwSJUJdl8DU1+tCIF5MQFFbFagrvdxyxj5N27m/NSYZyQ3b+uofzcGQ0w85licIg
fBkfshzB53URD9upokx3mfyW4y13qBxJ/HrD0mt8Y8THd2k1f2c7hcQOuojcVwoBmtf+szTSVzpZ
vYwftOX7zwSJOlRMAzI5JeAAg7CqDPsT7A27BKN7ocr+Y3g+tw9/n7DS4rfY0rRWd0umUiQErwGq
ogo9fhcrBK7rk1uTDZdQYxm9iuV1zqcR+pKnqdBzbtpZYP2839i/ku47/SrREd6Wz3wWLHCllLxs
89h/wmQpdW3eYExG2snKwm1EJHkCrFgkNhwj/CKC/oqieKXZjKfW9JImYv3pvkCGp00a1qN+PwN6
4XWD92YMzpKJSeH8+aZYejPRQYs31dXWDq/w31cbGZGTOnvumEV5amfVpwuM75bTIuF60voqy5Zv
ALxmPF+vmtciI62Br4Fy6DmOeYwhOmYb9osghLmiQxHXhcpo6KJryoPT68fyWlUdF3H/Y9cEh0fl
gEgKIlEmYJqyV3D6i2to3TTultnD5CssYV2pcpq54fKoK0nHRXp+Z9xXDD9uyDfUwQyryznKh3Wn
wz+6d2gMxoSurC3y7wUAg3njx3E0OtRfDQxiOOgoHCmW/UsNLO+R9X5TNyABxIfn+O/Jfvcw2Yjt
+DSNOtxm6EbuhbVgTy3c49rB/bUoX4BBPN+jIexqqhpm+PBdfWyqbNbO2JyznhB02Y6woCfRLMQv
AzhggUE2kvwyE9uDlFu+K7rqRk8uz3NaxILE90l5Y/lsiUQ/ea9qRVydXDkcEV7/dlw2YvADlGTu
zI/U6EulmOAkmEP636VH+6jiK8QtCEM/aPlJGIU61aPehSWu7u3fuSdeN8y8p9tS/WWWSsnN3L9o
mwOE8FRGdLKcXrSuqXlMRx0XYiQw53Fdd972AUdo1+NjKeoMTnTCWV2CwXxcw51VpxQkux3Zr6eI
mVplM81pn4pVBhlDZKfmemKyvWwsj16xQfUYnAS4fIL/gPH99j7mLpLAvNqdEZaf8cdIrqxUMSSx
LDDtd7vb6Ut5EQctu6KuNLz+S90UVstE8XeWUdWPhYVrK6cP6cxlgBL32N9iHFcXiZueo1vg8pAi
L1X+zwApYH/+d89pH96rGCKhHwDntVOhHDmyVJSzjOfKnMVMd0XzBOyosquFcEc2HhMvkiBQ3W9c
TfyAvzG47pdxAjCRuup6zbIHt7nLx74LLCyV1fBODRWko76Nx5I32XG+0QeZRK812lcJwo7OhfgA
seIjs8uEK3WqED8r1RltNzk3xaYdNkN0ehUl82P0HiGuREBmT/1n14moDXUmtDRWUuziWk1OsYjL
zp1GpPzU264bJXo7plPc3ljAPw2JeEab8W2U/h0INQR0tTlqTQtcqrfYJ4+UFqb3Z/9KKZVF0WBF
34C0uJbXMqSWjNj8NPu4sqXrqSjSQO07IIKgUCX6Pgdn7BHp08/zxbJteApgJQ6kE/k+mek2Ui9g
rTHDO2wso8b+TRjxzCJx0blxxKvUsOKAcNaBESAwR3/mm1+9H0EuN+maiV3Ob/LSWOLiZaH1LvCB
SBVo1ZwJT2ZC9bU5gdPetzc9tmyXWoFdLfRd9tU8BcOKbgNO94AREifUYZ9JTZoSQ6plzzvjYqtd
jWMcI9+9LPMZ4aHbAwXuUvJOd8Uc0UOOGMukoHwxVr/l8WNrVyk4eL+MIlxn1+wS+4S9bTmhifJr
MKDwnDXOgkJoSu3gq/0KTyybDslvmb3GZbgpqBIiZiEHOjn8d53Q2kFyHIGNdedO9vi2mD1YWDGf
fLPb3tmIPiKlNccTICylv+NKrBStV8FWxd6+Ec2j6yp6QmcpaQ3XOIujob6uFBAf75Gd0ExswseQ
C6+WhAjgTwN6D4FowUDddQsju3u7eNWISN014KB33lBfhy0IHTL32Q5omrAYG0xSzcT3EADQqHE+
CvJlgYVvK37ngekvyTFNXNQplfQwRB/o4WJNn06JCfVKDGLDZG77RgMzalVfuoHo7213rqkDLjcD
nWABW0+8IqKR5B9CzwqoP/eBmK6lFAlqFRxadDqyiNxH5KW578jK7QOYWPDMRVklk+FsQ46ZzYIa
hCKow1wt+L6QHa01tIOZmqnwSpfqMLWadKdatgipbTMdRlUBE5ipg4SWMY+oHmhazgP4nP8tHm6g
d15SS0/MCG6FMEaZ8wof+CqYeDIgqEaWDT/YLgqoq1ndDEXqnVGAzm1tktyf+HVWts3Bgtk9dpGi
wabHXG6JceYsNL85NKx3WLJipa/z4tMkC2t+H3UaS58OzAmntVXIY1o/xOcMgLun1AvBCQriTCXJ
LtR7pgdQyGKyPiJF3eu5vFA/QggTRiR5JV3dGRrP/a6LdXTHJVyKIg4eiIXm3l3vM3uuvZboOGpj
mJ6KC9UcH+MghWRohDXHj1F0GCxu8jR0LpHrUh+5hzxlsdkBUD+jgBjFHCc/YJgi4t1z5pd8k1/u
7+AOSDKR1X1tLUg8GQ4OyQvcd1IoivtZffv+8p7NMwhHqETO6XeFgoz+HhyuqOrymfdJpddCNTQA
cZlW60HMRYF6V1woARHLdiom3Nqj+srnRzh8QxRAA+j+UWm3rr+ykaumOHNyF2G6ZlRniioIgSmk
WaP/Dcv3egthoZ/zwmm4rQSyHbWSLx8TMpBs3FsspWKdK7xQYVZzkhPk5woZf/OveMXEUE3KnjEi
0KgfVK+csWWDHa/mOlEn0zWwbHmjWUxb6jrLmC2PS52Vo0W9IZMya2S51FJJ/VsU7Ba9jmrEfg1t
zfm9TLkdlDznRaIwrtAqg/+XZrJPFkCVRbyTnWe0AnWRYz/BTTRncUwlvzI5m84qDOZNnu7lkM4O
8uvxULoGNFxxmb1TLjXcECS1qzur8ocSU0w2phktNCry/OSwOljuWM9g+SZ3Yx5SyyBnktMaSJlD
QNVPYrfMuIsxKtPlc3wc6+QvPywUJmmY3FhYfhcbhQF8WNfZ4rWm4VrTDqS9IuWNAqio5pHwWMH9
Bi3LWGKebmYBXlamcVL6L5oAQKa3wPdtiS3lLBsMkkNPFYsyC/LsMl3c1cPnpSbhi6b4r91rCSnM
Ir2gMbzMWjeSwQl0ZpupGEsPT5UwH+NIoSJMYWumtUBMs1yJVR7WMBtZl/k87ZRJs4oj0nHz7K+x
ys01oQzfPItWHwERej67N0XkrnjFBQkkUtvAZg0SZtfMzKaZNaWI8BUhlRx3UiQxu8uuMKd5q39r
dvWEdWd/WiHo/CxNewQcZSz36ViuPnAo0DfeW3c2PwGdqB2PKLfEdoClOFDZ3WSu7VHWPD74149j
H46Tk4pWGlfJZu35fuQ9pPaUU6FHl+6krieExttxkPLinugisXmXqDhkQAy9z7kHcRaOgehWI/QZ
oLkEsecXo9srPTmcX25L0L1XeHQaIRE4Wg+2+4WbsV4kysjmH8oLvLxwoPFDSnMAwvPwjEEfHkzB
nlum2eYtd6abUMWB6frm7Ozjm+qBY12Tv8oE7EHcmFX41/eOAHd5QW5v+bucqi7IEVIivkEwaCmq
cA/58Sv/DUIKerJhCyUGNaswWsV49hrF7N7WoV3P1wGrEYhC+xtR21n5gEeKVDvZuk5LhIkOrOeL
velXEWIIekGBV4YKyMLJWciMOxH+Wds5N4qCICbKdHK5C3kZoZGRK8LeFHisi9eFskSiwkVj2is5
VEvL0LTB0uGXaQeempN2ETDUQAtYroSt+2bEXgB13BKr+lTons7Uihu1lPATfl+wW+Z+D1g6rcYk
b0THMcSiO+AXxVR52vYC6ZwScLNZA7GN5/DMIw8GYj4XE5s/0zzVQ+BLjx3Pyh0woJGyTJhCdozx
/+3FNLYvjDOHX38KTrJXsbhC5y+4/qdvnAFZibPjHPUaCTHX8yigzNbDfDxjlxRh5YKR0af+iXWD
Ry6D0V7jaYdlaMxMSG47+M3fHifQTm7wPoqbuRV4BMyejoytmzLq+bdscqzq4JwaK++NBXuVuJ/g
hhtNvsy0GFGQJCsM2pM0MapLFKX9rpc7vC3gutJCEcSL9QUy3RIFFJH/kcce83iOI0JtOXwXz4qz
hu0Q30/5VDrnNuC300Vb3SvsxC5FVkmi5pb6Blo7Ea9gGNuwwAobYoGfaQ81MsGh3rLIwGsxF9ms
fxj4W3a0gf4W2wYa9jbySnUM40qBFKuJwqyhx41UilRGL5eIUNQqS2yNZ9xG9iyVah3TzOwiB7FP
xZw4/BfD7pQ9D6pMbr021jABrtFrCLO3OQFZ4qqvgBSfdpgLA/HZro3a3chp8idDckDL3YKgCd8b
rkQKPZw7aqOpT/dZapgqUg7BQbkW39AMjED73fUVU+0VpgjiXz40qn+kh0K1N+mwe8HRmNEzVG5l
xgIbpm7vgz8BwBM5sNSCIVoztSS1NtldE+0tWMwhrd7sso/z5Z8f4F23cijMScMlxmVDDdG+1kO6
hBS24+BMgwRDXe0Fejtke+v7wKIIzIVIMyKmgLTeHrmjvYXwlPvlPB9URWfAPoCQIexMi+Si73CO
94wJ4IzxyBafIql9oCkGgXBn+RZ3Zt1KWXDL4grfwljWyQEm2QZyTEXTuu6Av3TB9mCFxZUD3xj5
teo5Hspdb+aIgTLEEZxrGP9IQR/ANCDj1G3yDbzbDKpCwFw2KA1IlTM2bC0Zcacqlf+sJr8+Y1lA
iFWQOaz4+yr+gmttVaIda+vnL7uZIdWdj85xb6cthrOaMcRJZ+ii3z7+ysJN0gp1FsFOYCI02wR2
zOpLIyXMbSm+sLeqNoGOZ/wjDeYH0nWY7HlDFSw9ovgvbDP/WXa3Z7G9KphtvhzSxOty7clpuu0f
cOiZye2vu5qCibD4anatAsG6EeSV0mLaHuOe0BYW25fb6n3teR2fD6MOXkpebz4/Thc+yW5twWdx
6s4DFebDSDNWWh89hH3hzuKvtyzkTUSlTStDE7FsPUBqZO3GaAHLN0yZYAMfGD8J3muv05kG/jtU
6YX3PQCYDjKVWXsqujCylu/U8bFbhrfMw14/4dpOwQuNZaFYLavsByCVVpgtcyUXVS9PkbCxj28H
4O3dLlBmXSEkdu4h+W4LuZPWDbWWUw1YCH9fG5vFFvkQPk8wX6rw5Xc1G1Atz4LZ6fmvOAkww5XX
/6v3sFiK1NGNocmC6s9jLXUEQla4a1YaMcfJy3zCEqzeTg1V6WcIJLE4A95A+5x9wG6Fv1xvYKfP
pv6tLQ8HzFqdFT7nQ+tx6tKZ8achMTcVAOYEZaWG2IWv+fJVV21gFBKhvm8lySSbaJDxTs2GGGju
L49BouCv8GenJFdn01Q+t6XOcrssIguUyHq4QiEb0QooxWGllBLjiLzsbmamUTw7OFXPl8uyP/uk
Yo2V8ESI310p09VPqXRyTY5zOv+cdLOCl5ZtZRpZjXiW4mroomSZhwTCFOlU3Ve9lci1Lik56jKk
fb0W1/4iUKtqKFF7q3mXcDdFi7KfyOSq+S50sXc+jiYMFn2C3CTbSyzDapmk7dgTaGGiY0SHFfuf
oVxvGCB/L5jbgcTVjIPQ6afWeLN11KPEMtSf4N1rvccOT5MenetxVRXuRad/WFI0UnN/ZMNx9Vs4
mhRXW7MzhUNRbW/OYJxo3cSYoopQIBOT3EH4vjdnbTUpGQx/GaNxlybdzP8cM8cmnvEs+OOqgWbk
wzXUhOSgjKBxxCwk+/v6Skfolg3O5eztO3S+7itfl+iVkk5CfjAOar5OnM9JIr9CTkF99ipKXInq
qvDyM5h+wlKJ2trYre4KO+W/YtTxi5UIUpJGE+a+QK63nlxKJEqLM4UGTEKSJ0Xk8tcyJnP16SA4
XkY52gIbfBJBq8HWZmmEddtdzQdnmxmPDTQlRYgG/r1hHsmLulLOJWlT4BsVDyd+JXscJltuwim2
J6tt2ienKzFewBzQ6yP9jBE5HOysfIFd9X6g792KT6ZGFB07Rx+/8xVxzlePzQENDGz5gOZrgc3v
iGbKklwYzyznXIn7TKWJBVU94ryDdpePLMuQEDecoHTD2fWI2M9n9yz9GmeG6ACNP19qMmLLQhqN
qXl03o1eby9YPrIrreJMBH4RYJsd+RjsnvxzmikRxTkYR5/+MzjCflz0weyvHLRzDbkUBpKBWapa
sGUqIeexU7XmqLkULGifU1qTiME1sISkof6QmwzucLzOzT4pIGamEz/RfTPnCe0sPtunZQDodtDT
hGkW/+y/mzjuv8deecbeSGzgBw75EkmDJR/w2MHcxnBHzfi03Q2CqGQ705fvsYm+8LK2uby5qswP
vE6xZJab0G5cetyduIEFIZnlZjDfk/rSRhYFT3F3aP3pFJQxFISmLf2q+fC6UPpvEgolZDMVblHb
dmmSBz75FiMVrCdrudWxwHWSGF6LADFZvn7SJfqOgBCk3dZwcnB07cSrlNsCc9se6nbwAGbnjcV1
GiX2Nv8684O5C8ajuFQRGir2SyfEIv8msSsSWRHCrTf1itC4PrlVxZ3vB4O9k+XwexDdPr2V5/Bm
MAMOCqR3K4AcJ/2bldk52enI2lc59K75w6xsipqWdhagReWkcOaEluGhp5HTT5XQqJm9QFYnDfsX
ocO0EnI/NyzJkHnKJ1mgN4ZabFG2NSVxEwHTQHprJOFXyK14NM43BYlgUEZcZ3ElrdJrrrmkquCx
0rvAUwLYbKyeD9yx8Mb5FY7YO/093UQ1vm1jkn4Gqr0rKRIJzUqGLwKuSuesh3V6XH6y79pngxD6
OXaMcf1YHKwddL7icJEsRi61A05c4UBastB7gtfGncloimp5r+VwLcn4NV0le1VrzmqPh6eUzvoA
GbSXDIbocdwqpb6Cby5O3QtWGXDkPYFlXFWSExEDIDAwhmfLq9xoc+R7tmQELlYwK0hBkge0UyZJ
TlWyItzd9aXqjcWMv2W/kIJKezxHFeahimZ9fFEBQTaX3IqwiQA6+0h6Yo5ObGLt75VGPZZPwywp
yYoHDegTQd0L/clvczrtYmOs9QDEEhOlu81y67+aVeea1QmF2TSXZ5FtHjS4oHxhiJ7QzziZLN6B
sGSQwnA9o1bV0w/Uq35mRjFQ/18tmNwnAZ5L/8LCRNH6BTt0DgEriZbRQBaP9xlClKpPFgo9VqLB
+968N4xE4iSp9AvPwjNCSrLg5MhYMcKulFmArnyp193gjceJfUbFfQkyvs9vGVwA9uzzZ/h6vL2N
/Uh2NuXU6G1XzeqlmykoJXGRpskXIy+iLfY2K9Vl68FWNN31ibPwlwIQ8rNahzbJDaF/WsrQ9jr6
aDIbVrS1JhKjTXVLATXGCl36q9ZaKJTusGi2e6kStqk8rfqj1xLilENi2EY96YTPnUUwYqhAOqvH
77AJFfSsgcCkoDdG1ft6GCCHw2fKkcK4MUYnb/Z7WJwPDDUmNLxjaZfm0UXk/moFqMWwc9w9nPAX
6HpOxvxqi5m5dcYihLEiiJvLnWLda0Jd1KnD+6dzedTLksKiYpLySO8Xb0tiLC/vTZ8E00lPql9O
c9YeuGd6MsrqMxXbA2A8ophFbURcY8XwNkYukUEmSPho9pt7qarZU5jJWZL0Q9HIJTb39saPSXIk
lmbuUftu7tofBBX98grBCV79XYQb+YO4yYGsAoZ5TY5X7lYnHwHKqgvOR5cezyX0a98F+Vj8zgo4
m3wVPD8mA3rLDq7oQoOKJxzVD2+IVJYY6EnOdONqEH5w3ppsbXd+knEJIzxtD7PAPRG4Q4veCMp3
cKd9Tk8nJb3u48iOxMORk/75W1Ep7QuZ94i64p/tv56hDKRiJl4Iex9Zq8LZqKtnqbrde9YDf1Uk
CJ8ujhG80fZPzKIATRQTMcG/yzfe5rVOCOQIaXI5s3lQEOkpCk2F38NziFUI93cqy8vP7qTSEMfi
szQaXsPhOC7JfYGx+un6wtRvcZco0obew9zmw6PH322Wpc+rcSBk8Ts0OiT1wDtVo7iiLCKwbRgL
ZfaMQgi6LlwNi2vy42bWegRi9yflPbCvj7Mmkmj0+M06kkZi677ajpoh5GBTfYAt/vdGOhsKTVY1
E421MGfKxHKTu7G7F0enSpsTSOQqOGxeLUDV1xChzOlOktCjLQrAO004jnTLjg3WL9qNVVe303fL
Rrfro3LwG3Hf1muUIWE1jbYaaraglQOaTvJD7fuxqTDofvFVRmLBOlv3uUk4ru7Ge2q284knEBgD
gsZYLMf4WehjnFlG/uGxxSz4xtOrgYnkUXl6TOA7Swue/U5PVZE7w6RGvjpcpHsfhsQJ9GuEb9MT
3ymXz1Zay2Ov4XIyO5vkOLKoJpdraK5fMvtF7d394vDiGJzD26vKYDNcuX8bFY21tzudmKvR6JD+
1FLflRytNnWdBe0u5fBLnqARmA/kjKty7YJ+Y3MytSmz+k+xIoE8slNs/MlMfaRIB9RK+KkA8DzV
HKLUVj/p6AJuskRO5GGEtkX4WBacWZTkrACmK5UjQz4qAW/m1pYA70yznJmg5R8TESZJn+VJEK6L
RD/8nvgFv3g0WZpkhgS9HwbBhWJEE4+9VyPLoXUtXVshd6dxdHTK8FZb4ulr7TMSdTRWJIByBrxA
OLI/t/pNk8ewVnzh3IR8P1HDTNm8YYEvTOBjh2qFYI+RZDwilcWivSpqgAyULzJN28iDF9pWSAmS
0zg5tsKFMT58WdosW75dbOIsAU6yzOOudwEZqyG1ZCJxQ4zFpQM5eHF1qw1yruRFMzPgy1hDgghk
1htVQ2ofCTuQ5wqZjJyF4MsgAqxbwj9gkMmF1n0A4GhmKNVEVck43UtNpteTETfTdcrlalYTGfsc
Jc5BqkHXN27IdwPTEmeQmoeNrwNQz71zJ4mLxi2lLylcRJYa6KSC2YA7gveVoVnT4RUI4HPyQPMa
GPOeWmS1eE9X+hDzxRI8pu5oCaMk9gCUkxSBDP6AvstJ/ZIFyGACeG4DdT1dYWyo2FuSoigCi++9
bk9s20275wse00KG+s+Fe7Tq4lbQ4XCjiPCzt5h2PSvhjjdq8FfzSU35/y8mzsgwtwntD2RD2E3+
TwaUKkUhBt1BjLFmFdkncuSvPAdtWxLD+FpYqLcLmPhzjqqVwyfNRzqdefFhO4L0mx7RA75QvxMS
WvLz6RpUBMi6mcG3TBr7LAmDHXsAzoQq+qxZ9Qu3ojufJ1zciMg6EQa4l7MjTSZw08JCDnqg0mQJ
qbQXfuWwcM/7QoR14hD4YpnM8GFZ3hhjQA4dedZPhRqMkQCwnLc8qI6C/u8o8L6FqrRTLNdHeplP
XWOuIWR+QbmXAiZl/Rog0G2Yapx93C47cYb0UNNnM54Ng1RMTwIm6msibUPsf1ySFxs4BqnrVYLs
o37TSUrhLKhB43y9yqA7TbJqB1+lJczCp73JDkPLWSDhvKsxJ5WGmEQBPc/zJlAx0laKrNC6oc0N
EEUnnv/shUAzraAjfcNc/ipbn2nVs7wBTeOWIcBOrg+hHx3HVcdZ2Y+joFoa1fuOOVww4JZtxcqC
YuyAsSQhUO9W7CWzP5RM27QXsuMy/PAfo6WZKXkrxPHpromdf+343BgD4h3Ci7KvM7E8wEigK8Zl
QE6BgNebLDKgXH5bY61ce5IC62NP69nR7IJTw16TTQGT/PJvhV2ML2ucyzKdMQE/mDIl7viNVqOF
l5i1XCaM1+Smt2EkdqIzNDm9LvzHuCrQ8QRmurlva6wS2sB5UIHCuiYcrfI6tflZOI/M4XadUZJM
iB4NEj2pCusdkK1S4+5I0oFqMgELJhkBbY/alh+nBVnrr7oAiD2KqPximXoXy42i1CgSqWAoy2Fa
3vNGan5t8IxFma2bjcjL+w8ZfLDTQ5Dolw6SxXPoyLvuM+Fknbodtlz/D46Asa5Uj7xpXX/OhvlA
DuayOgTnGkt0I4heDKfJPmec46eO3WHW9F4R7DV90pJyUhlCzjRlHTsU2eqdEK7BoHrL1uJblwra
567jqeJWAaJffUtbZ1N9OIuXuuRbPueIP3J+YYmyPWgrIZtIhB1c2wy0M0GpTGyjp8H5wZf1TSRL
X2cTiyCj+Rh0rkCiTF6dv01VKpFUlZ7PVGYSjxWibqrwbpmIBkE3RIIf3rd9FIzhKShXZYWFBwM9
Ptbl3gCzjmgKHc9pjczd4/rpyo/tbqG+62+0176QyQ8NLBdzCZ6Ueqv0tiJd37PrxkRE+gjcCMmf
ejQfrHvggcjA5kj5DaPw/jeXNgUz/ypMMharvXPExRp9ypWuODrAyayjcbedQA9Rqgg8pbvTdSNk
k0kD0tG0XBn7az8GzZwY7uSkkI4e9mJDcWi3OkLPlXzc6ngx7rXPA3OegS/54WjxMDczDlJa4Beb
JdZshYXNmL8y3AByRz3VIWEAnodb9yI3xBwDc+DArJsp8ZxQS7G/Ux/2npr+zNnCZMYw5KC2KLeZ
uZsLTcTzGUlYZLspGyROgwaGlkshieiv9bVV1BgGMueh8cNcctTQt0XeIpKV7q4wcCDnmszJSGyV
2tWFWXn2ttoGXT5bm3p7Whq0zy6aJWEA+y5TiYCQZSW3OtI87hLbs9E6nPl43TXTfpMs7IubN5PA
1Q6O5gj8tp4ns7y00pCtA5aEQ780F4+7pqbI7vgYDiu7QAjJz/HkC84QHkr+s5QloRDPBw1SR77E
0z8aH9/NkXHbcYGR0z7yGPhLlI7+nApsJgHYuga3apJomJ42NYrmt4yZl/Yt/467CSby/XamSqLn
/iIM5bDTAunk4G1SD3ggCJP2nOALmQn/Aaml5yLv+A+6TSw6v6IDkThpXuL5Sx2rSiMGOCgTvPyn
IVMj6Ujk2HW968QpDqFZicTNrrCU/D23zN3pDbMYmNciL3wWaqcsXk2kFdf84SZlA7xOoIVDqORz
8e7yEbBfOBWxGOoRt+rj7Rzg4Q5LfyliMt5GsYlJ0NVuXAs+AQlSYo6ttpKtrB4HQZD/h25JOnlu
so+Je8vIH9RK00P9m+ye2LwUwXAHehLIb0xKdN0a6a+QZaRpBb1ngcYUZyUfcHJfUNKx4P0uaR3f
ZpeFZEsSAZPE+ZFwNqveKieVTIbc5b7XS96iIKS8/bhtuZeM5aBc/6eR1ZSeHnxSg9QtKwvYhck8
DXXgQAgsRi0ouqO5tt0sH6lgfMG1lX3KSb3WdaXK0imghUrbfc5lsUmP2xXN6sKd5tieZTL905D0
DU8mJPYocozX5mf/a9jpBlGZyzfByZa+AJN7YfUkQsePSGs5dQkEaVWtMe+YvZXuQrNo0Um8YfKr
DaLcykOq03BuvSozZDYESE27xoXYBschkToFzsSHhf6bdlen8IjQKeUV8s9WQEp4m4VCWpmMHhmY
X1VE73/UW3kf+9deKKXlrBVXXZITY0hrZ3uIIKBpUMlfX1osYOdh4kL34JTQ092x1CioyFQgRGfa
X52KxEHkOQULceqi1bBpHI1O5BmjjWhRzvca1NPz3E5L+qheGjcocn8CMI9afOnZl6yX/wZcGQEy
dGnZSpPUc7mCRQyPw6mhZbdd3bZeaGEEJxHWV9nHnxm8KngC8ivIyEXhjFW9B/sVlIOcv4bKMzdB
dd0oAW8c9iduHefitw0ijJK5LNVuacOLhPkCe8w0z0MccOsXzf9dVnBvSaniJdI3j9n/tO+O9Mdu
NXvX16jDkRYGCAvP+LkGkti5up7nHaxDjqIzqr225t68N6R5W83oIdikIz5anVvNklUqT94J7eAa
jL/1Sq/hLv00/RnDdPGSk4vq+/LbJJCw71ezpwX7LZ6SVT4CakTRyvZTdfXBz5uQX3w7uI6Q2xo6
9nZDUquqjWZrmyP5pw22oOL9knndmIKY8QDRljERrajPGjmAe6kRHmJlrdvYH6MYjmtfY4Y6IjDI
1zY00xwLwuuHqWRCw94ko7JhaTVmb+hBwIcjJI/3ADLqMGS/SUlk+QFbEIkMSKersLzvEJLgEI7J
IwpE8XCitPwvwSzD0XUE5KlOvoy0BtObx0bJ6BYkUHUETmgfp6Ha99pKxjMuhw1ZSa2+bQ7Fgdaj
GVk6suD8dKbhslRzj8LD3CjW4+ljSodkr4/Ldnr1yPo2VFXprPhGGRytXORz5sWgmxO3j12Hyl6a
YXkTYLRlTxDn/yehW4PrbXFrq6IEWO/Q3S5SQzK8QJIT9513a2EHYgQ6ZqLUDMReFfxzOuTQg2v2
cbDQU86j5ME8XgjC4BxS854CnEfJZmDlP4f/2YEc4Nk7Op77XRnpESZNV7X7RYdNMwMhNgT+KeDD
nhDiXaqcKVFK1JegDLxenGH4kb8KIexrsVwX8p1zS3/2V1BkvhP1mhHdZBt3fQPa0daA4ovT9Kqw
GcnUS6qHTsw6s99EB+cxlT73RsiSEnZW3PrHAp9hAs3HG0KNB+DGrMt5Sh2EorRMLfG39xoAX+N0
VPn/dgXuGZCwtMIFYXLOqXYuSTAFEDJgVwfDdn1ze2gNp76gkkBVRmxjeykLA0aRQOyuleg1FrJE
6rSbDkldi79SGl+db1AYI0L4HsSy5wELYkwLsQA4V9D88XYl61OU8N2gzAHPZQ+waU8nXcRIpazw
tSfH/zg3hJUMXm1bDFjYkQbTtBOWd5X3RW2yl7PjOFWTO31Hg0fzu43KeYZx7PaGevjpvtEXeIV/
KYvix4mcZHnuJwjtyyYvcSH3JFvEWKB0JZ0aFNnSuJJhg+EycmZzE7r5rZzU+AcQpiF0gMHEZgab
pTMQ9wqv9rfQg4UDeN19L/9CZviOcsLixwF6TOxwkOrUWZeNzxqKUlWspb8HW6pNJ4Wdx+oekFVB
hBZyFZd2nVdci7RFiuCOz+H/OrBp1QxkQjjUng9fT5SL/x/td7fydp+RP9Q4bnAYKr6jO0QSD2MY
XGHsVtAeZ86AZZILEKk5kbN/mpSNVlISqZs3GyeUB8yQ0EgCoKxI1NF3wiZOOBnpPM8HcmI/MQnt
+tz4iOqjdL5H6knTh7YgZuqDsZQ+mFbGqtLBGxsAbbK7KCcPJvyT5SBDDUhlc00LqQl6y3f+fkPK
R3mAyJtmuA6Zl7B+aU/m/Bz1kpUeYFbXPIr9tY0b5Bt0DdH61n3FuHvOx0rbdXkHtor9ZolhGGZ9
36ZFLTjnEy0//pNF5YbVROqrxYCFiJjk9VDEnNh7Bu9AaHDcCpHUtxoX2DMWU4yjJXau4PVf5u7x
U2fH3gMABxyVBorhTlbj/wmpqeA/lW7LjObU8/sJXSNzRCaR3KGNv5w6A+fYkRhucz4weJAAGtOG
+4Yvi0Yw22rhR91H9jsYFMX+na7czsisWjmP7LgPblVq8Ym5oOZHAW1Ace5+u3e1n22tckJo7zs6
hdl8E8a1TGio3oWRQoDCZtS/r83DcrIq7l+naAG9VeeMYmt7nSWQKj+Oqpaik57PlNSvYkgT6SBc
sinTckNdlMnfMXr24rbKPvssxuxHVVwiY7eVv9F6DMqV3ELluUqpZPVlDNb0hijoMn5rtVOvkdoG
v+HZH1oA2rwkz6RO1AZLQgl/sQmdwrGIfQqXPm7TbYDGeVCV8uNSeZUoc7PNjfdi/tKdwPkfnCHU
rBaYtLiqEjy/Gpzag7iavFQqa2wA6xnKRRb75QCB2Ev1R44nFTRhgQhLbu7TebPTRBI28O4yjML/
mxylewFqrFGwWn/9rG1OHw+l2fTaw8TVmG4u9XrMdf8yu+C4NkIyt8reCuf/Uxo3CQoxewwa4CDw
Ynw0kjZFCbvfAvrokJgKomfjpKee/h5WYT2QNT7v8yjfSdJEYkj4+GmC0o/FOpWC3grxuN8KPK/m
7A554HHUXUmZPm/TQKvhiOI56oDQ3E5pYAOqdvSoJEzyjMEzqd+ZMRDKFMOkKfsOvggoK8VB+DTV
IB6VdvScOe8j+cWCRPNi5e/uO6ZnXJY21fS7p54OUYkG2s9XiKFdRxLOgd+c0qmzKJB+Eaid/Eer
IK+XqUuk6jUFzKEilw1Jr2MxoCGGR9LxV3DHX48ravlTGfRNA5Q81895NzonEk36X1vjHJ9eL9IJ
ECcgovwttfpDsYkzMjuzDmPcJlMw6+PEOS0iUAJ2Fzkcc3EXHzuyfovvc1YasL8+x+vc672S0MpN
6BtGush2rPeAd6o0KkfAoslsmACYWaIyZGm5MC7iZ++PZusxPFu3r6SKwewBEiH10mtaX4G7eMZE
oDsYtkIb+vQitSsOdeLNELBb2QeP/dApKsOhSonbNFHLVX5NlpK8J7Aq2wklKWriJaHPW5PGrh91
hRAJ32iI2shRfVpDDbZM8Xyt3W9MzHwu0FLCTnwGe37Bcrz5mSO9aaq5+l2hQ1JxxYptwcgZhL8j
ghRETkNgEbbivXE67O7eIeRUr1rWj3fiQh3r8Kn8pWiDuDTPaYvgSvrVTVtoQLS7qYF5VsntR6pu
Nj4+YV4wjXAWqThAyI8qFl7zT1bu74GACMCd8iPmz/YM1EcJLpAr/qd+WRJ85HaOk6ZIfEgGvYMl
gLKNpKZrk/2SX3EvBlfmHOBV+xwnnFsaEaG1c0Er8OOczM0QYuJgLvPojdZc2y7MUSmaCM9HVZv/
eA/hmSHUP2wTZEeOFHYLUJN6d+t/B+Lu6YzjGHrJO3jyDGvqXCvI4ENYhn0EjevgmaRI1KOayIDr
rrXPGvSMATtR8lt6a+EBxDwwFMwiA3JIURN3lFuELZSh//BdCA/G26FNZHOaWyIPSOkbDzEQKOCY
pgyglwYFE7DbZrkdEvMmhU9Io566WwqITmxmBpx6tg1t8QlScayNOmvf3SyigP3MhuBcrv7+heU5
DnnSj/Vl7rcqkoJ6phc4PjKxqwc71AuA7cLOl+hIDPOIEuXyOZ94mDyTgL0HcQGLUr8tI1uo4l9d
6o4LPd7xJcSFYl8/ayxVjwnX8C0O+wEwd09vm857m5ANpUGV8w9nPMgyhiTijQ44BUYXj7tsHsFG
Nu+JW8yfzS4PTNrV8Km9T613j6skRlhTGJuFKGBg3jUkcKZgQ9MO8yhRbBfd7iDmvIHNxgxNteN3
Mm2g0tTS01IKyq7ioxZCsg7Jsqe45OnKMcNuhB2D7PLayRGlCB+2hqv7ZWEGLM3vxAg+d9IhxImN
l4hmr93f5IIkAociCAHX3nNnJhxMqsfZ3zcppTUpxusTdlue7Q+K7TnQtAf8h05HD76as4lJeGZG
y4sJ7ljBQBq6VA1pQKXNzcxNWiDvIleZ8iEBB0v8s/CKIdR3rjoo+SVszA0Bg7jxtpWMd5zPTjCo
PL302S4tA/Vi+JYR9a52oen4EdPJzd/et6JrTEwj60ENmvlYap2KtWmcoQWC5hwaert5EJywCu8F
lpqpeKVCwtGEnR5euhN4tMBedSXwc0HNq8TWNvTkrDJ7ok37psiArI9vEWS6dm+th+YYc7NPHP9X
lkFLrrZ4FwjFBy414O7W/qREmX8l5YjdPaWyi6Mdfp+3zI/N5NYHsIspnUmFDOJtbSAA+mHmCwxr
db9f/2qMMvaURIDaTzbBdzZc94yu45ql6qtxhaBkrhYXdebgtlrrtLo+dXeTykoNRphudcPSFAWl
jdRugRXstJN1RMd/bsALjkTIBr1hea7XfPT2W1R5OyF8AhFBKKkODLensxaONlbo58mwFCO2RZ0z
hpfa0qeltYjCRD1DFLzMBKC/OYlE7GF7Kp2brsF16MeUK+LZZFGt036m/il6A0WNEG9BvFSx6aNE
dq7Je4HuxgaNVD6gGHf6DLqrQ1W4MHg2Y/1ojwzA4c5xXI9j8K2KtGTwgzpiFZMd8c2EtRHpO3M+
vGy8XY2Xi6QtZVXFbgajdFRaX5lpltbqrM0cmc9li7wdQZkDvrDJJL8ttKBPGgDJto/+ouo49g89
3U1NTtHr0STQV+X9r46E6ythm3yNNRlE6adgYOO1A0Tg8jC6p/M1bLlo4Msj0cDGCuvNpneo5KLI
8Oj/rBKsKgSYigOGjmllTmz1kq3BPJhySgd1yZ4NjmUIutoHlh4FLmp0tAHEEAy77LV1XKCJ5GZI
Sxbav3ZDm1PYPbsPp9oI6PVAVCaOlygKm8kGnMIh79k2Vyby966h3tsZq5pjIXJkZWqn9JRkmBFS
kwOYDcoJ3DgKZrwDJwaI2zqX7fDVE2YZc8qqf5NPfTwJlJb/H00X3739KcaA4+2YV7R4yjRVWFdX
N4pA2SAMrtrPJsSiRN0gyoTHLUpA+KoxBcJuvyaMEi5BVoWwk99/GluLOpilurZ5SbjOsVoPvjz6
pd7h004MYmeX9390FkjaEc5a19aCPsEPKBF56YIH8AssAV2txZ4jhEkB57t6mJaBlEo9FAX2rTYU
e3pORHjvu1WzhnPkS8IHjpOR2zoq3JUeoVapV7NeW4tcTJaP8d1uPmtfjQesvrya5rBy2tfRrAjs
NfmbGNSdT5wYqAAEaaV945yrR9cvMxcyDD2D7/DSxA5BCjkfyHcRKpNjUfizspRE5quaDVDKsive
/cKZi2vkL8pkJH7ktplgf71FEZSch2LgrkHIimwQI8pVwSOwdCyKURWtC857WexM+o0aYj1fJ+9Z
2rJZQzN4oFkzdLz8On9Wt5v+dEln4uuOnsz66YZvNTgSfD8SEqRj8c6PmS5j1Epj+Y/nbMTrIUyU
yD22CLs+LlOUDF6Qu8Gewig/T2Nl7BzPqWioeDgzTFw+fscshbtKZNJBPQaCq/rlJKEKiNkiRV00
4HOhoIk5Bk0tyjG3AwqSvOjqVxknkwfvGYER4tBHDhHNPbcTqX9IzUTjDnwHt7XRZUh7y8O6ewoL
ULSyQusKIqsBhPmr8bZVxPh6HQJclOiYeRyWYD0uyGBiQ1vWMVIvAhX93xZH/07+XrqsB7YHn7MU
eTSa/LYTbQpyfBc3uI9NaXR3AycBVDEhM7hWOaD4QpoPHOuoKLS6JK2RF6bwhN8OV6SJhOcnWNzz
asumFTP6oRDZg7V1CuWiFBP5HU1/xtgVKcPQyN5gKDn02nOOKfelAOTUKbzs13EX8X3FcXCZH3LR
rzgbMlQLyG2cjD8Dtq5BUu/9YhTJRDp7QIuTbx0tl/9ga5oAWWEorPjfPAuArx3PDbxGSOs+2UE6
owgt3L2ehoFkok4Szewnt5TtE75epAtsShRjHTTly3ik9kDHCc7QWh0J6VrF8sUFLlf3C8HElJH0
BFRzvvaIogA8SzbWsICVOYl7rcz4hhXTmpx3URJw0E1Du7OQL/o/POVqhNzlwfWFjyBeMDnd3HfL
3qdYIad8VxZ1GnPHho/9O9wFX4g8hp5WdJcZh/dfATOMEGB/22GZnQm7U6b5WGpaGcrdUEcwIRTs
Icd6hRQISWMGGQsJ3YSRJxNfPtukBYfTOcYWbJenDpIT3aG2pvgyspyX+fY+cYrzR8L1M0vBzfgF
xEh9C+upTtsWx9hdV5jgZcuwDDUZlCT5wg46C5NDHBlRo4JPlhYPXKgEdMvIf07V0DKormiKuMkv
/P0+r2T9IOJ46xLP2fBxATJHxYQ0H4fAfFJWFx7gCJ1z+sLlS/vxPPnXW3nX1YRCkZGKdQ8soh3y
ICghxzs3ZKHlAuWrYRvfZoRVaBWpRDhXDyM/xSpMpVP+vtDYPAMfSKvrhZ6k+7+O5SnAA7lg8G8Z
mLoyQuPC94rGtEC1DaOAEgRRJoN5Vu84VNJ8C9BzN9KeE3uAzdFnJMl5sdwThTohtk5UX1rlMZad
8sgvRe63K00Idqbx09S5rPA7C6yjSliOD8LKokcpPy5ip454uNbMl01LuaRlNXM3HOgjCm+8egtv
OBbTUBYlOEq4L7ea4VjZu+rqKSQ7mCHhD9Hbd3Zhb5Hmg/+MIQ+7GaxQsn9sUTo9U9qsn5TMVlxw
Er5OyrstiBKxg8oEbJFi8MeCCzAW11kKUOrgicEi2tkj/T5A04cQlIdlq9gRyQKs/PCD87yQH1Z7
6QideE5NzE0I6jZe6F05m8h4w7uEc8BVQUm4N4reYTGdbKKt5ZruyJqygSXn/Zb5Rliu9Ht0Qt2Y
UxbiriiTyuRBoJw5pa8HzwMpYOPciWo4eUWDL9MSGARLdjo/WVE2bjXr2WmYC2xoQtp1HOndj0g0
dTbHJef5GEHF6eVndKw6H/nxp1Duv2UzJ2Ysvb14ue+I/B4XlIHBfHIS72FuHRBi3GSbLomT6Xa0
r5Bv3vs2aALS67uV0lWCbXX9vuhUyXnqweXK/GiwRpuhD77CGQ5i6oAtkUQG5vUZ1kHBeLhHu+K6
sHabnEJIbVtmi4L3n08UI2gM1XUoyBaZpA7nBCNXtZ5d2JPBS2fcUalL0J5vBjBvFloaCxXDvG3I
F8Bb+PrKu8iy9KAigy6GNd5txLLKl6MeySWH4Dp/cB8qm3cobXC+UXJres/w0SHHo+ER74Dbo/WS
2PzL0eJfYG1RnHUBmsNG0gkD4EVrzgQHDkF3HX3EXPy27JOggcS9LK2Y9jtzgMpwd4kvjLGpnjVT
rhniQsN8bVLUM0LKrKzoFrOxGg3JI1zVGEiSQR7h4zSrb7sHzUXKJfr7knIa6eJnEwFzie/VRu/E
VhuGMsduhw1jobl3H261UBMoGovzYBAzaBd4w+iqRxFRp1pijnefOFt1pErOvUWYbMCkUJAU/ZEv
9bmtx7bdLPq9T2J/UF/hxriQI8UX8t9UyjbnBfle6/qw3usLvkrUkpXTDJWk3s8ToPhijV/cjQio
iJ55/TBVJ7a8lKBUsbpnN2zrqnryqii17dC+C+vnk77jchEkW/9JfDVlAVM8kWx1LqaJCRWQFAss
XOu/vC4PyjCY+2IgulaPRr9BxWElpDu8aPxlvzaL3IRThi2BK7qAiGFDOh1jDyrsr6N7G3TXZIIl
aT3v+h/fMNKGzZMT0dYWTwBGfZ92GH2Ogjfg5jDwtUYQTNxW3feeL4MLpeiq6RSUf0X5epY4PGzy
Oeyslyz6LjEr0zQkr2ppaJDRsSzmsvoYnQhQdW2NQuft/CTlxh0QCEi//J69NF5Z9I5c3RkmRoNT
oXp2BBQLv0qhA6S7LmTjSWDLX99z6TQd2FxDYDAmIt30N2sNho5xiRnWvrXazQmf5jWAwTiPgXSE
F/BaGdON0vmSyoc0UegxNg8XcpcR7hG4irXG+yuKvhM1kVpeSa/4L9YcGtcU6oa9qTXYgYRdY1Lh
v7VIjur0P775Nx2gZ4Y1gg4DE4woSOrqLNZ1PCSh8aRdZKVzgfbjcEEMDp40pEvU4cjQVcpbPIpm
/hmD8b5V/gZvj8eDg+Zsf+oqvpWiGDxV2MjNw57InLGFyTDl+FKzCb5lAEFAmEwqWG3iH1lCimYE
+zeSU2k5L5idlx0idDdu4IYFBaoLZjtvAxTbL7N+g81DmX1mxKSNE28hUYCXEq/ZOGZmkLLJ0daw
lMGQ0pUPJTsQOzBVMsEXTbduqGRbNi2bsVr+8Jwri65ebrDyZvNRTfrSIQLHHgjD/gxpYA9ZW7J6
ffjQ7meyWZQEue8NKFwJlhadSOzONbGOhG1pYAj+pL0rdqivPkxAC8TEoCyxTUtINB5RO+2cf1cc
A1SqxKtc5Hlw0X5MM/SmP4DB86ydl+gnd+2gdh6lIoPIgh0zNlcf9M4CApALP8W7OTyyLZDdn0J7
5plBqYHVg9x/vT/nctYPnSi6En+PBQYmUlSdQboVQtLyJnBv3/98BJ22iFc4n4I5A352XuxuQ8Ou
hmP/yaxyYXqtFDRwBOuWofsn4uY7DIBjcAYZc8kOYS2Awu0RUOaQlUmRWPlHkhiXh2ky12wmifBC
cnKzB3V0c3SGrw5qNPclTkYko+ZG7RIeok+FIsVMQT0kqNQZis68ImuNQFVmGxWLszudaZ2RkRYr
eU1gZwKO3sxHUV1e7NdkrRi8p+gqJYrVqYuf0kh0b5DppgPeTahHbEM3VBsKprYsHXcWt+PkXcSL
wGVNhRPGGXEZV/9wiCu2Bd5hndDbiInbf5OgooGzMOdAMO1wLwZVORdDu9Xb2DYLkbVu5ssQE6ic
OClT6cUVNZ14gZDuRBYO2BUmWwD8UiIWRTITuznF7JGuwC9RIZWirlTt5+pZxO1STh24/6mAC/WB
WqxOssxFPfxDaqGptUv8xMFostFOxwy1CYamvxrBFIkE17ah8IK+dOQ+ZA9hyNbr5neY8B7lZizu
b4wKxrJdDSi16K1OE1MRekdvqU2X6E1EzVcGR9LntguNCk06I2NiZ/pXl+ZWdz2ArfIeFemH4K7M
mjWyFWFQh0Y9ZadCZM3aJ+aVtFA6fD8J9ahVyLaSCiss/wj+DBF7riAVurCEp65q1SKbMLh7EYx/
Nv4Jo9YhBviDViVDVktx7vngA275mXSJMBw7ssxVp5MIhIVgNmBu1JjdVvg1ntkznYbvbyJUOXJ5
km04m2pBCouAV99+ILDfc1pT4TwYgqBp1uafnPNpU8H+Avwloq3lOd+u7Oke0OCsZ3wwuAtVLNNw
snFOwVPXN3fVeXyPpfmFBzKPn1iTjuAfxcj3SOtk9MGKhEM4xxxiTBMZXMSHlktfKjVSCaQS/cck
6EtlvGrqo2yQ5eIaqWtiR71i7csR1TWJ3Y50qP0PgYbMCoQSIzhbch7Q4+xrKNZqdnkC2UgfiTjr
/cpFqpWJK48uMG8T2NMGQMJGzsQr7nGCdRG0ncY+bsntNM1KEFgCG/2kIHNCqTvFMrQYQMhztaFR
XDT4pqiZN8JrnBN5tYOFBfVUpu/w2aOYF1Ewr1prd07bCwYMbc4WXlyGf2C5+doOpRkYCaAXuKih
MVGzo9SW3peOav32j4VyZbqkqiRwk6LGNMKV1vM9mMUSYfrElWpTbN6sbnVUp41gtMDkd0+UgcmT
CiMcyCBeB2OYMTZDozVidMHYhGUUA4ubAB0w9s5tbOjaNbEFjlPICAGEeZUPtV8E+zx14Ijs9Sh5
sjHpjgkqxCMkgb8g2xRzRE+J0zaDJbDuwaJ5/sdla9onOiQaUg2dlOSi35JwhHnSysTMtODwkNu/
SD2vj9qE5x0BZmC4GZ7uysjNS1OM3E1jvqIHJ1OoYQoTK2USbxRnE0vJTX2dH4FbHe7ofhRj2+pw
92MNKo1CPnjQwq5f6BeBM7nPxdggF31q9576ij3/UVnn385+xNl6a/4aisGBDWfkhtYXY4mj6jov
Q9d+P0J0AqRlpYlyAgLwB8G8AKCe5eRhPRiWg/xoDaY0X2cOaxAiGQ0ddA/ORM3g0U/S4t0mvM6J
LespzU2wlHWzLb8ZZ36rDxAYqV8L4NVveF61XtZGd7m/mTMvpTxq/F0PJlOA+ITpQ085H2Ugveqs
XmZghdzk4ZzaDUncBcqAeQPXN5IRC5VOjYbgZrdSK4CM/S9TqSb+iFQDM/Vcl1OEGcKbGTzjySEy
oLvNBcHlGGBbE0T9NiWG9w+sw6HS8y4XNYpDI/FqAB1CwIlF8bhwD3Y9itM6wse1P8BeYpF4mN1c
TgnMaxIk37Evxz58aj62H1jTfpCyK5OUyHJpE/VEfXxsn2KRXNkV8+pwdZksykARTeuItPWOXMxf
pXoJeTOkfdkRZ9NrnFsUFVmBZ3b1SkM16CwgRisxuXCT3QZsneDlohXEKCndJodOboJJWLCXvWQx
aPTicD2mCO7zLZp0VZQAgVKu3Rkn5GoOQX6ZGNqs7mVkoLndvWChOnG49xiS6I4tKXMnDrppQP9/
XOJz9vwU3k9S8rRs3jE2L9FVYuoMCvYvjoyuVEN3hEd9WmG3yRC6zO9I1Afg7H3eNjM4hrmSGhVS
o0/iNSJr0lPU6vV0LNRmPQrrvt7ntQDJRtX/F3Vy1oroOflz27nMnIBoV3QgB8LuCYF2smZzKfIe
BCJ9ryrWI5r498WCN/IvD5PM9W9szkBsP1cNQIWUnrUNjc/dV9JB+RUGBdeXBjAmkeiH2TPx3Hn0
SPFAphwJYJwssopTIeR2ptTVWAOizFFhv4UJnIsLdPEnHrA7HW6ixu62GfYxThT4ka23ARO1ZebN
08tz8VRDIEbvD9VzhYG1MvDSbEp/yJ3s+hFP3uXBMmqgGONKw3c6yAB3WjxN4+AsH5x7J4Wb9zr+
WjQpoZYKFx/70vj3JHOgnOP3t3G+Qia8+J/KcfDQFpDSuFsEufbhwk+m4j6Tb80RtHP6fFHfZB9R
kFsFFXQrcBYG3j1P2iXTOiv/hVkoxWmZYiYRgH563JCEyDicN7+1u2WZ0xgjZbKW+5dAeZjZpj/y
AwH3iYw1OsUSFpHDgZ/IguB9bR8m+vrZ6dUisRIwXL5/Fj+it56Ccw4tYmgXmEzCKBoL/KwVXSkM
zNZNAV39w26LVSAcTZwImkrYTNwntE/IOVI5O+TAtk8TTEmc/bb+RephEIFuI5/FD/xH3DQTRVia
S1ucDQ/9h43dZU5DyvKIWXldbjL930FGf4HPejP1nOZos/RZRK8pw0x2ZtOxZyCCncx/J9zB2aWR
M0QShybH/CTT2Eoxmgqh/LRCDzEu39ajgviYvS1N1pOCTZCtzd5V7C9aLly/5t6ggc1fCItSd60G
rQ7qgXOpkUNYpUDwT/n0pjHXist4hafz8pZaDHAk/4mGpm4ZnxEEX9CtWlreUibSqhNHyfJeTyHm
8I2IVAp4UQSlDj+3uOKg4KWRLcmEob1ahwAGZQARrXIJH+LTwoRqjbFk3zPl98cRwvqMi+Yysc61
1HFeL/vFpdWnfk9FDyaSXmds6UlP4BHWTZmYG2JNU6c6532ga3ssh862gxVECc4Mp9IUeX1tLz1r
Y/ycXoWzDtMXrJN0OzptgMYw4hizC/hGKw9+UwwBOznnUaiVPY423iBTcWw6sKOTXvM6mkm0boI1
D1W5kHQzurNlVyuSgRU0pLp3xtQnoR1yCT3Is8RRJvege52n1ytb4e7aO2W8ZmOokiPqZm7tkwGf
E2lcSJ5quYQXELQKJ9VwedJt5IcZt4D5wtJ6GXR+LVDH9UgjceHR1FZdHFO48S3a7gsjTfQj3Pbf
D6PVyCWU2kr5ETu9vM4MpSBfOVRu8+kXXwvFYbPY8XcuwPhS7v6L98T61wo5KRsPNsoIX9QkkSmQ
YS3UBbI3UxeZXPNBf3T1gUowJlJuEpPilZM/UQ2eVm6qOcEzGRQzZz7iXAOIe4i+SqwK3hJ6ZH+5
qBzOCAuJVqeJiiXgR01AFduEEm7NwGbHyKWicuqmMiQZGSwvkfy+WY1rKar6pJ3tIVCiQCfSyVXB
fx0bv5s3dCCVKWU81udQKuPaNG22SESxN4n8LlGlwgpk02QeXP9G2Tl0bx0IS69CUXukSQZziril
1SUnvX4vNkWkqb5Nx+QOxro30x24ZZbisqma8i8Le4bWBL/uZhFcw47QkrxmHAC2TZzudZNzC172
szYX/p2FtDKcHe+M5QuRUXaXcNaf3Jmy+ZwWzzDMw9ivIut5fBl5WkdhpeHaF4QbGbCdMCRgAp0W
orvd3/yxkEh541kPkDRHk56SGIWcapZSlarBgU9rCGIyxtPJQbDBwkeT55POF2Ycm6gwrTwxk/dd
9aMgzJVrRYzLqImMXKvFBVo1OGVZEEaoET7AeXiLXsc8eqZhbUduQt9juBlda82wxtbHL5zL1JZJ
Ug5VrUHwrVHmEVoRSFUHkSXC7y2xqsgK+M0J/cayXX71TTcv83iQt8kWSHMr4DNvQ3OUQGPbc+ja
WVg8R3qLJ2Ivy+2fNcyJ6OL5s+v/ojwwiY3SVmzM5TQ1N2JBbEzVS3PtGTk/g5ZWNWL6RQJ755MW
jhlcen4xdLvacQ+wWudYTyKPiga+toMR9czlhCL1W9TtBeCTfezSwU2g5A7fu3stqHZO9iOhbnxw
d5c4ho0rlGgdlp/peZeL0igsUCZA8LRRqJ+Xxfmrmwl3lFEU++no9ozyc414J8SK/OGNKxkCyIfh
PfI6dD5tQ1q8+sQdoYEDKQZbbfNvKBpfIm4K9MVCIqUIYgJki/NGd7LSIcqQBKYMVmXTGLTd+ZWC
k8ulwNeU+aemTGql1PJtswhb+PTrSqKn6/phq3586mXlz20pcMp19O5wr0+J7FTlHM3Zdj8AwWv5
OOU6w+MTGhFY5Ix6mzv9laK5bI4OoaBTMS2t/b5PGSQLrZ9PYLUkCdG1wUSbb4KZWC8Z3JcEyrBc
Qbw92IaEROfx6R0CBHf5ags+neEtRsejqh9TwWI1HsmUKfl01jAFn3H/okSmMchJuNNqH9uLnWih
BvrShVu50NrCUt/rnvX0wawRoHApB+fJI6Zpc4ICUsK9PLr83802C6g+93qLw3tATFABARR4Z+a0
j/LDnsNS5WbRyK0YVDR0AiUPjc0ydHPDVHOBiNx73VvxUXpQDs1AZENe2AgRrGUnJzEyELsklWuo
E+9fBwucd2rNb+tPAkfX45KaCEIwn+k09w20qpinXrXjogXqFQhSr3sRo5q5uzWf+fNChfAjICK6
CqI7hJLbuwTxlLj9a6kjxRP7nzY4anT/8G1qlIQDnPPAAaXRGojlt2GXWoM2DHyWz2U3W8Oa4DlO
Ky2Q6gSdwecu32VrYxPRasbkSCOI0U1KQyJvscKVyhVwjDx5XFKWn0iYF+VqbGUKL4wA9DbOqvrT
tnH4HD7w7Q4HiJUnMlF0LkmbHlGfWxi+4S2vq6/GmdUklxNDw5qymk4EZQ4RvCkLTSPAIXSVSG1b
4SC3N/AdEUUfXl4NQe1D4K+Z9vHzWKhd7towDIyfNYTV0Rw8SUBkKv6mxZ6YScAKSZ41AcdtqRjh
RhM/IAVQLYtq6GMEEb/jFZW14x51eY70Q2gxshocokL35aqV7Ot64i/HE/WLwL9QdHy9mNhWIHdD
SfLxjRr23C+ZL58OBZQFWBqHZKKCZyByw7aEUKqvQl718nj3U3LSDUJgj/N4s/dUDzV/cnhGxBh7
JT0bf+nApsgsmz6RQB/cqL0xwRup5gVpydoT0faYRxlqFX4dtwGqaahDjnUNWqQpGF51ootZQ531
+XidVTq70qWYyw00fI82kSML7qYTg//a7eyHQvXdKXAyIWSzAxiyTqsATLZzsSyUwnOo0226gawz
cPNZlvaugJXp0WoMbrPoSZDkx4Kl1R+GumOoTt8fy0MLCO4zx7Y8m4YQuCfqgw1llUBUVXp4jwSb
6kJwZ5FBy8sgR65fOEGsU3mGrCb+reL7k5tJ5p3ND98VJd86pX7TLyCo/84IQCPfS8WXEFbTjh7T
Wi775o85Fwo/6A0yRKxk7GGTY76Lt7/TiWN0H3IDVx5mtzD6HirTFXYr4S4n74jSc69AIj2CKpxN
q3Uxi4qL6ZfpjPOEDzlz/tS8Uf5OBDn/QgZjpH5TZ794LIXqBm1WY62SMZ5i+AvNzq2EVIZ7YagE
Yc3qwn+SOtGJhdE9eNggqD8qydSoHB+YaMRziIE7Egi9Pjzhrs3n3Ll/gwK19kpwyda+gNIARxG8
A5gLpTQvAh3agL4rPom8Aw74QYHtIScpOjlkZjF/jaKl+Vx7ujK52zyJbg/AUR2JXG3AoRiwmo+M
igv5+U3zwMgyJXBPu8vcn1rdxWariVz1KflGTZlpW54pNIuyYhmhllUb95PLxE3d7LcXWHhCQ8G8
YAw2GHQ+VWQ0/Nsn92w3N/59TFveluWqzJo7/nknQT7UVV9uAc1DHnGW7SZ5bAFQfVwhq5JbBq53
R9LyLF6I8/IKUx9eDVy7Y9bZsuRG0f86GsuYojMwvw8T//S1fIxKifKZZU+nBENtMaYqs2Lm4+i6
X6JWBxSYwWIzfS8XfA7Ztyx96/7tbipWdxSLuFT6TdRpMvRJIQwRmmxry3zrkJxgxFXeLu+fcmjc
M/IrvbcULC/EHy7vv+gmdZQNtYwwLcrfAZAhn7i+uGWcgDtv7rI4mZwXoaK7zNkseK9O4fBMwgF3
mxby4NurOYjTzFrgI8FNUms492MdjpvSjTkHImiY+klr1rsrdC7RGnK1IJTKczfqb3hEo9j4PNdh
8Cz2KM0NZzeVdeulBk2vg5X+M8XfNB4xngViSt7pSjocjuZ5Z8W2eBEmgBYUGiKepfToTUm580Te
MeKGD6YFci0wOddsCDpxSe3gs8kXlK+40d5acwKXZSQsQ3cVYETYjI/msDnA+7PmQIAwYVdOwdgD
UQreAcUBn2g2BthpNBIyUPijKTGXybQWItQg/etSubHgKXr3yvx5ENglNxNO3WCHnhB616auoJzO
0Vi6Ri4+q3E3pOXZh2N6mYQQucnsji+1QR+GbysJ0epxmO0haWISuUJGQx7+/16x4zPBlKCFF+V7
ArD1GutX/SPlUGAsxUoppGSqbLDGMpkc+p6JqF6M+IfrBU8sMBmn++w6sTKJXhx1V4SP7cNGOrFB
A7gFudwtjcY0L/3zWE9/uqehD4hutnTCU/1r5ftyCYyk7zh06Sac2iU9WM4PnGKRoUzyYcwgR6UI
03Nbh9+m9wvyXfykLJdnCHOHXcE37ZmvHRV7Mfsp1p1ZdaJ3g2xWi47K4SZUl6POoS8SLNE6bXHa
bIGbzfSm5bRGgNesn5iR558BE+81aB16jfFrtI8YZcvV+1nt2murueSgi/m+EEtK0v26ipnkPHeG
nL+DTHXKmQpjcFCwtvNeJBEeQMqffkIJ6cGxMI4FesKfzS9nI6Ya8jymfgi54tRGtKLbWgVIcYAG
1ozxHOtOQ4olH1GZKPr6+ztVY7bAFVns8Ewki/pW6XBPFLjR+xaChkKsyZHlXel4JKwqn4xKh97/
VcBpazp4KmBJhiITkRuFti0brFOjN8RmRjHNDarhqLlZeL9d1xbtcuYokGOHaTiX/9jKuWNdYwUD
MKxTd0h/TYJyKegl21WlJorit/78XXPadkzLNs+joFTpYJMoW+yQTlUIvyPYdkNGzdSRPXo4aZ1L
58c9A/4dx5eRe1pePSb3rRqJLtlwKqLXI+KIq4rERQwy+YwRdp4oGzMSAzg5Me4d/TQVOoX6YkLj
EbP8Px9C1xadMCv5llXbwx7pGuaOBJsb8eCeXNwwcV0KEI2v3Rl444JNKs4PFKla4/MUyoU5doco
0ykVqUojNgM/ZlKtFe1PJs+tkdm1OhnnXcOriXSdjtqiK4Qftqz3UnOYE3osL3+C/WX2DHcXl0Q3
RaQC0D+b97efGMZXvRnrd6QzrLAPCkOk3WKFLD4OGAYQ8h8Q8w7r3beEWWsrhRgUCsMUBGU+byBS
AzGdxNpL1Zjl+0oiUCoHyu8hBLoglm2EDeMbvtwnRC329IKME5liOtk+MPw3+pzh/vca6zRRiOsZ
ZNdquFOQOeiEeKfRs8+ScjqWWEFxAYOAVAKOpxVbR98S9RK6ZxllZqavynKe9B8fklPT64sSNwXx
LUhxYEVeDVbvyH4sSn0ZqLd+3TXCtGivaRnDR/hUgnS3mAdkoYLFnpUXqg85Dr+3D62baclwd0jd
RvlPkbV4nkKF5CXY/bBgPErepz+/BS9Tjfi13s7YciJkqi0mNvrZu7o+j5miceJcrtGVXmtk7Gfo
7M3dJSXbbtNKN8sOd5HcON4Yn6tQ3b5zRroVEjly9438MO9iWTk1GzuQzs8MKHxJwMcUoObDq3Bm
4qXyTBtk+qtQzDVLGcBgaYZCOMpiLrQQyg1ZOiW34Dae8ztpk6GIilx8LOu/HLY41HPb8kir05w6
P7NVi6hNJt62oyLQqNtjc7764R9Q64zxbJf4EE8MsY/fymmpUCE8wVmhOLExloBp0GMfd/14ERtV
+qYuHE66EK+RLZrC4BUOxW0BTvBoelpparILzZlcXo2g0cIxBX0b2YFakBcwVHHwIIhm8iSpkrwf
dsuMrmygCNsEhToeLEaEW/smciQrEadW49SBa/EUXHugzZxRYV3ZNHxjyz4rZ8u0md90t/oW4kuA
1uyLgfNprWO53NdjGWbYE4YSfnv59M0rimoPTWo5l2TFMAOd3sTOb1pSYuKNRNhkEnTTPTzbEpzs
hhCvhTTmrOcUUA8lOH5lxd8V0oA2Q0f3Kf49ZX4HU+BcWNqX+bl64z0g2B6dJQRByVyIBmTsGfMc
mTO/ar6XTMZ2zKpKsn3c1IAm8dFF1zn1XSy6ZHeXTTnrfOfaEE0v/UiMgiYs7CKcEGB17+jMnu5x
+LLaOIf1dVUFBxwLqCUgtORLLPT9IxPONACFPX6GYSK0DMEH0ReFTzj1pQRJVDcyICh9LwCnUmc7
A96oFJ6//8R5DZeH6DHqjwarl/QhGrE8sJYmIs8VhwdpdCPEz6KyeRPxaI2bViP0OL27aHdsAlwl
K+8tlxv5hmrGmvcqGQiPSjAjBqJ+RwYzY1J4pzXAl3Z/D9GJoudUo+ZeOwD4VXQm/lqQocHo6tl5
aO4WxHXuxsybWB75QYWKbcYApN0pj/YPcfWsyTZivsSdtsL+sj2ordssc8r7Ixypt242iCY1C4N5
rjkw3LedX87JAN096wTsgADnNPTYnejTMGC0NYW8wBjx4tLLftvaUJMu8Z4a2DZaPUKJEPFuT062
zSObJHi7hVE7bWRjyj0rlWJZmSbt31I+OChyma02COiS/UCtkTSbmFyAzUvPYISo1GGCJmB/0TRf
HapJeX/RPa2LoMUjcA3Pq6LpjpfHdb/+iuSp37HrU6xykOyMtCF6jAcTuyTmcs6kGn+lgBeXLF0B
WeJWd33EE6S5mj41sYcVz6k5+VElLHIav4NJDPkZhPVfm6i2B7Ux4ta4JuqyA/ZkctDt9ZdAo3NU
4+5SJdf5Jim4O6Wwcbao8IhIpooe0h8g7T5xf6VpIa10jKksY9JBOIhKa3ufdENokF57gu2MeaHh
W+h12FdGsULLxWjY51dVWmCxJANpzdiquxk9cya3Pbn6BSnHpkyeLDLCeUUOk+nlDalUY8GIMu/i
8VPRQ+recMXDreTK8sxOyKz4ZZfQhB36pFbpr+BwFQJZIEI2OiV+Bjam/5HBa4BOty4NZHWzcI62
0HRwI2oqjr8XbEYdl4PDMNMEbmCA3avvv2Mp8okkL1Ijpj+eommQWH+tIXAz21htk0e3w8XhCLW2
VMmcdeLkRxX15ExKGjxOMP4owjJlRhnBf7yNlAO1a+17uRn9+frKfz5kjNVIPBEJ8Q4NeJxSWbY2
ZqXIAp+pTQ4KE7SmdtawYsNpx4zworjZJLO/bxkrEVfuhMCB29hWfwRcz7jX17JmvnULy8Ve+u8I
qcLXtUrP3fkvVAvwElr0uqTuIta2Hdyf5aBmMEtfQvsZm2Nu1tcpvFKNGO4kpg7BaFn/JYl+quag
VhbpR7unG2/qE8dm1WvHZWUXgdGz7x9uvqhcZEDTuOPOeGBs4TwFQgTsPZfrEdxQU+rDxWkZzaeO
Rfpn35UIszgOW5YcIaM53NsWiTwOmGHuZ0RoThTOolEVTy5GblvKCNStewHcyGyWvGD0KGRKe6Z2
SEw/XcUAvdtIAW2ZUlqkY4H8ftaAIUB2q+IMQ+mXC7NR+PPtww2tq88PJ8fiABVTJVfT71qGaPfQ
4F7t+ni1yuT2gXXbmChBz7E+lqHMKrZ1e5BP2H60al0Kp9slW2rRC33oMHvrrsTwUMraQCziJSvd
x8MVcawSlytkyNkh75v7P2PwCVuAUQ/0O7TtARBmisO0GEtOxMx+Gkr3LcHtmjzfTcOvHBeHstQQ
A2UljoigWpOnS/ku1z5KOWKAKROiIU4gIgRFbOvMNO8qADa0o9WuF7Ptc7Xxw0ndUwS0FHy7aj2M
1eZO32BpLfTmxDBNt2INNHO+GexQFx23aXU7kBfoPDfMn45q3msVDqzIq3YYNmc8L4rGHFa6WOP2
gTne1cIHOcWg3+eC6ipHfOovWO7tGb7sFdRrwb0AQ/Q2imTPvA46z5tSVav9ZxCcTMhuEvXoWnbM
F74Cyye8tizFCHcUyamOfw07zd2lLnsRevLVv5ghNQsxA7MEodcttXuvfv2sp+k8bxbcyI7CBs3a
cobXQSBBAv4aEbK3O5CqumgdXuwyYKcDS5uZLoA2/X3XkUAdD4fqkkzPvr7H44hcRkFJOjx/Cxvz
V0fSfzvVpH25eM1uztdS4S/UQPcu35h2CmazUNO+bD7to5qxO4WcZT6q0VUF7Z0xYhLXqlQuP1g6
JxeCVsYD/xJsZsuoQAqbH/ulkwhgfe+CpIAA8+zSWgOj2ngHI62DYfaJdlKF4HV0OfoiINnhadDu
e8cn0ZYQoCB5QCVj/DW01gjvkKI1SHA3crUzhK1j25AkO7dCj/+Y3jgTY9GmjdTGL4PkaYmjUXYu
e9IdTo5uMVtQsSTF71IqN4Vgws5i8vnrRji7pjGOc/NqbNaM/9mYdSGQ7QFhnUwdYlDrfRFZq0BR
2kBbehN2yAvX8a76z77Zdbu6agK9rTBPQotvdvYqWv38/xeARFoBbJ+XoWh3JKWfFx6VwtQbYl9B
IyBRO0qRT/vjRLXAmheyTCF+eZFW+NtONDhjCXipgWLBSyE+00qomttdu28aOdkm5y7KjQDzB6Dd
LhTtx8utN1YDo1F51q9AZ75Rugf1yR/64TVQMsv8+GPrEm5RA3m8hCM/wZTgEC/dy24MP1k24k28
e1bT67jR2MRRNs044CVeyuiPUk+JAmk6BCYq1TtG/Vb6Lpd78GZ8nswDb+xkgVN1PMe9+S99m9TD
bClaASCArXHC7cAF5nh/rWosDOYEerEUa/2nxeZYBAOrFoDgVr2foXnU96FwmuHgZ0bKa+gYBNMT
3/JLLK8I0WFU9oMyUdVKcZH8YQuUx99IiQNieOo9v3GZSgu0bzBL7IzkywuAbFb5W47bfB+aVqdz
TToLyudA0wcanR35JsQYMljzhLWlm0HemkoHoPDEmS4b9k3U49hiFtDG0+RJueBqFepap6Ztiewo
WAmVVUJVB1u9PFZACTiApj+doj3e4moYKy2mR64OLEQZWogMfoaf5Dal3A7F0ZsPknB6eDD/3c+0
Wv/rUzKDbgW4TDpws1U9dfImNrsc421mY3RUHvFNkJHiumhKT04g92xLsWe2MhoJbo5y00YhiDZP
53qJb0TSGiRnDKF285gdRLEWR3sYuD4KBOkrqUkRf0PwwZOpW/iH5X9WAyD4TOMVb78wC6O44jlZ
1BT6LZUnQ6skvTDWQq1UfeeFl6Y99BL8Vc72QiYs+aw46KwSCxrxbxv8cUCab/tmU9B5X3SsCvGb
JGXE+bijniWuAkKFFiR3oeQZ5Ms2P/D96QMO7L4xY7k8eZajPEXlEQ40q0kefotxml4D1jQqZBJn
ZgLYPWZR8P0MvdCtn9T9qaPzODdHbSnPtChvx0CpYMLHLA20QvJNkyXvcR7rxsNMm4dyEJnEmUWc
Xm5B4a4nyy7+ps/Mnk9FYPkJ5Ykt667qZEtAaLc+h9iReJJBwPRTKzpuQWwZfBwbygmD4+ABq3sV
1BdV9ysdph+mtLjU8UCo6eaDVdn+bWJVk/voGmQ44bsTf6Z86q1Wo9VYniE0hijWO3WR/ZSQX3vK
7SNSUQqfas5zK/d7c10tVf/H+xeFqJ+PF8cO8tWMceu2hyL/qExuBPh0vRvCVVsS8FPWuV5UgLrk
Cx6+1iTr/BJ/CqbCS6IwPCvPgMyIbz4HQNnncpfC/maoCYLsd6RnuQNscr0XE/eQ13tc6mV3K/dy
sSR748xFA/VUKRBkUYm8HytlPP1ezPb8E4EcivtJd0bXd4zB2nsk1wQQyi46Qr+0Qr5NTzl1Gq0s
NI3KbgzG85yWPgF/Y59Ghd8rlN3GjQ1Zx7WVrAxB+u9/Q7dtHJ2WRmE4VePJij/2AESnK9SbqKGK
GM6921nbGcorF0JIvKsbjPUGhdmcfjFBMUpTl3o9+6Xa8BeAOg0Mugi3Uqze08T3VMNM4Ptz+PAY
Qek8wLr3xs/cVppdGt18r03OEmUFwgWBQRgS/Ry7ODVPGdQJQ8H5rTncmPaYRCdXsmGqe1pcPFTu
8rJW/s621TTphtSic9zBOcENvn1mT2nGV/DOwxXxuEe8k6Hdm9Jxgro0xz/ZvTef9b49uzhonY2h
s79mKUTC8BuWFT0U/NuR86J/xkhpX6HaWclh5qBj1rPSureVV4ewm5SAn1UU6Jr2vKVmJ+7Lj1aj
ffROBD4yYge/2XtKyqxULDyMgaqfjZ8RsD9uxaflxVSZIF29MtNZVkQNNunynHuxwwE9FUYlPHtt
XtECDn16U/emG5wdBHrvUwqktP64csGyG74J1PwZO0Xg8icteowlnEG3akaMtFZG+DBAxMDeHzMs
MDsUdQ8dB3Ez8CibzFneT+87rvSN81n3UsgvpdwU+W6eNo37gedoq0cw4aTZIuiVcWdLOcvCBhoH
u/Ae1DG+jxwB7EkVIgkPqFnCsFwnA8eIeK/Hv5/VP9Zs+asEHy/0ncERmK2kpkZyw577PcAb1q1a
811H6scjyg23QjihS/Z8m5serxKMO2+R77KHXXhXIc8MqTIMqK7xl+ceKxJV1mZk3zi+HjpE/N+Q
CsOy8yrMcpREeP8e6JXyTrr4CPqruULwqn7XgcDKtAajryhgcLpRn7XDLvHntw/XpSxqFeltwGLm
7SMgIoa/I48sDUoCf9C7HcUpXCf97Z12LJI3NnSA4Clh2nbE1YQPhrS3ucXNplw/Yaa0fRMpxpvD
IHzmQpMdNGahVhDLlf/1XNqGusRMYCTiSyGgJoGqSrXiroIOxs2I08sqHRY9yJUrpfiBKpBA+k5U
qYQJg01sy8D3ziag6zK980QT9c143o/L5FRd+4CCxTs6KYLpoj+COK1ZuPJqw7UUT4+uxIOMRqSd
KGbUu3IzNKbo63mYsfSp82Ev+chB8onVostCq9pBI+chjJmG0SSB8FlBGT8gy2aRvtzDSvyB8u6N
4Q22WNgO3Nxl71z2AoHBnRoBMuAU27U9yMRzJ0+tL0VJTuJ21lEpfJH9W7WcH8GY3PNAtov3IAnJ
dL+PeE+iImXwExCKsm/Zn2eE2HS3Ro55ef4hVjmQw47SDs/Ueym1p3anRA3YWLNzOSSyw+1yY4S8
80qSuFoIaAgZPXTg5J6/rbCnVkYnF1bdw8hGt37Xc4F4Sciuwd+HNWOTGBvZxjgi2GlMyw4UnV1G
2/WJ7KvAisC3lzhDdvuHUnUL4WGPy8/RiPDU+O8pJP/pujTJ4b+0LjtUrDi39SJYp9g2WgZsj+pG
digbbCp9u98Zvpuo0C2Mqv9bcbzTsWGFGt3VrCDKqLnxrWdXqcOr44aNY1ByRDo1kF0VoqWYp58e
DQfvur8aWTdX61gc2S1yhR1U6GeL5iMsYluMhY2cLzAp1sAiAqvs+NixH2mob1e2vdRvN/7K12HI
4PVKatKGYxCUEryUYWSga7AnV2T1lk1nSmaoL3Yptgu+ymLJHMgoDwm0gULjmJR2YilaV0abELso
o+TYiFoI9vtomH001/mwD/7+BdJZQYWpP108dx3heMF7B07dgtVbaoinNxD+h8svqRXwrby3xkeC
akuOk8z2jE40f6wmhJTZ+so2ki6PScmvulVgHq9rIukiSHZp7sU8D37/MasZ0bAfUqUIJOGGgz2L
IE8pPVUyXqoYNbEpWxqAYFJhsRTt8Saf8LaDPenFMuDFgeDgK5WU+q1z7oNLd6TIH3W8nm7MXVSa
jh2KOgIvWbsmusNXjWwVCdiBc7L2iaz1rklJqXqFUwP6AQwrVFF8FzQsipYz1nkEcdcoqgJLLgDB
XqSesHhtL2Xfy+7LBZKHdRTSVtO9VPxRwnhGkkqG/7XkJj/QYIVJmj1RwJN+7RXA/+9NVqaaH2pu
0IWw30hGSsVxjCs1kgHz6ueixlc3bXJxM5BYk8gvMvW4RAK+iS+h430N5+EA7mGDkg5h5d/hS04X
z/OhXveL2xMI3ZvSoINi+TM/f2UvJAOupJve2pclrYqMzZmSr/i4DENtXYLpLH5P15eGX2hb0a23
L7hFxtLDzynz553dig+/1ZcJ5GjIU/+lmOTRfqvTaeNpseWRBVioqvbTuhp3QaKDcAdQelLoWjJa
PhJHVZ0gpWZEMM+Bd8ZB8oX3eNfANdYis6Ort00kYR8eJQFeYgHloLUKMQ9+X7stH5haKnuE+cNJ
LV0LfoD1J9T3zr+bnO6bgylMdHeWJ1W5YBhkwu7jYNotBZhU+Mq4TeT0X6y04fQFhzWin6I7fgqw
Y2XK2UuprEDy+UUdYwS4HPW7/lv+wRY0XCE66j7UBpX1Sa+ioDaERRCJ7MarRr09a13P2/JXv4ln
vgCWCK61JLztRCv7XGpvh9GFYjMu+3T4axwxTei7HYHe7vApmUMDHpFDQZTZ9+QcpO0otU6dBdiq
6RFB1hpxv076+v/nXlqWduaaAA0ofe4YIDr9RrPuIaUch+NTqtKNXoHFt1F1TRCYrzyGfqbcozNO
2K0RKoCNrRmijMmKbsGMqJodoRrmUPAI5r3ASr/yvbMsrp6u5StGyD8gj122JPce38uTSGQOnZYn
yM6aeeFssxbC8pfwpSziTU4FYHvxG2aQiOCY5QTTv7vMjA6kAagAxT5viuAaDWOyE0o2MYIJX6gs
4eeFmuNRmbNJNMG0N8c7SYoy5blSEaySo9EvtDosE9xYuJyzrez+slzR33HTYknAWgNYaJGQZLx0
0HW7GhnAh1dGZ3n5a3LENiuHgfFwDeDVSgU/bCWEMfBcJk5PvEKQpEUcCD23Omeb60aWX2m+3Nve
xgdM/3EOY3kJr2SpiALqMtKHHdw1u8NZ7BG3OIQZ4awP11dPDXCKAxXNLTI8N/Az72WdWtjtFPUT
wXvZhqfxc22UMpLTnI2n26RBaKm7V/1mRc0joRWuRfuD09nFNjN8bJQ3025BJxMfn89ri3NYCQxh
b/XD9VC0PDpoZTJFVMvLnU24qhwiNK22qwb6sB4eSc4lwdMvJ3lJy8tUs01yC1R0PBDgFKz7/pj9
FWTcAq+1/c1SHZjk8lcO6I9SgepuC9BejZtgmofBjuHzc0bogwKBWETjWDWlGtlNXFRIJi8n4SMi
Lec8MxMtLnqg0OWz3k+ZjFHY7HRH3pcVesJ3tUo+czp1QT/bTcSQAO9+RiAi8A86Y7wwS/I89WGj
WvW81dB1aVF5b7IhFWy0P0Z/JkLcCptGZ9qbqRITujS+e0cOTJPA02I+JSCSa39AwvbOWadQH60q
hPBkUVnh4sg4Enpwf7nYoeweT6CVjNSR24qZYhzvXHICSRX9Ix+CzISZ4yQqeKnobrgtgo5Ongj3
iSFCbeQWLjoLyegfFeoxiN9s3Fbq02ZWAteMaysKngXRMJXmYrW6k39KPT97JJGVqgJudIhMm/1b
g0Kw0GZjRIsQnYNTUnqZ2/IMhyXb6WePgFrhOWDrcakB49LDYUE8JpxfN7teq11m/vGpEtN15llO
YjPHXA7aGgd1yIo0Lq97yxC+D5+UZziUuO1BTFRcEGTjseuTVbCfuGQGV8duyh9rL2Sp1gOg+1Wf
ThO/mxyDuUpwAxXeTcnKb6GmLkSmCixvam0NyLql2YpQb/FW/gWuTaqYk6aR/sXtNpL+plJfrGQ7
sP9l9C9jOPGOcBP9dUTa5SprTju4XEqfS34Xh4M9fa/M9BqWL1piUhdYyRbJg1pYOBmE8K3GEgu3
T4ZZrE1/Fmj6f9fEuDo59vJK+v+g6C4B9ISWAYBNpgmGsLjr7wMQuNu64qMpEdyh6UntImfbp+nH
UeL20iPi5tbovMA1FUFwzglwSYuR81mWBXFzMYOOSe39fmxAUaLsA4p4aFAy2TUxmBl3cQAEclRM
U8TFsSq4tINp42S9QqCIUjI1pGV994db/eR02yDLd+KN0F10/o7ti5FaPzqRewYzKmAHCFic0iQd
4i9Blg3daHIuJhG4Cd4GwbxT2Jh0m40F7wJVGPUdcHMm4sDbiV4CIq0tVMvhZDmCvdUqm8nUjQWj
aj6i0Wg79j71rw+WhICvkBk4u5JYThVF3ZvCr40FX+S7v31pJUCZ5pZMxKyA+vQs6/LIJ+6b3GC9
wTLFwA25r2WdJH0rt14dee2aAkjjDFT8XyZ2+OQRBq5tFyFHWAf44WQ+FKWlQEx0S/GdFhekT9m9
MgB57A9GBxvqi7R3OokZFC5L2ZACiMd+J2x4o2hiCrPjbTf9RwabdCVNO5olq/yjVFwLj7FoHXwg
Jg/5hOJKY7CgWApM0yk49kpGjHZkf9HiKg10DiEZ7DMr/FmQrEgzkYShVThRDV63jHK59mz0WArQ
5WV483vaECjeadEB7JDvysw4MGib06r4v/iwuQbD8JEGZyMuiqrOfXZpCWYOYj8ka3BiBJo4eWlT
75S1YMJCBfpegU6jl2CgbkF7KrDneCMmjEhgqZ21TjbDUFksIWbI5AIC6L/Z1XbmM1j0OEhuLEf5
AiL2ukzY99JktqrVCcT05dTsl8htpBWozYWmxuOv0l+WUQvlW4RkjCooArd7WCusKBg65iMCKvZm
xxaFCy6wG5doM4+k/aenRNlxTj9iXvLqM0wd32jalBnwESLlXsd/co+Uqs/dD6AsNM5q0V4sLqy1
yKRU21VSF7iVZ/Q4ALBWlZuz/snpDAmJfgjvojURRQ3Q1cRJDib70ZsAjUwYaDrBxaxLYEi941er
pTrxJPDfDb8VbrlRIhQE1SbHcnP4fG/se57ej66Nh0e0U0HyVRC7LTks35qsZUR3hLxW76p0OjZA
niEwnFYOdgrGsjrpXvDWafN5b8mGw2y6UtrY9U6RkhoArGlOxVJuCoc9hV+Xqx7dBJ5n8QZymtxT
wjMRxN/SS/n91SWU+U/kHhSLidAMRlAVIIgtHy+/Np2yxaYEqQPOgb/6FiNawmyn98j4VkctpktV
qmS7+JZ0gBVXajIwguYfAhuTLg4l6jg6Xa4fdNhutEKa5DgOzh9PnHewIbONuUE3dSjuD90LLEgC
kjIVBRJNVSj0TCg74B4bXl3XSHz5PokeectyyI9nbSTSX6mo1Amlb7Iek5kpAcmlEY7hs+XnCL7Q
HLZSn/sNadGCqgllsnC51ty/K5ysemAYmssNkXv1q15djeroeCgqGXA56bGYzQFSyeYqwoRAs9KJ
Q6Qv+aO/MaIk02oTRFfIkVbjrcziJLb+OtWrPmP4WVQLB2mE0EEM4zqZApIVi493ZBEM3DgjC4MT
ngipfB106roADZ6SkkXAjkrjtN/1DSK5drOkxDneF5iX8y7QkbjYtPDva01AJWDEEQGoZ9rSFDO9
Fde/zuWOcCBUcEuzX/0Snbdjy2MS5gGlu/tDFeylSzIzaKxdFTbSdyWhMzjJQq3TmU0T8G/XL+YC
CxJwimnYTXg5FC0rL+VpSNqmlOW+8cC7qrb5Ojez17g+GowdAhI5X8FUPrYoGFWyRQOcLucfcKYl
5pm+GPoOl2qCPpRviWaHPWntxdlgdSAQzLBApHyaCN0qNi59d2BC4MzqHfvoVE/eEM0PAeu3xXMV
gaJFOf4D+HtY4sLTfuwYt4y+5xNcWGpkcfqpL/FJ8RHu1yfvJ7ESOyjRB40U0PcBJbKtR4bNLQza
I4usNpCr9Pay/PxJ/yElcDP4t/r4+A7yay+sOG2CymP/Zhj5NgaHPVR/xfwl9CU1t4xtC/ZoUrL/
rSaa7DYun3wMeS8vDTKAcYm8DWa4fymwWeW5UF7G9yVrqgp6iAXjm1YX8gg78m5KC07NLrqQoWii
YJNVQpmFn678HUiuKbUlA0ieWopICb9PLQvQ/amsfIHeYvQn3dNFdxBGkgkZyFU4viFg2st67FBU
U7/jbqEMrG99Vee+RJ4egS60rZuRa6oxuDhYwt9lOusQBVKes/0YK6xtgzJa4sNLoCINw+X3UKXq
QjwsRfh80bvjMPZ4VtcpAWjeMqz/5TW8YSkl7BnlyIteertCeiynMGP18j2DBcpQvMZCp0XhfqVz
35hHhToGzEhp/fqUT8PUaL2tTGEqj5DRp9G2aZK5Tu24rFZYK60pT8f7elbInfiFfurx6UelWVHX
9i94OYfqZ8xrNyaDdMXS6Nn4ySX6pYeSSIFju31VSde9Maaq96OG8ERpMZ67cs+cpOo5L+ZxFXYz
Rk4QLGYaFWCP1p//fWhk61o+EwhtPc/x81Nwvwpdjt6Tx71SKqxHfWXhVG+zwnPkMfIk4I3W55YI
3SXB4f+qRVTEKoehVa34+1E8GP897q/T6AYf4mqZyQ8oZoDwh8CvYDrqrDSeBhmxWiUZ7JdcsCS7
NAHxNHnlGVxCmYqVWLv4PbvQoXkX2nTbnR2ve/GjZYKIx61nTGOiaVMfRkB1CtXc2q77h7YjplnO
1emtYspWtYYF79gsF43rC2pcbV7gY3wHA/zg08fJQPyIhK8earmye6O3VZoZ+pT/kxdolR2ow1WA
+/5O/1at4v6ptRaStO5zl5A96aX828j96JSKELnnSisZglE2xQV2fBWGHscNe9VgAY26yEEyAIFt
kvl9+kuoTkRpRnkgwKgEcL5CTAzf9aaqN9NlU/xjxmJX7QK7DSRDQbJ2jkjAtsGBEpy5Zjsay2CA
kk/H9AG4zhC3Iq2ZPHBg4PFmI2uBeUGSKpIN8GR4loiuD+S9zSkHGWgTWfl9xfyJ/vGhNZVa75dR
6fP1bt+ra63XIQaRNZRR/lNYYnP1NSGbFnQLLOGFsdcnDHRt50mxGJI+3hid67FV/Zg0YqtGFoVj
XNMirDpUicMveL/iXgx45FVoAuaF4cvrfaudFPfbkUJbGX34fE5GP3Fb8cdviqB3XCq1WKe/1arL
6HMLMpiueKEiI3g+OZidWvf1yr/BDs7+JM0t2AdJHnC8wkrPjb2qb2lKU46avpi4CPZIuqHkLRwg
30/I7jJdekfSYS78RsekxOFmRRcyYOdQTj8z6K082dfoIJdl0jaPJ9Rs/YuwfNg36Z5xI1aFLAwr
k0oXxmqdufskOFHccslAtVMej6L5EfwCioWCWMKuZBqIH+fyomdvIy1t+KSCNOG7Dbkt5OXRF0dO
KnQUJqQOwicxHQDqTkUF8Wid5Cs7fS17ObmHbQkbpvdE1iXrgj9qcFepQeQg+97VYS+n+6lxBfB8
XVfH3JcegLlaDkk2xDfFK+E6gY2QlpqG30WZXtBzqPyYzlocm5HqHOTPIzrDt2Zarlu/R1trXVV8
JX/KZzshX1IhLMn1do2fIpR/evRU/jdyCGQ5LS0fPPRS4Mr3O+UiZdrqWPkJD5OIYQ1BrbuqNme1
lqz4ksybWLSXFFH3XkqE/Qf85E8vC9UVVaOjYncj7qMudV5iWdb6P9/UaWinZEXPh3o2bvKv4n1w
x5wyaalL0n75JepSvnyppaAQGexsUu6hv6bQ9qlSHvUySE5ZTJZEdeagV/wa+CdLQGp1/LYPw/9k
mZJSjJwudZmQz2qgsn56BIsHPH6u6Q9M60qOtCKwnCI5gky1xIX7lbJ11RLVhw71WNhhENhC8k0L
ZERLUZvHOy1Gijksz/iDNPa4c2r2IvC4ECtSeFtiuNfnaTowd0KxIgR5cOX8Z/dXTRmraG0qKVVC
5GeNhCjSZ/JH+afhVZ2c85Ujh4a+bE9i7Xi9FrfpOJ1NkFcRxQvCbPZiEgUIbSvY3oyi4BPbrqxw
JbeBwUEkeTKskL6lbkMZZoxMpBQYH/O+BL6j1hrPiGXMFlXiFXSrYbdmvJ8bGiMs125C5l3+53to
7wpV5KrIycOunHDRd5rQDMor3k3LVL1amlEhHZZelivznHayTNq3MxxUuAAZOnjmA9cvTBzRGaLf
65ZYxWarS+aCs9bptuxHUl1VwajIr4g6ZYH63KFjDmL634wttCDhx/yZazC3Pko90EskN0VtKvov
Oa07BPhjQbXSO4MT2asTMdBYyvTfTSVFmh3u7peW2rlvQa2db/0Mom4vwYNz+J1GvRpaYPQ/f2fg
RgtcMmRzU+8zzv/05KkMeN3Ngd7fDT+HRK9qXiRxRcmp8a3wC64dxF4jrABY0tJjEtcu6225YTn9
kMVpVMc68qebXDUE3DPEogfLvdoCs9pwc3/WJWAKiYhnQzF087LlXuOHIUR2BTXN1iJBgDzZ35yY
N1O4UqzKWYJChTb2KFpUXYdYZieTmv68htQ0vCNPQMXMuoV239OUs/3IXsBHJDOOzafHw7U+g+ca
Au68lviN5qYLYQ5xmFl3VI5KyJYiVcOaWRcbPfUlRuL5IWABxV0oBX5SZNaXDbjicEq9f6IzLvwV
CwikT37MjSeKaRC4t8kjy7GaOTvILdinC0761JHkqsIdcE5Z5if3fxLPBFb6rhPPyDdlRHqj5ORO
+pjrbIBYJ44j9aoDZXnOoNWhS2HrBgJIT/0x1b0olvhDaZ9zVXKFbrtvNHr8FPOdWZwPQaTDKp0q
E8510/UNTbWZ8MCGREeT1WVxR0I0uZmObO2oYPWuiIjbBYQF1X834g5SPwO+Rk+MRpuQEUIzsw7G
WFvR+mww/2O3oVEgeSwhK8BG7EZu1ZXZ78uN2M8bx+k1SXI95b1XcaDDV7XFX43du5rbbxRB29lZ
niVwLybWowrOg+Kk0kDZLIxbIfkpGzKLDzT2lumnn+zG7uGe78X7gyPBxFNPrRrcuJLazUE3bym0
Q0B6JKBjczKQys4BP1khiy9HFkOP3tpH4zlk9F2x0O88MkOmXjfvdAAoeiXsWfrCRJWKrLv4F+jV
0yMcxB0KIuXORyilIdap4sy6mDOHvOADj1LDNG8mvBE7h+bwSMFDphVKzhP5q9J4AieP6S2JuAda
CXG78EcwPAsW6QUE59OCV/IsfnZD6z9wkGX5A3kTyqZUI1dNmhjM/VomNrNZRVS01DuYjVgemw6X
kLujwGfghINSmyqBJMqXXlUYIdBRtHcM4BkzGiMWenPNFikS2iA0b3VUKYcxb2ezBHAdwNLTdKP3
lvZupRLFIY9AfEoE5tMzrUg8S2h3JKiRy17ZigY5XsmDJpmwvQ8hnres3h0ylYc5ZrGj6i9KNC7T
GqX53Vwha7Q8xtiTOFlt+fhhboxs5P3Aho2zZtYAOhoqfXayFlP0KTnxK+bN/M3CO81OQdYVuvX6
xt3z6acvatynDNQQOH1SOwOnZu2ljUI13fW32oj3vJrJovUGsAdEZcP/oQFJspfbIDBzwgv0TGWk
iawNDPJTEhGN6nuW11UsaPp/fTHMFju3eZZoBOKrljwA2iPQDVzsnCmwE3ldMYlZp+jVRQCpXnTh
cYsv0yP0mVuntyvlje2ncDRIpfY3caCoJ6L5ULLZrEHrTLP0H+WddU/FMQs6aRin3TvfQ8hQR2zd
MJ4ZdFLG8EP+X3IYNnTVxW6esg+2KTBCw0OH/X+9eXGRhkhVJEcOupkiHBJjBJ7wVcXOatqLxvU8
Jzn49xSsXKeYiKpll5C4lGo03JdaTpWsvEwvxXQyNKoiV8JIWYSo69lswxchfddQMheNJOkX6e6C
q+JLJhDMw20pxXZ1rPYMgjKJBM1TrU8OdjPLg8cCsGPvH/taq9Y4hvAS4jL/XMf0K8j9AULKRGpO
GsepktOnUgnFhn7DiKmXU73ziW3Ee/iVOUPXEAO+xEeSGA+0DfpqXxhz+8Js8E1p5S95gRx1Bi8p
QeJaQxvcf4+LbADrhjkJzotzAOFybbd5hZ2hH772jtbe3juMoOsQafBFyYzK08uEq8HjMWYLGStk
q+D5YIIPvqTFJJOj6/oZkmokV0x3w5nJZEpkzWvW/ZiJo9oJ9wSYlGFD7Uw53UxsXuGjCTFCLiDh
qFiqWVbwKL+Um3je6ZdOFiwug5ZxhWRIZwt1r7ekAvB6vTKxndx5B5k44pyfwjGqKXmjXW4brzsn
wZbW0T7sIdixaJIYvYukPNb9pIHnfxJjR9vhPlK9ilcWo8hHS7TxMM5pTh5RPyHQ3cR+BI2hbd06
oLp2o5KIDfjSR2KUn+48cRfn8w+elo90DHyci9GglJfUA1S5LkKGX+KZox302ArpwrwSN+e85d4g
E5QM2hJyIupMc6mBFlMed+lZIIID1Ezd/xjdno5dTEybAmn+FA1Kp3/ru8me3zPvOGWEeh63zkRf
pEorqOzJdpKOFyACEIoXNJqiXn58/0X12j3PtNIL3p+TfdzgxKWt7P4ojWba0UteOB8AwKb2jEwO
aWI7lRaXb6UD1yxG2pLdXX9if+XDhJb4kgSNkvKU39FotwMUo0AY46gta4VF+j3O2wDyFiIiLsr1
B+JlPbFpvvBVd2EpRt0dbUt/A6ih1sB4MfpBP1ilZTCbLUj+Db6xml6Yeq7zZerQgxN85MhOlDAs
FF1b6/4Zc4zJIJxfvpVhcidAk3HjfnzKGjFCFyUL/IxI8EOw0p3tFKvarenXv6hb+CeyKC1hMPgj
ezh3iStDFim5J9AyrC+uHQtArlfCTVDQcqmALxf2Pr5rLGE81YI3ovVAPU3VDfFT1uso+HqMkwM6
Nb1d3sj1WLiaIsRtNVTORi6Cd83FoL+W1nIuQqJZ9vn/0P1zw3+p3bB2A+65znHB/IIKn42QYf4x
kwq0CSJx9AoCGfg49LkpNC7ggeaAZL9Hxc7YnlpGWYkcuSo+8/KKetNGXceYUwEl8KsXida6Yzdu
MUp7ewY5DQ0m4TN7AAvP2wgWObe7xy42sWG7orySDPiY1vC3L/E1R/vO/rw3/FQ9adGHi/apeNf2
TVNl+7bj8r9jjkeXye4yHSUEIBM3dw/N6BbYhj2LcyhwfiMx+nmJTR0Z2gBEqhxPYVm9lGXbl7KR
VV9aIfp3OMqGtKV0hmA+yPTfdovyXJQjYJWxauQbcfvZTteR6VA3QOYwnINmVqiawc9QRvRTQolA
nqjwG2NVm2qLn4ldpp7EVm941dfm5qlzkizM6gKp3hB3BZ3yOSfup7CCGXmAU7U2SKqfdeg/6uuc
cgpo8HD2+6Ow/GsAqjPLmxpWCjZDtmDd6KAzfGawaPl5fh3zdn5wmnuahRQFmppsVduKxEglmMb+
CB0wLse+kk65YpXQsns3GJsIfWfPSWbmT7JtA7uy0T2/h5Z+SvSj5K3fo7ljAwSr+eCZooG2g4Mj
C+2IFZJpLLdunIbY8gqD9P0NlFUikyPU6IMsgQR0yQrzg1012WrPadiO5jv8ezUzA+O7Dl3+tWpH
eoud/aF+197ACQ6vZR+InCcKwbFWHaoCX8ycF+aGYNXa9WjdYqgi5oq7PRdDOp7vV0pjvDD9F8ur
KN7JSg+fSpsJ/NyoagO+LBMS2pM8DZoiceyXAON1usymgX+I0ZoiS8SsaACspMsbJglUA5v1IDYy
HmpvHOPHTpFuF05OByWmbCG/af7h2+Z45h8St5I1iitN4qupw59bEx1C2WMWEvcgiM75TjJlSQME
bPNHsuf4ZTSulpjv3xqBKe0I6jH6gj/9hn4y9bE+sArPf2nYuoyP/0VPWpFxo5cVeDU5b5HR+VlG
XGcaikYTsEwjPqW8yySLYfi+Y/oTih6wiVZcOYhBpB3riUl7f6/Ju2EEoEjGnJLkqhHD55XT8G20
oSI3tTIZ+9H6HKlsYuyGdXfeCjLoOBjRAaYF5bLmHSv3ZLOWEZx6eDoLCYGZGsXDykYS/Gzcashf
p5wvVjGXIGzbR515ebQckjo25I/F28PSb/Xy1678jbCIxUzNIownRXTAp4hiJlEyr9LIe8KyfQu0
GexVJbXe5KE+updqIJXCdsXUFGZTPsOUcb5czq9y/Ro3EHeHhWlxGQNzk4qCins+aOv/XesL2mh0
A5SfKJSZ/QIQRgubU3VwI0RX7YVDe5eAKcHSefajaCM1VPWBX6d8nt9C9C4H3Fq7SwvS/kd9pZmJ
gb6HBPybnKYCpcdTTOfKWXkYizZvJQXtYD3zcLrznOvUhT9oOOi8Ga98kGXW2axtDkp29+hMrz0e
eJX/jXPZ84nWsQv1Cr+APH+904W42WB8+PfsrBDSX9I5wXZeIij5I1MQlUwUcOJDRAkTIClBLIvu
RnJuUBPnF5vC3dad1nRFMWbxRp9UVdJKCYhOyOHuxhTre7fxXSR7yMnYhiIsCZz240el6hNMcTlV
FpZie0W0m23Dj83gbgPDkBRyWimuH8e1tIkTIYSptAAHADu7JNKqggR6bKTBj2dBKgdJuDeh2rEf
QFsPPuWO8yEUKDHNsaLYeqVZbYvJp0IM2ZS5/BqeCJlUs69F5RNkR3VRQPTTFYhrnyv3brlwYBBI
wO6hiishUv349Hv44Okeguh5hO7uwMSgUQKjieNzMVL8PUQWoKOZEUnOk5DjU6GkdqjWjhK+b6TF
Ba4huc+QKZI5et3g9vH+ARGauJgb/cSCVGAOR3a6IDsAwBwDZ5ivmSs4y2JsPhBKML2fEVT61Ltb
4A3hzwddgDIOQZFEM5P+F+ow8/+kPw6QN/cysz5B3RQ+PGdWvPaLU5yZTUNDX46FrodG03MxGfJX
Wli+NNKq7IH48gk20UghgiUiuQmUY2SDmBVgtXVjQCWw6VQVraI7ZV+GkeHVCAy45WanIwIGCMi/
BStysYVHmmWiSTvZVwNUD0JKQHbnkSyqniuDYW5QZDupVYAwHT0nkI//3zn3i9BLJ50Aw9+jRaYM
m1OyTn8frwhgBym6TrDaVgstUtcicz9ugT/0bXRgbOL6U38LybiA6sApMb9D8ROT1/ZPG9pnzGgQ
07g/X4lzIJzU6juHy2MnuqgsvOfHZkSpVWeKp3/6vHTKpC3w2/8XfEnP1ja5zb/nuqzPErRE0Tuk
cTlyBeXY1wXzSOit3/Tla6K9K7aKqapx82o2MUVxgYtQlPc/ZSiUxHqbP5hDkbA7wJ9n3InegGMz
JsNe8HYp0KbHSmR2Lo3V4BkEBbR/1BUvtlbfTmcD6WAyREHO4utftl0Ys3f1sR4cqwquOZK4WTA5
U1m2Jm5zpRT3eoWqfpSxZce1BlARyPjua9K183pi/tdQ2uFZ2mh6mtho/I7n0cLwAUhwdt7Rn8Pe
f3Fuq/4bqm2+eKqF2MMcIheFn0PnhkQdkv83H7Ceq6vxHXYbgpDmGGrMrbg5btLBMiYwWfWdaXbS
Kq/bjZbyk51GV6SYpL+4KZeNX4wxn1/TGssRK+G9V8mjUdm8acnpbe0wGYkDYAV0VA5lBhPR7iKz
an9fzVC1igJZ6eNOBnZepXpB8St0cQYUKHEeOw/ZR4DBthJdI0seBCXGDaJdopcgpBgoYp9AaQXe
d8lpZp7BBwaYNDgfn7zRqYJgQmjD4TNbqbZz60qXu3M6VlUFlygdC5TFYHa2c0RfuWrbEqOwN2G0
HNqjfF7PW35IO0Ej4u4VgqTT1RzY9dSn5QbqpYSBanutxsPQGM8b9wpO2AAGZTKQRVfJa8+atTMI
qArhde7peSGUhhC666Ov9HkZv75IrllVjqHGKnTs8qKPKb/PNoXUdkte/BNHPJayCHLEZqtAmy5G
3givumkqOvSNx9VVSWrKRyG6yiYN2NMxtQuWVm0oGPrK9x5+Zqab+oikYa2PQKM5gVMj24OcyzXE
5KLdaJXAdY25g3KcWP1ns/T7nz2txJyBzyKunv0mb9pkZWie2ZlxXvX6E/i1dKafDicqroQhbBy7
GCQ+MiAipa3keYBmD9/572Jyu/z4BRYmY1cvBDcq+sI/pawLRcgbTqGbrXTyQmmL9YIPW5ejmH4k
asIMs4H/kInNXlKrae55jQmAYcmihjsAmDp1zwRq8wxDRXfhlYlVRFf+7VJyrqBiF3iRHqESpAg0
eTqd3wLBIH+oVdC3dTJ83uefXzdpF6j/4w7nbMiW1NXeqWySHvcHWo0ozymoqXb7HjdG2voHeKUt
+LGlOMwQa1u8xaXEBkOoy9MK5IS0HpxbqICGpjmWU5hPiY4tGVWEuVSp/Q0rDOFbV5KbWu4dCLe6
l/Q32ZtA+CAoQaGT1pzdhwtjpT3QUv+LflnCtK/YO60fS+wtvoWhzBCcsOg+hr1+0m2a6PN4ETR6
5e41qocFbL7C9rIRDc75oWMXZuOFfoJK6MUKsbNSw81wnm6c2ahwd2aP0a10fRnALsvlZwMEOFEW
1ut4cNy8U1885bwdOjec8s55K2i/AmrlyxN3dEyZovdvb8CSgoy1kjnMS8cwBgDjKlZ+V784DOJi
ufmH61s9a3qZult2vAFZkfiOSgv9aq/kh+otcybLi2X3Kw5BKjtO6x9qQKrIeePuwlOf0nQAHHUK
GXkAW6RB3TS/Ty0/pr8LK7KOS09h/ExK875Dsb5CzErKmcy1bb1AUzRkfa2ox0t5sCR3fbnoIYhY
7pHYUEJ2ul1Xg8akkMJBeoAVbomxaRwQ7aQWAPRkE8znmma/Jh1PzlemqFq+fT5ZtRNTabjNCqSV
JCcGWJJeo7vlPD3qIn3hik+hQZWKaH6M8XRXYyhWkM01FY6rGu4HT39uT+xWtCWT1D97gTzYg2wD
w/e4AiIzXIh43Q3QRbFCkHbxc54MFVfTr0crqEMUPgLB0R/Sq30hZ3Xy4jTMx1Lfk+XD/Q2Yyvfd
R4fVTz/JCKv2ddPcOAJ3TRtfQWJqGwc/LSUEYrzpETUvY81j0krhJDk7ZxY8lib4D6MaRxqbncYo
RxhmAKGyOgNDUcO72aeSOdVqR4rNaiF+brpej3cjhWQMNyST2pWIg8JMl8Ujb2zVhclh40g0BV/h
4i4f2aBKzm8rm6yJOxH9gAwuMT6x5J1+oY3pcI8GbQ3nDpfrTcDPnDO8t+4QFvfpH3rm+bIq6C7j
WQEgc0bbuIG8d2QjWKpT82I7cSC632ObSGbxgM0diEiV/c9L8z/aDbFlzYswQWml1XOczRvb9Iiz
eTm1xb7g/tc3wf5gMKBeKJthvDM9c22nT8Ahjbe9C7geYLG5SWlYALufPTMtAgpLKNN/uQopFDxC
wQExJa5gHl0msjitE7ki8kSSOOd4vcVLnhOx0DB2dz2XaigAltLLbYyoydwXdvc9OXzO4Jtzj5yI
od6gKLotEVWyTRyCo0TSxhxLUUl7nasvXKeaU0E/rAZHDks8933OKzULChBufATTs7edLd7LDyq/
r/I0wtuoHkyO3rzuYQVpLbXvtSgu0k82pdz30UWu4fqBvf7Pucipe04RqhX4mzJoBklVLPN5biI+
4f+5gWgxqcvIS0jh6V6B1Omuf6mFm06TVJbl7FvzU3rT9QtNBRW63C9wiHh23FPdk0jkXNA+JKyo
1KFzALvkNu1OutF2x+okPQV8l5Hm4PCX2lkkM7aOZe4DLwpYC9/+m2GNzJlB6T9TzCVcUxJRr2gx
LEWtYJAN1rnW1H2kFnhosAem3fm51adHlsZ2hTCpBZLZZKHIdJcXCR35nL0mmXD6IHOI+/6Jpzfs
dwsisFxOz3XIqwr3z0XyhCqgxtpDUGbcktgMrd6ddLRznD8frAP7Nmq0rHjOVQ/kT3TN7MQcDtMX
e2Jr/0mBSY5P9W1LndXIP6tqAezUQDyIauxGrek6bP1ryLtJcjFY82K6LeBvnmDsXzFv1eIHhQxV
gdEYOyPxSyIIG5G5+OA2wREOjduq4KPhqG5KY/sfl4ubJRdSCkbBLOmyOHNiiq7WsyOXe83tFsAP
o4mt/7c2aIHlPr6mSXdfnWDESr7kmn1jHzkCnxbDuKe5Th2jFDFG4YW7j8X/XSFkcMswkiBzLJmN
hdOdxhcvMRORJGPe/HGGIlEl9ygXDka8RzghY8aCgubwCTeyouqEw1UtOcDA5XzrHrmx9unYsAAP
u7Ut3Dsk11NHR18kLUAEUtWQjQJ8atM/GT3HYk2UR1oMKZbDLjx1QM6N5ygEq6mfIPYEajExLX5h
2olFbU1xksG1lUREee4CsKhJ3RatSk/cP/QiKgGfWnkjfzw/nrachIeKhgH/wcDrNQ0/9R9sB1a5
mb7HMDtp1OxqRvHePXgk1gA1YPfeRqvF1GOJgQSvO0l9Jz2O/NCiaI4UC+CjpZslWfw5CO99XB9z
r0dZwABqPo1Pz2YJJeR8ClCf9LDZst9FQzocusWJrc7IewQzDOKTQyo4eBUwq/P/slSFDeArUmsZ
EFZsLIgx4vrPDwGyHrjiwuBgtcxDkaYP0BahuN1OLlEgaS8vk1PHxnPsfcUn5sapAAhk+3sJ3T9s
uiP7o5HhTURJKorIHIqLCqaETir3h7nPs68mq7NKbpVAyzaAYxLfQ6Kr4l/CQT6gPcOBWaPRtexa
5D3X4OngUVPwVH8IwOcK8jJiAiLEuqusKbqcKGQK2alXe0Ujao2GsZLoKZuRJaZt+yScBObcqgwF
jGyR+Qbt9s0dGm37ACqHpejKgluJBtHK9RnovWv+BiVxR3k98EhphfmE7SfSAo1NXMcOD6Ne+Icw
x6EChI6rKYAtCy42EYCVBfKUDArrNXAel4Wr9FJfzxSxdFJXxpP20EX8NMc+i6mbvQ5TOIXN+kXT
05HGxVY8oQJ3dzDuMX7eDEm7q+zkSvUWtRSvTUXB2lDhNeEJC2woB29nnwquqq+nd/bCTNQUzn7r
PG/mNxpQxh1pFVSAKv7+gwmew4Xct/Z0/VT1JZaPenPmDLApPd58KUPd1f3cebSk/QXoKjNBkd4F
XKhNdTklnCL1W5+sfXfEy87na2C5G8YKEDV0fGoRxEo/5dK856nT9o3voXDmxPSaPL8pEsNveuoR
UsR1OaAZQipNw4FKSEoAawUzPikHDgG8WfuQmSt2uQYNedu7QU9pxVhnf+wvTvpSb4T9/rgygOrM
gd+xYuxAo+0BhtHMq5q74qc2a4ZcAmR1uOb8PgfiutyYGU5lpiBKjzz60lOe24eYzU478xlvCHDu
PGZSSBvvtu1UgAyYoJHq7R/dP2ojGrgeQ/W3Vz0gehDBv6QSbHidTj3S7tludkxQkMvHl5fuTNQE
eRXw5NvPtfpbjTtO478wYLA9XybzVTtvsMNdhXF9kSGKBs+UjLEp/Qvyd8GcoVncV9UiP2clFQ1w
woyHQXuAuR97dgGB1xzSuFYkQPHoG6xx+XbfMJrt+g30G9MDkCuW/BtCrLXi4InZUlHNZnlTMuZ9
Ws1MQDopEi59vICg40HhhkiNnJZo6C4GdQCoYJShvoEGAug4XMCMCeX0hiTukcw2U1987FzBnJEl
e0/dyDUlHU6tY1024wntfVOl8DW8wlBZBG5zkPZbkkOC1p1rYmgiAl9Qx6cdh7rmDvdTOGxIJegC
nZ1IFvTPDBG4w7fJZwROdnQbnGqlk//TaMIGBT2wifUD2QbgA0KtLb6LrbTKAU1i7F946uyLAy6/
Obd4ZNkMk2YwEsTnldj5YcjCTYt+RWKw2DFVyevW824E6splSK5COstHxjwxNfHIehedmPUT2X6D
5grfYsHZyBK6HwKssPQZgeZw9jeLLxrTB8tHgOWVhfDh30y6F3i3bd3//4gnnioCjskcaVQeH+5o
K+9bG0PcJ3ndO8WPAgYC5zMTehpuigkMgP5Ko1CmMw/xGy8RNJM+QadVJGJlwidfJb4rGq4SecxA
jrOcxw39i3/TvxKL5E6RraP2xD2nvivsJvX9pwmgwMi8BBaUf/IsVjz85vJwyZUnuwEvyqQYgRns
lmMS1eq+Fc5WpkJPYVbRlOEwBCL4NYcIyW6ZtkTlRCaouIYjmjXVPTBSDCuAFKbtNBnF/Zw1oxr0
gymP6oMLfEwd6kRACZv3SBdnZufi7puP+mdSEJkz5E0n4N4gpJ+Yt+841jyLLMDVNRMgLXNNJVss
Mj0/Cq8CjZy/tfWY/FmtTGQN8leJXy2KyX+8Q0JEXLg4jnmgixQGzx4vMO0a4/Hh+jCWLct5LR3n
erKwUeqFaBcWr0gtdoRpVRyYWCg1uAknuh0ILUFCRXFC6aihyynmTpb6fxpTps7K7ArRQ/7N6LAx
LLD3Livre/BrEn0QNgm3ndxK7AvJP1h41ILnYauYJeayy94hSpLF+yC8JWFYYYhcYdWjvNZRI42n
Si3Cxm/DjJLzwNKO2JiehRTGPY2zfZiaCXv/tZDozBdV62VOdBVacimolkByw0r2lrJCi1EYJuOB
ZW2OWhHieLb9JJuSLnsQcYr6kzPYTYJxXPjcsvKD6PQTGQOZgweCjqdeDkpprzkwR70Fh5v3hpOZ
t36I6M+xFpN5lTTRqUC8c7xPoQdBS9ywVh2lc3IhsFVd3My/nR+60g9Of85DZnN1oxWUe/GM4jlu
Aacd79KBoAZ9VrmfDtbRer6CEqo40r9U1YXz0N2I0Q5bzdYH6kzd+6zN2mH+Yyzj8v8ho/5WxLib
Z4aOobWXd7aTrRSYpP5EmJHtPLfsaoCAhEZLEARe4Ar/k5hh+4eMOikgWXJXprP9T6H3pb8LguEH
w4rG/PBU8RRvHIHhyoVtF6jDYSAqD/UlKbOxQiDa1lcIcOaEyKIJW+VO1cAL6bhB+eNViBOkiy5q
BlC+dA1AdrdbEb0eNbLjMpONR9Fx9IUHfXhXqXPhf0/+FB8RTH/wMxNG8LFSGuD4vLhxiNSMkewe
QE/gHmxdvU2nT2yGpuMY72C12UcrXVQaHaXmXyk6vL0GoMG+6Y5GxF4ctgmzMraiW4q9easZCG90
WZSUSXQFgwniMQiaUosn3+VKYRJonqrqIRVzAs8btv9g68pOUCIMbWrKxjNlB/rvTpNca6AABn8i
D4EOqh53juGG/XaRonlSMEjYAFyWVy2+NbXlOJJzU+DA4TxR5rmj/VhX6vhvhNyKpCaGlj9dL4w2
/pgP9nCzInPcSH8YEjqHx9i6bNe9JiUCsrpxrg4MmVan3SzE9elMoOy5gwhoTcTU0EigShF1Odlf
1d00R/no7NCQspq0V8DCYeTYR0p7oxgOSHQNdoqYCxJpMF3usJPtYk60Xm25zUChQ1sfSUIoQ/Vk
qXjL8Fjof/kSbOV0gM9ZNQXZE6L5XVZrzDxgc9DDAQfKr0ppV6CZT3mBX+6J71cGc715dpbD52CQ
Pv0gio/vtix60nXimJ9kiBpeNISldk8JYA7FUjUjYqrFrWaXAu7XWiprDlzBNRcx7NRi8Y8lsaML
t89sf1DTmyShn3Zki3nVmAmSyZXV0bz4SUPCoSoY0t6CTo1eNL8ADT7B704sLAR2K2MdIM/Ae/L3
hoAhDjAMHPZYu05RIB46CbCe24ivesyOH+LKgoveBHWRwT6uFrdL1s2I9dlNOcC2AbOfa/vYCNF+
JxjtlWOOsoePIffT0KZ3FOq0l8Dlhnas24l53klhxm+/Rp6XrT5ZwXSpd+UX5b2mNwS+bofUg1lZ
U7oltWVJXQNm2HUtstAMN3TmfLV26UJrIE9x/ufWY4A/1T47vUfqJh37ZbBUTTbN30OTpgoRb6zV
shrB5209gg783OjUDTuFrILSEctl8K1+7gBXskYyAvKG7j8tyInv69b9bkyi7JrmsXsrrufanPp3
C+MhmVN7HZaO/bA/TL8Z4fb6u6XCGfSrgoLShe8gZhxRhHppWU/BfnCsHRMZTfPnIhTpsfBC79Oi
PBncsnCO24r6O7NlEFwdrwSv+m3se0HemtcTL+r7oGKjQYbBunHdYn7229tUZnJah1rEB+4qQlzF
rLusmVsA33erYqMUKA388Bis/FGpmOWoJPeIAK3/l9ITDJprPS7rXuO0HIHy9siNTX+Ytt1MC/Q0
DY/CAcUbiMzj/KSmRgIkCgpXWEnFjB7htxh15nVuhNWF4y1aioTGObRlxDxhr+G8T+Ad/uuqVLku
vb4VG4cIteNaiC0Rw58XQ0cCmoSBJQG/hcNPMHxZoLyGd/jI+sZSEkFlKbPiSGpvn/V54XBLWwem
PeE6FjFCKBuZS2fxuaK+UvAzlLTu/Ww5WN8igX4QnyyxujoLsLGBoV1re78P6wNS9qA14YZ/RjTk
ma+Tc58g4BNjP9226LrHIQ8JVOzrhqqYimDVuoOIHGnQyfaWsMyFo0BMwU8allkR5if6vWQSTOO+
ayv8HeqOT+xI3lLVwBJ+vJuF7uK4DU4BsaNHoQpxGhlj048xxZoofJeeXYGD/PhftDnQiRhUeb2e
9Hw/wJawijHuWDAlxQAxym638CVv4Wmj9Lb7O+p6eGQNuXa1fDF/7LHk95L/w555Ft/avUlPT6L7
7xFwxVNrjF0ffeZfR7V+lLxrUe9L6qodbYiG1vPDpkwHe94AFvI8va+04R2IY/wdQ8nFs2a+WuOr
VbbeYp0CdxIRqV+e8Ewq1NB9QijuKjRgywtvMBYqZJHHiuUgYoFb8QaOcJz+lq5x50NGzHt7xmFS
Q70jN70XG8WAYmOAhPGiasH2ZBKVxlQkI0Z4l392w1PLp+MVI5YsoaMOtmW9+uj7NR5qnI6OHuQC
p8fSqogh7Bb34udXIV10QcsKexEkaaRSn3nmxhZxhz/GXY9tbdHPOabWFnrWP7V++NXyHypE062c
MuZUDC0Lr29c/tKVY/bs0DPOvReLYWt9j6f6AnyIoGhE2w/g7JacQhl9SDvcqiQWBhcfXecukrKb
XjjNdogi2bIyhukiALoSbr4TEPS2i5jk2/AN0AYoFznxgM1c7CLhXmscudoQBGUz4DI/ptnuZh30
RD9o/YbkW4yfoNEuo1RTkJ95SHUwRCh32xAeNiBQDiLoabypJuXNfWF4Y8RmyQHGzT7C3KzU3BRx
jyL99uz2Q54UeJgFhQ8E4Y2KAUOPZLgjaaEquDay3W0MWNpDevreyaut7OExrF+4rQNiLzhVpEWh
GJKy9MA3+BHPpo9uF7oseH7ngO978MrG1r7d4pV+X9qHBRNfQPmAoPcxj5OX6mYBKXVWmxCvR2fg
sKRuNty5sMzb2dVJrLnAnKdEvxcLx1xKMCJYvyW4VgTeyHbTMGn7Moao6zFEoIWHcQYXXeYma/oj
5L9myK9T3nWt7kj3bmlHp915GjBgxYudzn2xRBnjwET5MCMU8apMLVps8FV4fA2yY0mjfQqCem3o
PIzNoZncZHLrCDuN96PnF/Rf3j1qOhclfe804iNN+n9mQet4jfspFrqIscdq8+OLnA7lo/Y0Kv6D
xtfqezICN3M5RzMn4ZSFCGsNG3XmCRMxs9nSp7jI3XT/WGUTf/qFffOqmxWaaX1CVywocbtNgNVZ
kMbIWvP5F+eBfpkIq03apZh254A7szrWZouxhY899GDBImETVJgCqWy2fVbRLNRS4HYybdNoJli0
ACKaF9ObdqxXFrC+ANW6Ul2erSNtIBoJMlaF+NpBaK0Ya0UecV0Gp/aXQNAStzDXNfZ8/rxPfrVz
PzA5ENnRWdqPbwDgPhuZNGNJe3Hn9F4UH14zVvlx6glwE0Hir6poCCSmCBvnDWVeWNwyRAxHVYvD
4zoOuUzUaZGDR+DOz1JKeIpcuQkMbnm59eo2mafpazyk6opSg4KYLMgz4G+jmxCfbnd1oSZkgXV7
YkMzPI6SWD6266busKy1JvolXKKS03Wpc61wmArVND5qYz8PyarOuPOc9KLVgX6ABqZ0QGxAmlwP
I62PCKYwHnuA9nCPzqgKuZ4D0FacO41NJDa6tjMcC4EQaWFzoAlcWInF820uATdje6inNq5SSy2L
XGHiWwXBYUwyc1BHa5FaMwOZwr5crMZLWK6s/SXJlP17idCtNFtyd/cRo/nfeFWMu7uNPJfSnJ8z
LeBr7ZFqz05d8XtrDUIuV+ThHxagwP9fzm8di6bmgUEXIDkh+Lod24f1tvt8K72+QvFM+1BzF6/L
8trkbcKcq9QxcllxoFXApVTD8Jgwhn2GeqRcIqVV7jqq7NrAZXaZJf95I3nNr7v3PiMW41Oj8lrj
GeiZjr2gjiu40xsrtp7GZoZuCWEdPSkRv75rqj8tXKP7NYW8DUKjGQdwu/0Z1tm5GUsy6/Bs4vim
xi+qZhIJ4rnbQDi6o+BQIqRHV81qLmxGDUp2dADgK8L622Z6C/WY45Gu/9FvaQBDG6b0X3hjr87R
F6O6/mTkB+EIwA1Ld4u0WwVRvnhr1lHSw9drFdsJoAXTs73ApQBURVJ6AMNYRyb01W/eHzLvLOKJ
6jyIIDdAIVxzYWCRfU0CbA/NoH1pFftshsE06SeyeEWk61h24DynjKXf/Bl6VnU54lgdpA5AovMG
b6WVH66+b8SfYAty3TE6gAGBkAbjuHpd8AFZ2XmiwvSd7BB3msdhSY6Y7uGz1Hfc8HkHDwP2Jg5x
ZgQ1OsqXYytCqFF/s/2tL8+ZjtVQEWHfRP2+M//oCKdW7oOYAAhlzxzBhiavYlNLRzrbhMb779I/
8r2jWu5oP5WDNVVaAxztXjG8oatURhLYH0SqO8OJOm8nhqGRKuUMbYWU5eyj1EvSlGM3qG9vDQ5x
7Hyvqb/F8faHAZocauJAgG3bvHXoskcLwLNpBpCHqjc+193X2vv2jkm8+y6nDn9ytqQs6oi4dNCa
+f5EiSNNg8ysYObilVcmbsIDugzzR9GWdtzKkpTy0MT3W2FV4qLT0AiwoHvunASG9MtcL4SbPh9n
9F2YqFV0VLKKrM4Js4Nixb7zXFtJM+zY3l5IW1gHTJkprIxgL51bUppfxg8kBebTPiEXO48JcqUe
3jgfr/xy+Rc6q9gGg0DGxvcFx/caB8/uGS+Q265777cm6j/LU8MS7MaUkl/BiI9iy/FwQOllQi9l
nzyRuFOIMx8AVXocPg5Mbt8D3/8luUqNy9hNnjvw/7aqdWw5E3dGZlcbR57yEwjY1/nBggNWQ837
z2JF8o5GcjhGk9kYV0GaoGlvtfFI/Sj25LGTQPiApcBKDD2FV1FC3C6PThQLZ6+7xE37OQ7DEWBZ
G34c1iQCGEhlnLHw7eaAn5860deOMNMp/8B8gQVAgz8Et+f18+xSEGWcOQQQiHCckZYsF3D61Rx6
A36IbBriaER0iZA1NvFF5IyzYkma7sCW08j8bA782nVQBe04MdAj/vQtkLw38p4NCXiGDLxhCtAQ
NRaeXaGOxakIQPAf01eF6jYjk6WxG5TduxGfB6WTXzDL1mQ9fSiyhgZIvVNBoCJknXSnsp3Lc3GB
SFdRGG7fpKu7cXil5mVe43K29Z9oMqw6iZTZ0EgvtTQ2m+rhhGOPyQXtHldqY0X6495Tq/rrNykO
gf6m0CJWXz7ZhS37uUsaO2iPOtjPee7ipmWbdSq8mx3zeWOVFWkmbXOr7L/uGxOpfOXCFJiy3Eu4
AkljiGIBReVKX/b5hS8wnSs43u6xll9L8GwIz7TnaVjCBbwO4ZtfmEOP70srM0VjmTDWip0wMQhm
4fXdX3Bbqbj8LV6/GTwdZZvH90nvw5kCzKfdaXngbaTzZELsmTbCB8mIUl+uKsCr+U72aTYYQEIM
zU5iHXmi82BWYk+cSiYk5rHpXhPrM2FxEqeT0xDQOReepiILuzMwO84QXs9s7pRy37ChglxsX+26
0vWS2ONzN9EwK3A/aRjWklQGMkraBbAEIgqlxV4TjI6H4DQoQguhrHVQakRCnAQBTm26/SJoZOhJ
NXAfUkiHpHcJgWoSK1CwP9EVU05MrRg3Y62VHp6b28kkPC/4tkdQAP73FQAUnsmvRICyvoqhCC1m
QOfnnTJmLVyYsVixOkro/mZBJYgUMV2SsNb7CTSexeN2SMc4OPrYem469uv1d7ZnnNNMhvh0wq1A
12Ey7K9nazBF6d5NzpSmP+cM4og/9BsAMxu4h5Z8aoW9UaKuFjeWGd/5j8hZvgVYP3a8TvsjJLYw
bcOiS5anli2c7p06HdRpRH4sJvTHs8/MPZNWdsmk72+eQKtCalpshgby2s6RRyAHiGMG42ugWx0H
v3PSccKsQRMlrw3/+44v9MuF+7xrXzlbWpPp/aR/q/PfiUpnFTJQHMJbAW+Oc2ueDQAtFI4R+cwa
Q6T9uV0RFfNrz2UuDx0TEHqfkAK5scnl3X/Q4BY9BKtQTMXnId2GZpXXjocVFvQid0NCMI4jhzhW
HO3RVaIj1xTgWw5cdJWjM/3InFtSQvDze2fSToAnA/triO+Lj0AA3FxRdgfK2UicEptOpFkvFqOd
0EQP2fyfdVvZKwlMxbXDNc2XVdwVK+as1CSn44T/7hrvQTaOdHYICe6cJyP0cAvMsTnXxkqQFoUp
3DLi5iU8H/Ih9xAixxBXU51r6/24IevSR6U+lKus95ORrcAz/w/vIwWz2QEG9rUxMA14sop0WkwI
iUBS/CDVbIXezntoO6xfqWzQeA/nJJvBFRloLdIWxHfdlbkfH8vShnpMDqYewE96aRJmdviGk93r
yPMTHP7Y7yQ5bKKDre1UPjYG4xP4lJ/JJAqnNkVw0XiR1oTO8HYPcfuWdRlMSzs+NOQCnNn+b3co
mjxDX3nLqbKmqCS8/X1dHHH8DrPSa+uJvCMKC4e+85fK5u1sU5So9xs053aGihKDLKJva+rI12+f
U58ADUwuH7J6q6R1YNEtAOGsv+Jt4qaNE28tTqilXURAjdPCmYWv3O2tdygirUdXW/bEaR9I2PGV
akZOhgnrVYvKJ7Q6wynCQNdO4FslDxKsu09RpBIR887DmvTGLwh3S2ENn6M2MkwqsiEbeZPU14q8
cOnwI8j9JCcx4Qc2q9g0dh/FGkapEwT4rap6KT1eHnI4HlCVfHTGPY7V0kH9/5zHU7Pl2Cd/rN9R
2L9Pdf1SsF0DhBaZlv+fn5ZGvrTseZgveDe5pgRNVMPZHXobA5tAyQX+dsqRjPJP/BRY5L1FziGg
OISLTBpA5+a7tVdvhBXUVS6PBttcm+D40LRBHaxAgWAW9eQDgQVCi4tdjdDxhJIthQz+JWB6YNX7
4c/NBzH//NpY0fz4A+ULYoVeEeHAMq2N4g8d1K5n0yI9F2JnRcuLwJbHstYCmV2a2MkSaMSPolBr
RYktew/GIELDmwOd37VWEk+Qd22VxPFNo8LwbpvdTTXkucbiYR8pqrVRsrMcrEHZwaJvSvyFEuyl
bk9JhTk2TsnR3WN04fVISdpxlct9d6y7DYdSt1U13fD5sdT2mPbI2G6iUy6ZfbARldi+UjqVwpgl
2Q+vwqtlrWykjjpQO3ooM0X3dKIDH81MAy7UXU6o7Nz4SjKFqQraCIeqoc8SdszfzfktxqhwliHM
pQYYuVPyH5u7/uuvrv4YRtw9F0FaI7/0i6zoHeqrssDPPU/j/EKEzRRf4Lde+Gl8IZzxDWaVaE31
EhCJ4hxYxjmtobg+fTVesnq3WoZvuijBwy1JDG9b5f1jGyqFqIboVpKJB+9m0YECF16+8uGnkfOW
3Ew38TPqw453mFBi2gaaxvpRvNeMJopN55bWuTmyq4JJ3DK+U9T9ZUYL/xFVUq9r+b/drQyOeToE
o59EvnYudwL37Ug4cQx0EIsp+fN/nhcQgtbxiyCSAqk+CLxLbQNX3AUv8IomulVCC4tYNy2nogF2
wzFf3Yc43nAEqAEelbWsBUJ3uQMpAMwbJETy1mLEZZ1rjtTr87kg2IyIW09jvmqyhEwk3fRrrpa3
jxAd3H9mj3NS2lwPqhoiYjjo4YtbrC933tWcEFN5P+hvLu3bwMWw156014A4NrSFcLgq6YUCajl2
v1N2IMkI2crO0bnk45O9CpoFoHzqrvus+gTUL8S+KFXEdesZm35Lre4SIaCXUgdA+qfwWIxL9/vn
LTL6e0KT7QUho5W7HM5EFe8ld0kaASV8Gs7K9b3JeBklWqplRuWEiSLbOZMUwzivYBGaY7Vl8fIH
yLSHR3uxvI5yk2ubWBWI14w9XUeeyurSMXt8tDTcbaZyomTcCUFS0Gf0+XmTw8OuK06fU5vwEzVp
pbHCSEQxGs5hMgpBtqwj0qOTOZOJaLGqG8QwwGgp4v0TPp9a6CTU0fiRAzcAH9/unO3xp0qMgHNp
a+h8a68OjlFLZI+4iq91o1xjOSqXzBAhcOhAC76gYFo5n/d2dFUHE57ey4dwjzZrEKzFzhn6I6Pj
eleQji+TulmQl8LlTXWsxiZ+JND5PsywB7bGSFyjsgEjiKMucwndLEERhlyQbTFi7QBev3XC91xQ
YFvxsMl5splVYtIO7g5/fzzTVkp08yp02oqwL/6L+yOtFDokNHekEbsfoY+OJlsWL8nm2YXmXHcJ
brdY0j/cXOdYGpdbt+OEG0eQxLy5G1gWdUvKmwlSQLiS0XXmtsQociKRtdTBAUQeter296AIZznw
W1wuBZHKkuJA68nQSz9T7UbjsxyFBlP9UsXDIsQfxC8ha/Z9nepeaVSA3ehLpyLtdJ7pode5pw9f
HulYDCOtcVGduT/n/TrHaLOTFvVwKl+HePCrzDVF/ER2PCVUTYpudSAiVsCscjAIh3RyO9FVgL6Q
8/rGVv/FAJkRT82O28TAH4zSUqqf0wAWNp92qMGsbRbUFsu9M/eU5aG71+IGTbCMdJ9uy+ThIJH3
MTulSkiunSfNvuMeqnWN56JSwSWD0nd4eiCyivaylArx65dH/Z3SxwCA/tfFnRR4G4/6ZaB8OpKB
6WjEbk9bri4Qs+syJ+wjt/GTgQc7L9DNMc6wb/Z9TDinkkxxJJj2EpCJQkl4wPd1t9E72qaesBw4
u3S2aFfgFNR6MiW6N++hzTD0CjM3wdFQ8mPWPLHp2IyvOn8CjyzigxjuIf0+mEy3WIvUfQUZUevx
0aJJ8Q0vtah3RSZQcIwIjGRd/iR35AitBA9RXUo1RhDPHCHocIjFwPrsEL1JTBpEXeAZWMkjV2hM
8IbhpHjfF8G4cZ7eBYwx1lvUWkZGLduOgDAtdnB6/gwiZZuO6VjXArHc+XrxocbKI7OP+BxgigvU
S1Dcty3VzDZwNkC/TzTDEBGwVpB2mZib/nN4SdNuNy+eTg/MPaXEP2d+XFmDyEivd+a5bFd03ffA
QNWs/Qd7MnOe2OLjMKs1UZu+53wlL7YtAXi2e1OucRzlW4RAZhRbjl5oBQ4pTlP6iYpZHOQttL4g
AKekIM5N7G0/M42v7bjpk8qVJMc8EkYHKa8Tc1lKohwMD0VmMi3x/y+f3SM1pMCAmznFqytUs0ID
0tZz7t4I2u1Zgk/6Zn/zigmixBfs4C9o7xuNAmRtJ5pobD6E3LTcjhd0leMaXzO3RYoXVKYQ89J0
F1YBYZ9HgYGMBOTEB8cQytExy+DdJivII6K+IAPKFX9jZLMWmCYBud/16yI9EyzBeBKCWeP8+vxK
GFQPpZWiJBf2Y1smptAUpaPdu3ANoMNxtNiPY8Mo0Vq1cy77R4jLhobxfuCsDli/phFv71KZBpc5
X9MIfKyBXik2HyR8vsBBvFfY0ek13bRe9ULg6oHlXMQa6CFQyUn8zvLvhu8HHcYbc4LesPsz6khu
MHstNsVQxQ4z7LtzwesupMlA58kMdZlcc2MQlFEK10QUGNgAT7aOAOME1y7HkFstkpMFcj6YICna
qJLx0cPhJzEf3K+YfYOIczV8G/bxSmE6TeESIlVgwWvlH4r8ptTyL7CuhKif9yklManikHFsFhyh
zAYTvpZHO8Fo84rRBmN+t3c+1BCG9dNVlFZqHH1CeB1gBKEqsaU7Hz9T5jgKXF7LavfQNzJgVlTC
roDU/EzrZVcwm5wubk+U27cDRRVS1PK60Zw2n4B/AEqXuVeaBQ3cr/3pomJ1vaxAYi0O+zMu5wby
6IKthQGmq99vryKmctO7O1YgvQJfcq5IlLaEITblfcxxunKCikCEVVM5g7JzA3K1FR9c7TmhUnCw
IL/PruB+iGUzoBvGbnQiM6sjs4kpYmzQU9PlldJzSsVs12zAixsl8nMNxHOR+PD20jivO80aibJx
Cs7K0mIAyWFoBdaLgGezPArzLU2UlfvlFel9GolwG01k5/q8Iqpf11/vBueBs8+i5+p/Dmu6k3OG
EbJDYXurOZcM3zxatIXHc/o3w/72EnwjBV6E7XV7TlUd7LjGTK5X1xXOr5GjQXt266goUAGrLinn
ax4dFqNGXInrQd1rspvL4DI2KVeX2Ts52goTwqOBhBX49gci9eBSULtw7TZ+ccyqtQbe1rQq+l9Z
u3xHfuP9Ga61EdAOAr6NwRe0VMRUYg4eDvQ7Pk86b43FKyaQVrwyeqETmtcT+AfKoUIF2vT34iE9
x/xrSjGYMZYrllgK3znTMqiSrNTcF9tRFfUl1k+9NGfNgR34NCCwScgfls7TGbVoXLKpejMtcwft
QSb/45HO1Qxp9MR9oBJ0iOpZx5mZmZVXROZid5jluPZgxWCSaZb1zUOBbZqaRm/vn7Ed0SWtkyZW
kltJqpIFj49TC5VzvYcI7nEW4vg9f1Lz7afIKwbIQhnLA7HIITyKFSPjekx0uWRiiPYiKPIw4uj2
F8Vx0nrtvdPK583jf3V+fxnJ5lITHKqoUJj9GFfHrO7+WDB0hpcpy5akcnxX3c+Qgl4MNxAjOoIf
MRASpFwikOkqFBgwWOlOLWqDsZ8c3X3iJuLI52m4SyFjfFwI5Ki1JcB7Wx/5XP163++vsgoK0cPI
cPdIzEMvgOjcJnDb7p9vbFR0LL0ry/PXVTWnu6BS07iEcNKDlwufF5HbL8csg9/qbVHCyuqvu19X
CkvOzaDYyIcdjR3Krr4v0jwOub1F+d8WfvvxeZjqCJTOSMn8crysSMEBHBSFfzJoB9f/rm8by72e
mwBpcMlKP1v6dRZvj/Ra8/s1laHMRK7jro7WZgpH6TEvB8pXRl2N00e+JZD2osdWz0vRahcZ7kf6
U4Vwmq8avD4SAOAy60L0eAi8h1FWfincpDqyhzJ4ghaXRsuq9V92g1CIxvnkRG5lZ638mo0VxPS0
VmdoPzabXtL2/iSe6s2uJvOswkin42bHjDI4qq+YNI4KzMzoBEhjIWH5K8Kr3W/indKCHY0jieej
Jmy7tUQbeJmoZSwWA2pVR/A3HKfGsg0sGqERENcw7jOzzBxYEn7RMnBhEkVJ/f2ry3ONaTMhN3cS
5wt50r0bDotX3O4yNWaQEioDi5KCU7oLmmBk/MjZwZBoBHVZu7P6bCKDNHZ0oiDoK7GKn9m2/aCl
3hEkES1LLy9NtyZShBMXqu/ZF5wbJYUvIe1/lhA88tpjjXU88vzCOywUv7aYzu27C86FSpIWEe+u
Tx/8BC78olIItwc413R2i3NR7PgOsf75EufAty9yehz+hxA8c3ea6RzkoedW5vj2ZysAVNJ4ipCB
Go+KJwWyULYYLJtCXaucocqTMfUc1Smp5C7VxY4PJ+pIVxPdNX95jWgmUXEruQtOwK6SmdTQhsPM
xUbuPFUJE0d7F5oHgsuQY6J1j0hNCXL8pr+4ivJk+3nqQeRQ+rtd0s4yqWRTCf5tN39NZneJHXXm
fnIh6EVzVghvz76yynjqWbGgKq5ZeMfRDzPwJ3R4y9wuq1d9WvW8+QLHEQSNQRyRpbSTvyw0SEgh
bFohroUYIq5G7vAOUJ2DQ0g8Sxv4qpPUL27KXT2bJ1LJD2SIGCGrKY/0b6znZdVmWyQBE/WNqCty
B2zFysGwge+lr+Qo7B5DUH4tqayucxj+pntoNeYxrNYOvsJlnw6o50duGY9luP2A6pW5EqQvyhn0
/nHXuI0jfIlqcRsDyqDpe1XIsTHtFlUdCMunjO3tyElpLsimlFqZmf2yumLj3o+2S6vbDcQvbUre
tIdVCUcqpcRBHYi2JuvnMGUs06Oa2/ujmvP/E7+5LRIaQ40+uxMKYWFRqcaw4Fm3+REhdLQYKFlR
7BnwoJS7v9KyWFBWx12esmt5u1K8cvMD0LqAMXAfTaF1+MJc963n/4xWWm+/wqngUM/aKiaCsB6U
pqY+07UFrt8wHi0d6ZhxBboGPFxmRqC/bAq2qey9NqkDKFMdmN/U+rqfYsHK5GGvtOlY5kAIDmR5
qXWDh8QqJHFwXk4zEvoKDvlaiYKD4xHzR+25kAAHQhnark+LskCmcU1v8+4LvqeT5lcVphWshQBW
25WOFukdf66dPVqT+5TEhrr+nYEzbbS4If5oDDe6IQzco8Z/tyrX3kdQZ2Ev1Lip1vUVftRn3PNG
MKImi4GSKt9FisYHPhLcapsTo4BnNM4i5nOcrhhdx6012+dbaN22nyODOOFwMSvgLzw2AZwoBikk
7Q1cNkfk1KZYG+GH4a9gdZw41qEvBnb8I+bsPFhIXyiUWGc1l0tI9eSPps+xKI7luFUZjbcUxQTq
jPENncHPLjuzVr75N9OJ+Ubfefu2GryIiYomwfCuQm+H1szlX9d6A2zVM+qslvxzYJ0otYXC9LaG
C7n3FdH/GKLZ24zMjRJVI2ARlg/oWjZsrcZBNtmC5p8cnQXRIgUI8vCjph9gmTjI9h7nOQpRRQ59
gkys3k47UHEt6Wv+ivIv6qOlE0KkLOTLxctwuf8QKa2U+sCg9Bcd7hSH1aYp1NVA6MBnyuBJ/aHQ
XoEi40T5bFw5iz9yyVFf+Cj9e5VQ7kzxMeWUw6aoa9cxHMpwUx2ltm6ZZ5fIxLGQ8jwh+VnFhfgx
StLM1fbJXKIsK/iZi3G8HSOPkavt/MhPFM1LHCU1NQjlEvgGFVt5tVNOufLu3YI8zlc4k94NLsGj
F+oCjbDufL3L4nVS+zEDALp/0IiAg54WIbflqUZB3We8lzHCUZ5NxLbIK0zM+bgSs37Ng20f5vBo
S423ItzRf93rkZfLlCThCP6aqzF2ecvmLcmAAbDJoHJRJ1gmmpM3IaclT9qt3mdeSoICBcU6rsIl
up15nNq7eRrUm2l4LjZNLBPhKTsl54kb89PEspnceRmYURhaF9Tg3N+siQAdkOT0Phc1eB1/NyOQ
IAkC4OU6av04wbSRgsIpWxgt31wUNzzjXQ5sv5qtIhF6tAG1IDV3dm0UaZX0XNwZHzUspfSJ+pJH
RlSL9AtVADNzVKKZ29T+SUDpf7pZ5qV6QmucNqZl5arYR8UTI03GVBBMUAwwRCufO4BrKxBd5Ky+
INCbU3ge1V6ZqbjWOJ89y0C3MBW6Anhop/s+5D59kU4w90+tklVr5FUIaPgrPZElj5Pkf/09mszc
bTB2Bl6ec0Ofp1+0V11OvLe79KvaZyJgl85tFtlvJgBwNWq9MkfJHuH046osMSYVxGXmI15HFHSd
Vmm6FH97vOY9sn4ILViOJp9WudwfhmaQMB4Uh0ApMCtoz/hzzZ+BkBL7Q2CR5Oai6NE+DfMq65s2
urZlISe+Wh5G9B5iyA99nPneVjSRXEPzSKuZxMqaV2qNPUULK926vESwuddR4+dSWzpUZniVJHaV
k+/YMXi97nlHMZPuNPiSUze3IrHqL1zyHd48xXIHTo4+xhb8H7Zt96MhYJ0j/Yfjcrm7eN2hu/Fw
nvSjobtd1xhaN1kimSOkA2PSYdi5Qzj0bTW7UPLPw+dQluewQ1OaikIClFGNmvxTT0vVu1Akpf84
oeNcgbDXoI2RAvMzwKZ5nzG0L+44+M+WG6fWhLOns16sLUz+LxSTrAJMymUd2DEL44YSMeRo5gkE
l3FOFCnW8cGtn++3eg/Zto15d7O+QaUhEq9aqKHlh7fROOmLd7a9xubr2SVZ3VXMpx25l/8/9hoA
wRJnq8+Q36rUg4r8Og3KxXlWki1W7fkCU8xbMsPeVhs+wX2uTxR38NbN3jRokSISnEdQLwwwFE7l
VUtrC52dyHEoA22UAqH+qZQdl8vgNas4JO265IS4Q/lIC5NlU69ChbvptLIql7Iq2odOv3EejBUY
uB4QtAOPXK+lj84HOboext+7it6O0iY4hPX40ZY7lrw21CbvaWQ0CEwtCSWz070f9NN0LA/CK3HM
TOT3F3DEediuVwe8bN+5WWl0JCskFkIA6N/vP3qygz8PNF4dY9CJv2AkPc+Xm2LyTXpTGAxAUkHh
89rmaKnrJoPAS+XH1onv9W1O6wxkiEbmpOc9xtUrVtddMcqjwpAs+o5yOlf2l7WUufpb2L22fNvK
IZgwyQ0Ki7ooZomAuqxDkds1/zkB+6OgAirOaU+GUVwi7O2Hor3ILOeFx04dyWx/b5R9ferWA8jK
CJa/ccXOxbDXnO19Re2S0I+T3YUx6fBH4LhpPyAnqIcc471m4w9urE9SsSdSMHhvFCgB1GH/qZi4
CtbVkKQUVr3oIc0tDD68u77ti7r1aSjqDwohXcmHBPmalf8nM7TvFMN5sdatgm8R7l9eBzzINwfj
gXpejbHtQWILb5PcapzM2NBbGt6anBAiUzVnQqjrOzdcdFgexHI21cR1tCM5shIs3XTCeCNfWYVN
GC2NagYklOVnL+nLLyhhSWd+GJ4Sp2w9KStjCYQEyVxF+4AYrSE7e2xaSUqLlkwsI0NBCMsqLsam
4Hpvajznpf36CjMvKtEN0rsRa/ZAo9W0pwnVKP3QJ1ttdhPzZPW1x4d2I20JlEIYDIafs247gPTw
OPAImFtBmnRVD8e47TktVoogGe6q+DRc4kQmwnPSgQhKaovff9u6Z6H2MysdYMHND+9eLYCS1Mal
UtAW8qQVt4GTi3nKxJuomP7/7J3XfWZtP8WTVyBLaaJfeuhyt8RJt8F4k/XujgsV2RZYa99y+wyy
tZzU2FMXbWzV8lNstcEMgeCrzLsenV9/YqkQPqNXzqQ74uPQwQ2yRhgNn0+Ul4ALfOpxY6ernlGV
ulZ7JG1gG54mesA53GAWn3nf4cI/K57zpm0zcXO4/xz4SpZMRH/x4JXECha9WPriIpQ5FMvyxA7v
nkE7l8yFoBHpZFgfuxjuuLA7cbAlsHuacV/RpU6hleMSM6mRnZ0DHiPItX8Acn3fi1MMFROoAu4O
q5ARHfHAXthX0uMc1SRG1hdByZeOF7SS0edsik4a8CdflclkxJvo0VNh0STZ7VTwu+vOsmzvDuWP
ig6aKhstA50J+EphoNeNXO6GKbmwIgF5Nt6y8CSV5RjNUztuhkLPw2s4t0Grk2Y1g6Zhr4aILwHQ
wBgyFRWCqB9nOblSbt/o5oXg4i3VizeK/ova+z064YLIlHSQNzD76tR9WblQPQmbhj7ECPbbSNTR
+kvZQmJIGGqaAgwD7wB7zSVP5FM3hLUaT3P3HSCQJHFC+6CZ/8qNHStG0L4bTc5Wnv3ezMgIAsz0
HOvVjJj12wyUIrBub5k2eyWY9HWy5IcFYdliuvSg7UHSCFzYHGf0p9eFzaNug/xlhepHN3NRCtXV
+tFq0QsoNsr0RYy6l8AozDYzXIdZB4AqC2UwOuwBN97cuDGJkFm0WttqJGAnW1F3P5w86s+YslO9
tEJx++gRBRR/7ujqzyAojr08heFP7n6VYebBEn5F4QpTfrZBCTGGXKfmL9q0KHbWAwplUqq0og5+
mHr7FrA1mE2H/VklrE3+9apYQ/BMAflfDlwWV+0OtDqjN7w5FqRGzSkcuiZWaptQXEsKXRk/jd3n
oWqfsbNrw3cHh8gxg1CJIiZYNZFiLHncAwrZsvhgZdXLP2vF/dreT6lDvigTdrjNUBJ9pRo9Vb88
iW1g1cojK1i6jZd/lwn1pd4x0SuGBm9NJ69b2RMR2ZouN6OQTX0wHVo3b05ysCO4+icFpG1fEi2n
r4WacX5d9zDj+ppuiGV1BsKyKYK76Rx4wSohZtSbD4mOSYf9zriKI2EMQErAckPTS7xjmloWAiQN
pwu1Uu0bByOD1vpdpnsp9URl3EgS38SkDi036C0QI+fsB2iO6GnL+LcQ/GJHWJl4mUZyFochvzbL
H5olbpAbJcxn5wrSJabkYpzSPyep4HLcG1UTZAKB3t+9rPeXUfT93CmMtrp53sjUZOiQLXzv0kLF
JvPoY3DJ0WHAjqDI1n/eGRwtg+mk/GWiUK3pEbzBRr2M3Fk4Hm70BQ0zxb0F/2ncrGFNcafPu+Ul
8lbLpeLmYar6bPhiW41yEwuO6cVaewEU84Mw5/tNzPVbVmGLoO0VRC6XgdGQzEAJCZET2Gvs6thU
gmli2efd2Kh+g2p6sZjUckXGht7E2viTPXL217hNvPgbO484vdUn6791yYgpy4UjoVyI/LL/uSne
dsy05akDyeO5I6/UCkH5kI5yU7ey7QZ8hNnz/xPyqFUf8onO52k7waSSLdfVwelGs7a/JY7Dd4CS
UAqnA9HTHp7tnjOpQUGJXNIazmzKCPgpnVMKfuf4srmQMcCUeA9b3RgbG1OZEksLtDUb2S/4hxCB
WsXIuX6UaJ8zYb/7Fr1oj9JYRvph3jkIMY5iuT9LfLsNU860cnVTCdBXrboVgWPi9zV2n/aEFcHe
2zd1nvmrYn08dR4P9bdTUlQBOLRqLS3G5EJtXN/Kf7roSF3gzdb9OubxBxPqwcEKFbkneHinRjSD
Mp09Gaxkc34mavB4LC5AKmvxtcBH75N8QxpdDDsLJSm/Y+2hc3k4bYwtpT2RCR6k7nzz5Nk528dJ
wCsvqIKeaQiYBP5YAYCCDNKnGYfiq8jRmrD4khXL2sbimiFbKIdbrSF/S5QVBCqbzLF/TB42Wi98
QzXlvS1p0YoZSDXV/UlZXnSBk7PKqAf6Ym5yjb9N7zUVFi2S+c2xhR+jliP8xjcal4/XYl1XziCp
VdF1zPqW6ftuAB0HMBCdGHUU7N96zTYd8GmOVCdh/je2kRwGjQnlRCJHUC/gIQFvxGqe1JjnAQRb
fsTDWr1FPpBFrqhAXjJJc0LwQVwh9JdCwznfrJM8ew10b6PSoBFGenSXnWaYYIVZmR891y418kG4
ohhNV0Crt67gEvP6s6Ed+K4quzvQA5RLQFVjJR3TkUzLNA4anwLbRklbk5BfLqlU1lyTkjClSHcT
ycaWSIh9bxVi+Pt5a2tI9ApnAvIriJVmRQqh3ZCqqXQUVNZ/N+/4qmSSN9JyB+EuRoq66iRf+P3O
A6c+tsQPKIyAYl3CvDDarw+cCOGPnY2W6Tp2tpDUnDctQujPSSuwkv1cNrt70euWnogEqW09MI0M
OoglSM9Dkhdxuj9vxHI4B8v1Ueyig4RaWmEC1ZLvi9GFdO6Ibglns7j3+kin2MA5415hpY08rWWh
TtaNLy5jUj7INc0+19xAVGL67240YHoL5cjqguHVib6TOZTmorQmMZxnN+TDcC+ynmaHTvATned7
RAV29EQLeoWzQtBySsMzxXfUCoCL/92L5BZIf+/44hsIFAtopzn4Y8fr1b2g1q3enxV1PeTvHAWt
ra2rYnMlc7E9VcgpGPQ2oyUmbzEgPrGMfBfZmdYIbNC6tPaDLFQImT85Lx/VDV9Im317BVAVuS6r
mExc3rxnKAgR2dR2d6K+j+mYLuHVrF4ZeCK7TS7OQkNDv19Y4r7sn71yL5d913USU9TuXSKUUFys
1OdP9XIkzdCun8j2Sh2GarwfRr47LBjyTXEilkD2Srbutd7Zri4DpwQRJ3Xqhs/O6MP56WlwBM51
6FkxjcWkQKXU+phUpcoeoNZXnzBVr0U8gSjTgIOkKl/5SET7PxUmH4sUn3n85jSBYsqJeWS55GD5
PjdTKbIZ6h++mQ2Do5QznJEHe78rfwT63nnCW8ckJciLhC+AjWOTbH1KCElCICki8mRUEsvYPa0i
JcD6TNZRtAU1F1GLCEQ3EYD/BMeEpEjWuWpkOdhD4FpGxLxN7TwjE5fG6KRZxdaiBfJlG6WumTpY
GkHay6BmJ+yTp7KmyTRALDtt1T9oT5W78BghY0+A/Kxovt9LFm5i1OgPOjrzuqhCyfIYxPYtLMEI
Lu7mXkTSJTBrtB+wX72hId1Bqj55uWY55aHyDZyZ73s7wk72HPO9t1QK9aDlMebq3tp3dMR1Jzxm
RVCNLh5EtlK2tR75cKX6iWZk2zzZlCv35AMddUmu8jLRd/MvpwfWhxHdrGjOuF6zsdrC8nlzj4ba
hDYFRjhksSfB6zvS5me3B5UOKWHXyzO4nqmQ3sDTevokbyxvmoGZRKEnSfw2Q0GT5lJZWy9+qQKM
aEiklg3+wPhnlNk7ntel2zYwdzhfDdzNZnUw4F+qgPxp7qaPpwIa+RVTRrBwxqFpb1d6Aydb5xd0
7hfFyonRBytL9ft1eMBIOLdqKzUeMZh810v068lFwfSr0awtdQN6WYWbFqZbRZw9HpgdwJE5zaQq
4NOURSRreEb2nia0U3Lrc7CG/eU7ZUGOQVlYdkgAGfN+b2ry/AZgAZDnlxKdS/DPUMcqDdcEV0nz
xyfh1riNJW7Mr6idg9Z/7cHBVzyemJsvlnHLytDc9lIQeEpLXrF8N39wPESA0JoemrUktEuFQ3mG
I++mIR4XOV+mDXKVU6pHypKblUjdVTkTl6fOnVjdng2duov3Mcy6NidUuIxjdum10RQDrmkJVeol
BebtJYFLU7FXTXOr5ms018NcPByWOQ5Q327N5t38MKU2lyGd51P5SmQ5OxGjk1d59QA+KFkhzVzr
Ltb36k7hFLxZdMCs4htbqKQbW2PAJYg4ZkCKlCgv02bQeJitXdCg1EdqegUs0jLm0jLuzxN72uOg
3GfR5wFA7cPlJpIJw8MnTAB2rYfJFnJhPE+9zJx+yOMkArY6ki4LiykOPd/ZFDt4gUrwF5KUsytr
rCyguiWOaboF1nsGNLI7tFYMC7qgRe61xBm+spmqNCk5UPYQ9e6KZE6vGBAKu3jDWbGimQ5gf08k
Pmm8ogPdLaG8k7Fgg73Ax2kZmOGR01FrrjdAhPUoMB8fxNhFeV7/UgPdh9+IUa3/A90ZdpALbkIB
CS8LRhpUlrHsc0kmApmjWQkTTgaeQ6s2QfLyI0ixIAWwwaPNZdeTw68ncXpGtf9OEY2EdS1iFfXn
hjR6yV/2lp6DquFaR+opmN+/NcXm3NFncOjGb4kYksTBHjHFuXO6O5d56LrZ/B1lYm55RFq8lsh+
q4QugAFu0QfnBPugE0xVBek2BqsTxQ02n/U0xu7FuMcOG6flak3e3hIq9ehX4jPEWZ4Iib8XKMr3
GNUHXLHTSiXMO+lXBTNHIs9/sahJgpUjV7HNmTuzboYxd2t1vv+W6cJED2QdMmIjLFbakRNFmRmF
0ATGUP3fKmHaZ15VC5+nSoH4wU8ZBjFKdHDES3yIa1lezRTkfv40IDAkhI63om/TICwLgoAm8xgN
vG7jp7HfOQOOQiqIzJtB2CoanSl/QIrcAjnNRz2buiWd5jfAeHPpMSQyHCaj4Zy02seblKzuqnwz
Z1mO56DKD9KLwdnmFcWRqi/BofVGaHASdR4dW+XSHdMoE4bqfeGKxx0fAzb63YmGTUg60jCOGc18
e3PaIMSX7BiT9IZrVArFTwZJGzTOqqhGY3ooOtpoPo8kTISGAfIvIoKTMfpuIKDKaWncupccs8Mp
4F9CWKyGJ9dMc7CtlhATn627CIyo/Sh5PnrbrR/Vr46u349e5+CyWg8SaX1qRhjT5SrZYEBssOw2
nMTGlh5cD7C0Rq25+1E910kH3JFhsbZ4IPp8urxuu1Dswqo98uqvdlRtlZ0SS9mf9wY6USDu8Ied
G5+jNWHnYLsbWPko/rnB77HHNKxfPwuBmym7UeDfdSrPM2A8NjWbG/PMicX6pUgumshBc6Xn2Uh3
A/dM0c/Gkd1+scbbck5EhXnKCh7Zr094OCbvJfW4myLBDDf8PWjlfZvjaDIcTBvqi0EtGbepwPDy
K9rx/WB5ZuAq+UE89alYMOedalGoB0SBn+AimoH4Ij1KH6URSesmzxHeX7g/MXQeU23a4QtpTbqn
p5YzmMX1/ayU8f/WKmrqTM4wxngoHeSNexIbKI6FPtfo6BGZcJOPFYC3H5AhlFaYdS3VMZrWDmKv
qwjVj1Xm0U7afwsw6dGLQtFFoPZkwurbDB1OndXA4t4pgmD+Gc0EV5INnqlLpEW3pq8ZgqgHiGy/
BIte0WHFRQWkNZMGRHx3zJWzlcydKyTiTs6AGGPbQtQSa1LaQm/8ooOlqTKwbCaS7T9ct3Th7KL0
l2sns+ebz+jpd4Qa9pkgpcdVtsb/NdTG7alyv9I4rVU9o75HEkHUQ3fLTuUg7je7KXNiOJ52O9I4
ncMJ6+uiFU9Gmk7HexpvyYbjA1scrVkcDbb8untIoCe7bJqu9SBv1xXtxZSJ7o+LPMtFFRAsSPPv
l0XYnvq1NwrSxvzrqMK2oINxxoZrwC1ilMvjW9S33cjwrebxVHjkdTWidw+JaBuO3Sf2f//PmCRX
FnSuSsC3xfsjgRn03IkPMBiCGlOTUMTNQMwCorUc4wpqLDSMfFekG/J6vY02x8Qrkld3o6BEYWfg
mK2DPN0SW397E7lw65RZ82PKEv3suTTysWHAsKO283nb7w1F10YJKx8qg97GkjNd8ZVFuriR6GPF
GITJcMo60YgqsK6UHNErmyTP0xi2JQK+Twce/UfcsG7Xd47a6iDBtQ7Y92abecTN9osRrB8VNpz3
e88RdzADYGqoLyf9i0quLm46yC/QhCkFO3wGx5xACtRwLBEw/Tpi4b207ZYgsztNp4xlZk+ikRV+
s2sRHZcs5B4MtYGCYsfnUMRzxG5SC2zevzdAyozatLEChMPQb662dwjhxDuelJ732vWaGH3e8Uor
LwuMqlce3VMhW6XD8CZen2m7Fi6DKFkJ44k2vhE+HtM6FdigPLgZUdykLIVYeTM3RdeD3dki85nk
Y89byr2iXeKvGC4RR5ClerbAfc0cDKQStX5t/sjKZevigE/4zopUZ3XCLJX4w3h22fEEA6cmKEsL
dwphu6HS820s21EALeyqVVOLaPRiZ7CB5DYQVPW74+mAPn5PAtwsEkt3P0Hf1QtkGnX9MvCuG88i
VIPuJXzCZjjQqVqp24XpFZIwyeMFt12u5XQvHtD68olFT1YydTa9D7fGeIvoGei46BZcoQvp9BjS
uU0H9F4FdHa08JJ5qtoRjYFq4LZfsluJkFvRWm49RjaClbgC5L5EA0hsSf2DZ8FJAaIgryEEtbN+
utaP6iOCMt0bqBNGXRi20qdxggGQormGKOQqoN8dfEub2wOyCOQ1s4XrJQ8YBMto4Io8JmkFW8XI
nj0ZWB+MrINq2bUYplzHofwrArwqTrNVE+pUYeuQnfpwRGSwnehz/u9egSSmzRqYzkU9b68EMTTj
hTrHBDUmIFoY9+VFj3+IREtYBIU86JQ+EXZjQdnD9Seq/2Xzg7+ygU9O313p2rtqRMIxJHF7BeBW
hIHGi5AInIPwctBLJ9XPlLJX2pJMn4JTmslBl01dSBAc8vW7/M4bDH96E4I0wIlSR1Fu1dwmS6AT
1LSBo3GR+nyqpPdKMtcxwEtnKN+pVNesq1R9Z2OCWm4IjuNa29y66IjoDjqj79z98FStwefUu/Q8
mvIr2w1CaoWrY6uc+15zawMLUdhdmqL0juyGzeTP0L1T57Lmrz28wXeGNvdX0GV64mth1aPXQ1Jb
HKeNCrtLPEljj7fqYWnDsKygcFSInnxhC2+Fh6VrhGizgIxbYS+COr8DxQ43RIPQQFHT+gIFx3sB
3tw4omvL9v5uyU46BfEEQ5Q9J5oZS6dKunMykefRfNZIR2Wi2RRHsIfKwiw8LvIhEQf6hxOcla65
oe7ikafy8tO3kheGTxaJPiL3rSwV7En62TXHvlqDlGv9xFysF6T/t/Tuuyu1203VTtGzgt7hGg8+
XRTGF0prCjT6DEHWyKFXIDIwBNwKGkh8GOl0FT+E0ATc4E1QvyC7oC2JAq6tscgECAc5tNVMWkt3
sXPo1uyFT4inESz119G3RR27H0QfrIK+KTr3AFuwLUJjtY8Bd6A0tzHOL84SZBuTCREJDl+C35vC
848LKdBQMCH6G3vdjhlKn7bKX/rYMwd/rlRYAMv4A/plzOTBPq4N5KxWTRt5s4CZsSEvART6NGvD
1iInnt3PuJimLp3cPfSKUwys3YaZ/lnO669UegBW/Wkz50JqhiDRB4BkYGbCry8kybH51IXYJABX
U71I33gx/ixqoA2Sc8+xl6dauvJZT3tD7SK0gfTCwuSqVKHrWtjPlD0yAGS/uGLnIO1sPP/3l/lA
wr66txevsVDdgS63vYyLehNckvB3s+C9iFIZ+J+FWD9x9xyvGRyoLYwJrGyj06QaTR7X09nW+pMz
KgAh/dVsXiExPDmo3LNBdghxds+kmBs0Y7GcCLd9tjiGWBb1YKcnWNKSH+IcPIVT0xrJPi7IIGC1
5hi741904Y/KfP9rxSSU7CSIOpHIudEBlboA49unuh4hLpjc5E66vcViyCSZJIH9f4MqLhgluPKi
p4vp0KvO4U26es9tWBXs2tfUhXLu56zRQPk94UZd43fG9wVyiFagaDR0cNubQBxFjGxBuZIDAmdY
VW437D6UEUxjKt8pZe7Ym7UcOjpb+H8cgTtZWclIBJhfsFwca6/VEuqoaT0uoBbi2P5734dM6xl2
Aa81sz2rkFgm1rV/H/ZdsKATLOiHVk9hJxyUM0cKdsNUmhFLV9WffuKjIMdIGFNB5lx/MezaSCYq
d1I2Dnk2qUQ+MaFzCE59IhJ86GMOUZ6nmeIBOpJW1AJ9bw+03UA6TVVZ/g0SCygI/CmDSHmQQZ6y
dPW03OF6KjvihS50GKClkFeF83L2QTvUmpLMntDBK4oCgZN3JSGliUIKc73GBuih/w2ZQe/8WZKR
qhpkUyaCkgAu5uNwS8wIYtvuyXgoKgM5b4mTfc9/0xReA9VvsbXI0hunHogbLeZLUup2aggk/5hD
bq5y8jPI/zpPeiYErUHDlWjryOSJsMXWspSeMgWrUvCSPGHaXoh6RbH/443cBFPd8ztvgrfwtDfr
ElbbaDlKBr1705lGzKnocKcd0ZMh4/FEPKpSQlmmyUmFm0OIs+JKaJzHQ3wl7k+gcLzIx4hbvRXk
TNjhgO9SlXs62kARfR8xdgsT+RjnITvi3Z2nYFtf1vEN52VR0cHhdZEO0E/dUOnI6rI9sIxANVVu
NlZ3w8m5JFQ1zOfdiA2BR3tLY82YtGoK4jBeKHRWENblXcb9uqg2/boys5ngeKEdSOGnGc7wlMcG
4jlhnzKVCEZ+pOeePeX/9Bsv/031SfRhGzQbSVFsY3+7gt1m2u2C+KAQg60k3/9LnGg4NJ15goSn
tBZ4U9bObjrij4bh5VnghCB05kB3MJ2zaFZsInN0PkKzziD5H2uF7oKqk91oISCMAUHTFkxirzPz
wFJbOKE9jhVsL71oSW/1IXjVjARp8ctEKjFJyPXnV78htDg0f5mq8gbrZo/6CX0FNf2rdZbSSH9l
us8FeN1nIqFZQR+4uZ5L09HMaqJ1loZIC4tT+/Gj99vOJkQBSrJ0Cc87tKR9+Vw5b0+FRuxeFT5i
MaIHZdjkjUTEHNw60mBw7DF0hYGBZMPM6lc8fEdVDRQNXR0kuFO9EBeCCdnSVJZjPQJQLfvmLyXk
0VOXO9dMxJtQPjjCydHnSBGSuzyeeUAdlbLWporw6nBMS8kKzMPekfxGjESmJvF0mY84wvyaN3Qb
llWa/tlFmXK4HzwNsULjznSL9z7NujnUgbzgLyOFt99FzPwm5IMDh+fyaWdbcHp3InHT1Z2YDHVe
zLR9ZbcyXm2AB5U/KTFIxUDfWzPcacc4y7kr0hpigM5ljXsZA1XPAaSPg7i9a90Mj5to82841gwY
aV3dpl1692Wkm//I7nNQmav2d5SgdOx+xKnxwbypUHGTw2RrhsFgFRX9RolX+ih8lnFkDXxJnZPC
DPdppydnYxf+xhuFalYY6NsKaQ4yhQoTUsp1l6r61M4ImkgYTZMf+P/MScg29AohG0AnMVAm1ELL
7XYQ5RDKvMzrav0OMRA/mq3CFcyn42bSvjVXDhIfcs2v6detlHXyqX5gu+zTZxUYHdTWPdyZxzUl
XwGd9j3283Ch730K5hVLrtI/VFMB1tnlblpNGq/TqIZrngkjLyL+i/AxTCjyUdd7TjNL/hvD8Xw8
vyJePAxOpmN94v1TgL+tkRAI6I3U+WgOh9IND62XXWPXxgtwvqOhKi3+VoSQL0DwLTYYqhLJuYZb
c7yb33yhNUuhVK46HnWMU29os7jOJZ60DqkUl6eCAdv3JEnyOzlNt6WLeOsbU2CUWCGiW2zlKyG3
gkAK3ks1VQUDiKTTG1mtK3mfAidIPjROPfHXxbsF2tphYYFDcQUd0vNIzBAyYW2qcFaKqgrBpOo5
8DYt2ScoQtgvvPlL7ybmtNOnfw+LGgmMW5Swboopr+TE4URiFpbXXTsa3eNbZsBZxPyDmCbZzRuf
NkYtW9FIzpsCucnLYh+dIvYVQ0F3A4XlQ3Z4sUqTSjR03SuhLDIbtay7Fj6VpZg7Z9XEDmvHmxQr
rwch9OcBblk8ziStKLpc9fRxSPvmF4KMt0yF+jNmTvHiNqYQO/aj6pGGfMBeJp+DV8tsDoasFPNE
X76B8fd5qwqdCP2YQgMwqOMl1TCFWb01QqpjD8bmFrt66SABNziCaBSyRso5edMDTv4OwPPC8m+d
D1wfJHZGH2/EdT8TH9H76rTxbMFLFuc9Swb328hK8OAN3//my+lq+nX+Zs+CLs2TxijR/gx1U5fw
OwwjkIjejfb4H/Zy/SuPAoWGl7I1uqq0YNve8EKPxKS/UR+YvdN9Vrje6C29P+RjnYQ6jvToFbm/
IeVTptkD7DcAFOykKXcTMuuVmTH5u29HOwoNxdZUYhgFXS4oTNfi8iMgNlVaBSg8zqy3lz6naoJz
UJ8L8PcgHYKW7aexNHYFEN2vap4C9t1Ho80vaPkHzpWDVGYmKodU19RSQZeyKthVlhcLZ5cnQmRZ
ztyMWvPaZC1G5G2XqJS2lRcfdqS9x0PtDF7AAHUn4vLPxRc6JG34Gb9otvPCJvebZnAwHGmnKskQ
O6JTBD5AoAfbAmGiFgqZFOw7Ra6TZKqLdjLF1j0qjiv9NRvSxlKbESXUKyVkROGg9dtenPLUM4O/
YwDcAMidpWRKHpj6v7kC+BVgBqhyB61NF1/gKMEaj4gtm0On3IpxvSEYpINOUxsPcILAxJUYqxVj
hN0/Wgp/VX8TWuVAcD+Uz+e6FO4plQlB3zEuvnqiMDSoPTLmP3+laJBcPQJakXeZ4V8cBVP92eXJ
2BPVdTzNA04VA7byFuM/WcfAJD4bz4KDabu7gHL0ZRCC8+DAt9hLBaGqgHgRfiebEQWWYtu6U464
lHDEUBZRjnbUJpETwIRQbwOQt+7k3DoWlOhlefgo1EjkKgkqmsfjhA+F2XrF/9CO85rgWRXeZPYi
kilNwkU4KmAFQq56GUtwb+PtbYyGPXGww697KWIQtR264SRkGMkcL2cUiBFleBLc4P0Mfc+FRnPH
ZPuEHPNA7aGKJIiJSszrCZbeHFh544J7wzwcFIRjhKrUj5OIyBYHH+A9hmJf8KgqfI+d7i0/IlTD
OOX/Tsyp7bmczHBlo/12zsrprF1Yvsx28IhJHIaTukyLLVFwvyucd+qGbUTSplqs1J6laF2Z4lC7
6syjm/XxKhyBSWBq4FP6dLpJ9RRooA/WxGD2XerMvw5JCy/7M1VW6bJILFh0h4Ch4XLaNJagsFu1
ewpuX7veCmsyfC244ePAiIebGRncLpA/ZSCdeQ/Q6uQJ86CxcWxsDg/QesbPLPwO/Bvva+oFpu8T
9FMvCNAoECH7vohEeaCxZHUfFMRMo0ScQlVgfQJmQpfbeX5XHvKIIrlOQbQ5kjOtr0+hzKtZmdPK
qCPEo+4o5dEZ4YY2vv0CJct7ZJ9HrmA3ewnRkcRLyMjOMs9NHW225HJtdD15U1ElRaqmlmPaQHIO
ejX62DcXdHXgrMxGq3K3zznBDhGJSnoaZ+CkDYF/AmAN/pMdbexh/R8zSSY/ed7gb7Opeb6CIJY3
wHoH+WCLg5ERRPrdQRsaL7tcdLVRCnkLXA4pomuv062Mgn1O6CboqmN8XpSzINv9PYuO12MejGPP
klInymifYr2W+QNJaQTpATdPjUYeURiBrK8Yqc2Sak4BhE+ZgtqE5eonGI8BTd0Sc03VZkjAFSe0
kp+4L4yhnSbdTFIoP0xyCLQWJTZiXUb2NMT71w7wJleQ9UXl+gWayFs2o6Psfb/tJOQiyyj7c/5N
EqlQv8OJfZiRdVSH+2vEuJB2FRISW70yLDckqt5KMdh7rOcVx87q489YMfniqgfzUQ4kxGDO46Zz
gkTjceYOxYxUr2g8ZAis4VZ7mGBtVG4tTGAwkL3+5d/LBGsOTt338KjxdAWsMMQmTqsJIoSx0L9I
pLptznLFUiCzqMGx1YZuaCG/xLdZnpWYMw9OtRe7lE/VaC0MCMyQFafMAlzHx8Ql14kT1B6uZjln
sYz8KHL34rrQZ9R9zg1FmDlPmkF55fRpR0wCkxD3s1WaKr/4jbcqzsErnY+w0I+G7I8cWc5Yazyk
vgXSD9oxtwA8GvLI4clJMG/iQWWeknCTzPtCfhsfd80d/jyJBlg53MdE+dpuSRhndsmmoDIOLYO+
4QN2jIjbEGko8kQK2WVEhMa2O1IyruYhRY6Dbm1mVQFNAZrNDnAInupRUaQQuIgvcRmtXKGRJcyd
GaCjLcb+Rc3CUv5/g/mhL7oJ7bOBvDKRwJN853NZZt0BTM7+MNDMMwpH5thNsifvlkTBuSQ0Hi+Z
/x1oKv26wS6nYK7fIv0WNCa8S7CK643Qs/OBZ8prp1TNIB29lrGIznfcwOzZR2LfWFivDTl/+C6i
12IPk5ZA+RM4Pc8dpu+q+5F5zZTNba/f6CHoM1Hfb4fvUATROZL4SCy1+t/HhSJeu0+VMD66+8Ng
sBJO7iuHgbaHe27fR4ROtdxwyk4S6gUCyx/dV+fMzwFN739LZ9gLKR+onO3m92Z+c0uBVVnkn3xF
bvD3MykurWc7KZ92IC+YbEAa2zRY9EZzI6/ejK5RI8zaeJB2JoyB7sTsQ0FB9/AoI5ASLsVSfVny
Avcvyf8UagvNiIegopOEDe02cljUG2k9XoU4CmToEL/qh0tBTD3y7PAFK0da8CrkkLlR31I/aMfL
I7x8Deiu/jPd5fHi5lXTRb0KeEVh/2YktztbOFZJcfwZmBNUQixcEWgzTXYoHyJ/ZtF1qGRhm59w
uboYgtpUKcwB0tAjHzoTe7SSxK7Yiu4QAOvGiwMC4+cI9/hIIBh7g4lCVRtl8xFZqRjGB6/KuFb6
l2XCWHHkFi/MX8yRnglNeFEisMX+B8s58iuYVeE9pmi/92lp79v0EZ94U1xZR22AiO+9tMy9xtKI
ysmERArz9JEGheNw2yYMvo2rru0gFcO4soZ0i613DQ4dvLoYPr6jfIyNa1FcRROYIUgrgxK6OZBE
fCvdYEjUMOfBSDHyqs+c25Gnq9M383E71fklW8H/roiLrCVo+itkd0qARcjHtxRhi1L5IbrlxnHZ
Bigd5NO1d5FSMaSqCcqAJQDCTx59LGFUUswxXX2beK2Tzp4YtQ3ct79cGxOR2qdxVFIJvHsTBXXt
96lUeNCBWFgGVrFohpMbNlyJ08klqADRcfj/vGmaHOyB9G9JOzvpgqsm/aYDvOICbOhTv3ArRsp5
5B8shvjARXjpPrh7RfnKXqexa1MIkEHOhsrqPc+Xu1QN02HpIpb293sL7gRkmyy5Y8S0r+5Gwu5U
Nlac2pA3C5WQAVQ3CYED//Jx9JzY0XJm5v4BoV8r/PNFeqWaxaOcU3ewCjBOVaXRBd3rEx0MlbIF
KmhtQVDiUrhzZ5+8Fg7e0+4oQVjS0sGeR7sSVaUUa62GzGchFrxurfg8u7CguXCj7S7DhCIZlvx0
EjnUHRFo4FcONKdLLjlkNvvV6gy68nBu+VwfpOps0ej/QBA48cwqI0yxyrPtHEsCTbpFEvvvU0FC
5It4onY4iD1uZJPn4y3EV3nE1u28ObTtSgg/AM/r8QLK4MfuTxXcrUa+2YpEG25/DQxuuJU2BW5O
eJvB/0sZhCa95bobVawY4tPHVVXaNE4c3Yw0iB+KO1+4DYjzDQF3UYQjyJLNq8XKkAp91L2wfkaE
KjquP2vbWBn+9ybAqiG9mJRx8fvKpAfi63SnF+Kf3eF9zyQTTX+I76c92z/ujAlQcMMogFptAtCY
qULgrttOk+k5DpnheSuiLvbzycaFvcSooWdNTJtpyT11QtcpLyY78dXZxKpKfGmvjWQGsIHhKN91
NrHVvKdGHOpkTLTEGRbiE6k60NOSpPQhNGzGkayPvdMx5VaXkDqcIHZoZoJfs5wiL+q5qY9a+ytF
oJ1SCkATUUR/pVQYKdHYhOEuw69WrDK84p2BBhUh/JW+ispR1if5HjxggCAU4Acwz3TmExNVhyVD
94YCgs4V++eJpV0TjuovRToPXM2woCFXfemC6wV7TuHm6pItcFaP63C8O2TttBIz90YzkOGIVbZe
mTlvZwvOKV19U0nsTqoXzn/IgMMQyKGE3EgbzRFsrXf2v8UFojUCk4FRveS29LzqIafrfdOI+GnC
G5SEMRo5fHINmYvMHKLdlANuRswgfPY9K6GBILCd9pwesKTrvDMQMpMAxNJOYZZLywMM05CQR+yY
Xa5Md2IM9B9XfkLr2aOy1jzlD/Vn05S/SmD5qpaSsWrO4ykx9zVnUAqitZ7WnlKXKBBK8ZeIk6Vw
SjUbFq42MnoVGZbedjR/qsxmkQBoRAJBUKwuyyG+0Qex9S82MRG49h3gpTv15xoXbAOH1GQPIAkK
zwr9xRC2aektiujXL72iAqwDbhaiIbCBRiBX1kgKtyfNASJ0j115ZpfzrEf5zhS/Z6cFbfuKXC6a
I8340HxgrYVKUqKMNfwCOwKr2DSmlAAoc0E8J2eeSutZKupSSKhb+eik/XCtSBo0/1sUt665/Nz9
aMGkRllBKbt8cKPO6n0L7igirwlPXm14cfTXLqLFpoF2y2vAyYy6ooWi5LuXG13rRXTB+zFYtZKd
PG2nYnV4DG6lNf1v1g4Vx157PjG5K8JipsRUB3UubBz4Ti3OZvbxz2biG/nq9obycGGINcP+Ssmj
V2tKsqimVcbuQumFUOciGOV9+j6CtgcnuhaphL5p92zmnXRcBEScSjSpSgXJ1DZkzeyOccE/c2G1
LnSTjI13c+0u8gDIBQlm7cNiovgO36dTHfCMgnGw3wX3uAmhNo/Wz9Kfk5nwJeErXv/M/Fb/XZXk
iL6aocf3sOcFiVHGpGZ3SEhlrALzY+oTMq14qJnU6DGhoiLCsBeB7BdK1CxKM4vnQgJkHts9yuq9
hZrbhvpArv36hcSdB46vhNZoStEb86nhF5rSCa67oWP0axrtaW5AKLDftm2fRh2sA1cSb4WGRPGM
+Jn1vtPr57GgJS7w6DdQtlcgr1JtsPxrlbWswNmX0AjXUZ3vTUY3pS9VYIRblgNo0tc2QhepfcyC
Pnfe0lnIPuE629byFhkbWUBX7aim4i5prsa66CNiFjLS9Y9iaaVPFdTlx9C+uHolopQXsvy76YAh
tvTc4Qx9wGGFee5vAOe8gpUL7QJf6jeeppyz46yFEyR3RHY1UvA8Fl2VJH/xDTpISSXvTjbim472
QHltnlgBQ4auI1ebyZMSaj11Cwzj5OgCidTFUU8ycWMUDWOkGM4DtTyhB79qL9zlsJeAqXqR1NGd
2+qvO5SqOyNI5y4zQulgQtthMBQrNwBDTpCm2jjvCLcN8WhfWZUZY1tQQkY8RQyrkhJfYpmSAQwZ
OsHoiIIvX+tNR4Z7qZWFHuO2xhK84QWUQvY4oQBABr9MjdUTiYI28euEIMrc6D5zid3dBn3ahJwR
t/WUCyr5vm4ZRRDZl3TavSO56v9o2HuBNvhBoB76DB6V3UZjlt1KGRIJ85GuWkIdjDP2oUyn3jyh
G82lkLRn6FtcXp6RbHKrMThOM3KrKS7MYDFjEj0SJTdF1Ux3ytnuCNdfAlGEyNgrSyyOLOZudqh6
ARyt9NAVTWsXsaZymPn5VhtOnfWknL8bJlWABolwrE8Ct2vBLsloxCMslFcMQoQALIU1XUQVfHAd
8xurWFbOVaN6Tz6gt0dPfVbJcjtTP9LrvSwgqZ8QaST6JnEjP/B13OEnyo+MDCRVmJgDbZ7kdVtr
sFNp8zR+wo9uzgHIPQU0TeLaa0Dt/eKi9NCoiER2Vp/kFCkaSPC9yNLKSg8ncq/f2JK/kBNPgZBU
31FrGfVgqOms3+9J3Go/lXSSUPVfzLTZZnZroeVi1cuRKXPzXHeAkI2q4nmSN31/0h1eFT8j5u9i
U2+4BxlL1CoVWaDrCaTQPsGjxyr4O+5h4+MKPeMKVxAdb+lkm9sQrtnC59XdVRc/ssMu7IS2pYMv
LwgGoMyjTAJTXq98x8yJggajJ8UiEtcEMwIbspDlt7pMuxsGPDx/mhlomyABxOQ5HNmJWkLQKjNI
gQeFPkfp315PS+/kUFT/oh/4unIkSik0dvb9u4LNJWQ8vJ5VOnCvpc/Whf/bPSwsBHWd2Q1WrIZj
NPQ2y0SulB3PD9A7VsQPkNNr3TOaBujk28CodC5S5mH1vfV7SEz2NM0CSMdWlqxyuz8cPCeZNHyS
/ICqgvlZWXYeMh31WCLljfWok5cQHzSX8fKqHKF0iTS+wHJJVgGysazhTcr458x0yIRsVKR0LCmJ
EVdax/UzPu+wyGA6Wc7WTlxQqovWjYDmCiUyijtZvTIs4H7hDR9SfICASKEj8l60gRtxsnIzfxPD
a6LqV73D9TdcXfa/DaKZl5f3jYcGbnn8roJjx0zSKVpQWLXVDJEpDwThGQBL8jHAW2I5t/Q37uQJ
D6GmciODYHqM9MXalaz9jo5dEDYPsNukIXsEAega8YzOInsB5x5gxyhKEn10YKoPaucia0cRv32K
ZpgfjrR6yi9yahw+BZLkX6DHO3Gj98CKbpCCOvRF1DZuG42714g2BAytfdD3SrJt/T/0EKuVX/RW
9MUWRqkY/cTZooG9ODD3xCGbh9rP5KVB7yY5vD5zxem44xfkocp7/WcVk5P+3ZXU/yPtq3PK+Be0
aXFM0DIHhG3UTnGbspmdX4oHWmZeMqaCO7M2G15o9eJYbkUTYs0XgAGp9sFZHYo10GenOpazUjJV
MxY7V/MIAIFhR5lUBYLNVY1K2HR2bzsIaN+fS9ecWstdo3k09dR8ReDYfpIKWhaORoe9O14LJf7P
xsxo2FSL6EsaUX1Q85adNt+w4/ZVcHaOvZgyBFNcgjba+Btt6iHnGmzthnI1yzaBu/NHCNyw1Qc7
lktbTsfsjo0iAPwH1NnwIM85Opd4SL9Ojvth6aYsLSU6MIY4Epf7KKX5dDbS0rcSXhq8mk1kQTUq
G0sTtJyfcYm5iRu+zgbTXrcI1z+ikWqR8ohHQIuxxGubIAs7a95rurJHPD7/zkHNuCR5L19r8oQT
QGMo8lKdVCRec8d0kTNy9GdeCXm4A4ZGmktKeoFA0j2gmwmtivTL4A4ubEiS6g0mxl3Hv3J/oRlG
a8U0X/Yv7ZM8IYwgB/r53DBG8RazUo4aBuuro+31jSngLHNVM+rS81e+OK+oCvt0oQk3fjWtKqJt
wY/axUu0vnHtEP3U2KBFw9K4L17mdCRyOkDE2uHt6Wd0IW0iBRpHVlrirwqqrfbzVqxgbHgpeQ/A
XyeyWQsv584cwnjN82ZbBlMoKkn6P5wAdFeL5ABhlf/JXUCzFruiZXuEU2kU04Ti4XQv0R1dn9cj
WBlFRppb7qCrt6uSEIRvGbHFk+2oJfNk7s+pecX4pn+YoESroijYSzYc/dEM9HRjhMu9HfKC8d0W
uepodqcSCqVo3SedXrQ6ArEtrj6QChpDa3W4xpIeb4PVhmXNDhfpU3tXxuElQlsSvKxK1aDuRc9i
wI9FUxAiUQxop9PMvKKBhDHyt0kTKtgwlfkh4yLVDjzqiQCPd9G1SrTusL5MGBS1kOIvjBoY3eh5
0LyjAjmHZgFzzchETJFg7qRi2MhQ9LmvBgxXWas16zZEIrN6ZeMPEVIwG+rYOW5SJiAeb1u5Gd0C
xKsCNFqXIFVhhB5CivboFv86UDgPKSDyPdPOoMrxdnCNthzp9uXeoYklDQ+LMlcy8QfxSPiOBxBV
cNSodEfPTZZwsOsTPZwcruY/IE2QkOUJ4+1wblyMQBU4oAJoGwPljPb3+GZW0pZYUzZhZQgyVL3b
stSOqG2ULj9j7o3uzLX81Vl/JM5U4bhvtGR+FocPCkN+q1ynltVLrSH/Dc8wNMYcGJF4oVA9E3u5
ukL7SR/xwKXLS1xwb3XbCS+J3W4A+X7/AJb1BKPeMBaxF1C88uxCErr5osNuC+0wjEgvx0X+mLmy
bf0NkO/Uj8mNJwnv+di1o3bKx38akcU0LzYWAwsq/zmzesuxuhqiEiWLffVkPkmOoiaB1+2nJxiG
Ym1Fgn1pPE6cm4cEhm9rI2iz3cnBdmojv3LcX4mJIkPAJMyMh6ausv4BOFcJvxmvAf79PJ4MOlZ9
LemVjPzIdhLPs3ZrlJ8DEFHIknkOX37DP1nFjc83rDO7I0PgYJbK155Gp/5x4P2YwbGnMp91Sqyv
l7zTCu8hytS1Q+TnVHRrA8dpDP/oD0aTHeFFFPt74oEXhynG4DMO3BwxO838S0EpYtymnzjZwQQT
DGWsGnctl3ZJ3KFSAmrBMPhzKOzjDtYWWeFqEETQSFAHDAqcd+AvpE45r6pU5dVjce4Fzw0F4d2s
9ABqic4p4At+MGvnV31BYl5ng0avUNOifVqBqbdwaNaNw6zLZtUf6m3NsTB3h8BoN39P7go52zYo
C3ma/sQ9Kcbk8VCApLSRExCgcFsXAMF/tOMPsaPJYSikMWzqVqyZutMOgHb0rGGwGj7gBqlqraFT
+7gUcKXkG0VdBJijILUu+0pneAco9cGr9nf5foroqEFN6UpPJv5mCr40NDlxlsnXMFxw+HwoXUx4
hmFZBEXHocW47VHHPBysG+Cn/NoL75ks/pCpvgLJrWmkEIvDoTwHZ3R6ZVgCzkZhGuxVTaARAW9l
34xWwi3KPShYuGE5Y9jrQJHg3l8mFxbs18WHHAzQdjbnQFoGikRP8l/bmp7+2yMyRy/INFzvLLyh
/KP2D9hsK4LRPXEhqlWY+yhWrjq4Fs6UIJ/5jaPjntOfevk7mxcFZ0FaeqzTsk28tHt9MSNpsztJ
8v3q+y89uMkIBX3MWIobYdWUF0zH85Sui92IkUSuVoII9gmQw8V67FsibS2lX9nlCAkja9IDh8iS
bOX9sAGE0h2Qu9VWdkx59fVOgquB1VcVEnAp+MQjt2Vkte80dv+S7hjyI8TqB2eoZCxkBTpF5SgV
O5BtL2/dErxhl6cGwkJfsdzc8GPdRN+rRa2SFtn51IldPcKB91VEJwnDTLl1N+flIkApXKR2MwWU
Y0J5CwM+x3r6Mx11UKrewTdDGlNZQNwTP+yO4q3hGoM2WcETiinFEuK4hiXb8HYpTBllJFIcx2/b
dZSWejcHy0HVQZUCK4qqK/krXtZ6cNafgKQ1j2ZJdgXHOe/sfcz1Xsu4Z8r5paR79o4tTe8oqUdH
SjSINtI13GrsF7UepdrMa/builcdP1GM83Up3Ps22LTKOAHJ5YV9Bld8f30hGP+QPDL5sAfBjZRy
z0EyjVsXMSoIIS68uPwMMqWI8E9T8254fQqr4GZ8aMN6xieMmNRFr+GpVJdMK9pHIUGJz+GndaQQ
GNizXEVY99TIQC3PgKVhg5Q2QabrZZL0eY8lK3W7egjKa0uYXzgBnLHBk+6FHpdLuFn6fXRzaegy
RpyiVbaGdrurkdrlnKbZ0ZWHdQaPgYNI3GAAGv4HFPB3gv4O299Y/lGvMYiROfMN+dLQmMoFSlBC
1wR4C9DhA+yTI+//uyv5oXfsyjlTEFsu0Uy0avoOSPL+Ew/D9ENURFbxzlKc1xos0kWkXM7Kk7q6
7+xX0/iNFZBHZfC4H6/qBDHMrxR3Jdq8qIGQzyzOjHk3Os9nOCxZxmtbYOCqXaOR3IUXyO5BXN+G
8/60ISjzJLWBLc4L5IIjQFP0Sb0w8TXcjLKhSr0aq8SHaX81BTVAqIGKEQ0xFT08eyGlKWnXegtf
hZCbEkRc+IPhiO7Xcsw+byK5eVcVCyxmx+WE7qMbMTEKfhROFRgA3UpECmUj6hmsjnZRbX2Xl4Wl
vwHlAGIswbZDvFzL1v8jTBSP2p2RrMCy36qmLQpzBXpwxBypuX3rq+CRvbwrDMtLJh3DgByrOrFs
z+Vb2szwxqWuVxjHK+VqaCHzFOMg/DdUmroAlQJBHAYCLSWQrXxllfjpjXOsRKcdmXBSm5u+IOvp
pB3SKwmr8CC9vua+aqnKiBRmxz63RltehoX0U9AcL0PFUUqFfgv2MoyIf59s44beZjbzWFDF4XFO
UhCIGmlizlFBBzAGb5B7IwdSv/lk3k5F2WytYSKL/2MiVKpXi0h47Ro6AhRRuQAy1MKA1oGZi61b
i6GjZeQe0ohqxaMmAcVGR3vsW16FimRAMQ4a6mRh9d5e/RbW1hFet/vzpKPFZlTB8fvf2ee6dOY2
LIYmobRF731/yQCQoBTifPP2J00tWtuBac8YAUMaUxfNOuOFzX0MzfVyVchduxncsb5I+hHnxq/g
l8BFkBXybNSGuRk19iyBZWU0vNdCaw9IZikQI5dJu+tGPF1sTn0fuPicx3ftdl4pYS5FncnUzchX
UGde0iM46I+ZvKOD6ZgkTJarLqgpfkUpE/osjYC8dB+nZ2iZ/eqb4OMnlbZSKN0G6HCzEKwPdlPo
MqlVLmoQP+tan7xAQFawPheiJta9vhnbbyFP3xYV+hiNxE7LCWZVO+n0jR3lGyuoeHCjFyJUzSIt
jmNiTaC6eJhW/cOIiGciy96sWYQ5ot+H1sB8fBMQLromnj+g7BtAC0LWUO3JZ0lY6MaORhD/ezqB
PJIRIcrEePoBhgj3MkbO3LFzH0+I/ig9M6mmDrOYi7doaUHpf2JULxFIo04XEJNad0V31GrkLz/P
TZSTip0hFgg73wFda5hLw3ghMgqZHY6n46J/982LWOCfqro5CL9agpbgt+oCMaFUOvZSzM+0tbIO
SfXzW69H6O4GHoc37FkofKI2q3OKKbN0h9cvQzEf81uvdgZjiDt6z5QkGJTyFYXvKfK2RvQ6BPS3
qNljm2d8y7o1jwBrmjDqFd+GBvca4ii8HcnLjy9fbl6MaG4zZ5H5OkOxf1rnVkDdJlPWbh70mBob
5Ofz1TFD/sY/1+RB+ZMCSmDZppkM25PkpYixxbx/yFx8ZoZdyFdokRE1dBzOE4ggTTFeBCkDldDr
kLe73pWLCzNsmazv0gU1KCp1R7FC3FZewekKfacRiQx4AnchyfUkFEAmfRtjVUmp+8PqjE7xDz2L
pQpTJHVkF3JKYwAG8jd5qDYKnHl/OXoiySQnSJ2ZMWA+eLJCJaCs/J8Y2n8MzArY3Kw8Vrn0I///
S6Fmzf2tKZGMPDHstAfR0ewQq8g3uQ/UzS7NfTWP5ynFnegzhL/Avqu+bfr4bo80MHql1Qd2PzFS
cSYl5MUS5yipbZGewRmsIsN0EkypdWNVTVHwMWpdAJOgTkFWAu3cnhVjjn65j4danCjHZRWPakIy
CbrU8+0VWTWioc5kBAcaZmxGfaGIpfyyUxKZFXDMwQkwah6wtBeEFhrhphfOd7yWHuAjairn/h0R
yWKbd760SDxOhNs7Jg/8rnF1dcOSjbAO/sQDSFcZC6hk6hDJbGlDIdbVeMl9PX25+PDfYqygNnO4
Q/CUPVekEail8u+RNOMtJWMaMNu5gH6sGBInE+3BhBA1NrzLM8FwayvDTQA/g7Z2EiR3YELDwJy/
3V7KGEYrAlAPTZlTBh80l7bWbEx/BHFDiBkhBBAwvI1sSNBmnA7wSsWUkQ8QQIBZq//711CEWIr7
OFmGKOGBUGolYPBeda50MB1GjuKbuCs4llQpNr2EaEU/vXZK9T3lYU7fCtoPdf8SMDF4TmC42bdF
14w9IwhEHaiqgbj6vMMERlwrZJRU3mUNSYYK7Or3bKO7xLc9UzGfQiNJgfYBiXwuFUdNWx3Ogi6j
H9mrcHAbA3UOORB9Z95xPl1HV327/ehM8oFpOH/nH+/iYhzYbk5m8HdkYNc66obvFaspHEzHAlG+
+iva7R6gy0NRdaF9J70eyBgy7ndAgmC+uU9/Kt2qWW77Cez7Gzf9Ky3lTRX2OWtUEsk2eZ8m4RVw
WrsfhSnvSBUzKhq7Onn+qOk/EakD04bK+lwlg19sddcAREwbSzpRU771Rh4tb/qqCPZsKnAPOa/i
UbglL+5HWUEC7IezAaY8TPeC5WvFV4cKEQfqHjJQqtCtrjQykDU12/c50sDaP/7ITFKfZ3HDzRUm
/qbJEc+8BHUmyA1HxZ7YrAZM5T5x4/rfwPKmRqmC4fAFBtOnpFQCKnI1ffgjW9OltHbTERoZLxk2
KtFN9npmaPwIZ+HZAyiO5O946p1iOuNkyBLGAIvMm2CgY7lCelHWgxROyCsAf07UkzanIlX5/BXr
HFfP/OgC3Bs9s1ZCTqcNVGUYlJwBp8P4kRN+EGdqHO9JQzEBq1zEFxqsfyeRhLJBDXKsyRKZXvJv
eMX1GZlThf0DN43dIjdCkoBQUubtBtaMROCj8Zd1UZsQ0gDUgBvTkWkGERpJjU20N9Zw7euBd1Gu
65o2PAyV9hE75m9naHcpn8tzYowKVeREt2dW8ByOkG1Nt9865Qez+WfDn/htK5xLch1Qkq4av0II
5FarI1Efm8EB336PdPP734a/LaKPZetgazX+orWHgsYNUDXuiXo5h9lAP4vyKO4wsYo1If4ARQu6
bh7ZyKqkFjRimKy0FeSmqPp9+NJ+hDGRThk4icccnXouDTnTgdFeTEAG5WKuktWcGtoLos78i/A1
oLw7NL3X+fMnFPFBvCLCPu93SUd3SUQw7/rcqQLqfLu71CEATD4mF1XHOa/2+NSHtOmWkWWMVzqw
nC1R2zZGCK5EDwRFDq0HqE7Ed8W++z8pn6KJ9IBTbqHcetHyR/j70vZPUqYx/kSK1JbnFvFaXmFW
DTqGMzgtTDldByKo3sfgfLXDbP8dI0WhVnBC73biujysM2f3L5yqX2qlpXhMyYTryE9z1qkKWfSz
sQg2i3kc3ogQ5UtDQs/7hiOokOu7wVa/apdaoJeb3OYvJgNX4heMALZZrMeZ6E460x4ifU0WYzQE
Yi5uOKZ5ZYqPDZWj4Rlvp+mtldJcSYeASfAIu/FxqVHhPtylZH2ZKl5AVpyFNTdBoaL6Kb3D49dB
rJTKCKm2MFnS4pCtHVZl5kzUw8YnB3Tl/MmFt0NondHet6+IIlZdZ+qnMC9L086xGQOK0Qv7U9yV
K6GOHM81vEIMiSWtyRA7divjacB7es7MiQQrMvOpArKcbEsFhlPocWYpAMqQ+zWkoBH9uMDW/quS
Iq6IrSnjmmni8p2WvS6J35SShLPiAoonRCbln5INGv3qb8agm/UnAAY6Qd8NIkdfOZaHwA4u8p4+
3nJ6EVVr/aw7njdNKaBOqVFrfNF5iwmezFOI1ru800mSiJQijnLwFQrJcPnRHY3vpxAiCRsRq1Ys
/TX/O4nW/+8FjfARJw/9ja09FcbIGCWngIrHDK6f/wBp/l8MyDYvJyuJ9O8sy40GxJ0kyM37wIcS
Uik0nb91FiJmFY8epDwk//fJcnR1S+7EtrYfb0RwBOjq4NFV/fB3J831s7XYtpay8ww6G3qmim8s
PtpsY6kCgJ9QICHgSKP9yfsHcqzdfqD+DjbP+xUHFiLcujWxyaFZEdol+WxBFJl07umkHiakM3O2
c/n4rJ9HAZAfXC3HCnirbVzC/4JZgodgFQ1PWVaLngLg+rbWZ2w1usAQr0rOAKCnrWHwF9CXCCNO
Iqzbt85c2Bn2D2Gew9qCLfffdp/FfyIxpD6whjxKBdtGm99P2bNyVCNggHx2JPVKdegYyoG26mTU
kmTcBcndh9FsEBB8YoFzfWgpF8d6fhsqakxoGJQ3JH6kA1sIgXhmfS3HeTWbd334m+fDIMvPOxPF
Ryug4I0t0GEZL3OqAp+aw/yAM1lJMrvI3pssvf5Ngrs5azo0wu5olngVkyke0dIHYf9Dy7zcjQv5
FGfC2cE+b/ljeoBb6tl9QxrvX2vWsJ1DoXpPs8CP+U1Pm9DXgz9gl3Lgq+XGJX5dtGyB7pGoK8UE
iIHA6i8AKbN9DyBXf3+m6a1VKiFvQvTDguI1NfSSz+GS0ey7Ak/9+JXBoAlpGZwIrQ77SOmuP5tv
edvVH1ZrVOh/G03sYBwm3eU6GKIy8qdCn/yOt8ws0sDMGexhSbX1Vfc/QcJdKE0PzLUdBh3XCSR4
WgA1FRjvZOti33yK4rd8Er1exxs9jnvYB41yOES/8Gyk2y9uZwyueZSo8e4D8hS6vW+1BxVqilO7
Mer0NQVdAmjusjfRXd2+WFflWDvEzsNQxXW2d4z+/Ah6rwiAdVgiDWlrXeYdivx12yLRxOJqdSeY
tQBNIamsIhmtB1bmUKpB4brRef6i2pT77i1osN8cdgcz4R3vyjzzg5155NMUHk7QJaxbb6nMb7Yj
1ZVeX0ymzC7nyO/5df+sH9jUgu/8bG+INs2N2eOBdMSYYP+YqQF0RWdi8k7QDAMN7e2PMlFKdZil
7eGQ28QvmNZQvlkc0plxKxebK2JWdf66XU+jX+y8hRWGK2zGuobwtvPbMNKPNBHMziXhnDHNOV3/
AZHocsUA2nwD/SEINnbbngfbIIPwkkhUEmdfU3AOyK1OLdEdxuMZkLRW379fWGoBQngtP14DIVIA
PMTkWofI+rDu9phh/bwwU+6CMRE65Go9MwcDKcw1fnM2NAiQApGukIx5J9BGQDRiUganA2FU/O+j
n2xnAJkAVkABOPXiuotqd9L4+f0xlqv0U5LJwwa1iF82I85wc0x/1b7VLrx4Xo+zed5NmsLltzwu
eNjMLUQdvchoOI22JMiUjXRUhMTeYkfCQ4GUb2R0rBbA2nfh59NTz4NBrmNwHoCcGivpPfWvShMZ
LUtgS0vzWMOM1ClBorhy9WwbzB7r+/kc24xkOf4EdrRnLIIlAs3w0NxBOauWIRUrrmCiUFZ63Jt4
EbbzwcjlQgHIXuTis1g4v7C3EEE6ahWnOlzaZK2AueqKgk4bq5HECyyRrTlUyxBaEUmKLulya7hZ
ahseJEVqvtjbSTzqJy6EHoGuMchMeMyiW1TO7h3K+QLg0xE1ZDaM0z/2+gJ1Z4GnVH6IHSOLLekZ
rs+IpEPiGr3jDIWj8F+lFxoaDkFsD89XlAkrhy+fVF+637fF7p8CB+DCKu0doNwbQhxgm07IGHsD
kPyJudttbK+UXh9Otu37dgWtc9uHnULZrWJ6pMu04vzWMEw1ou13wrB/t2GqZz7Us7B0SO87RdDL
YQsZszLm0XI+gc7Ju8dfwNWsm07rmXO6G7jHnoU5MvaYjOkKsZ1lYIn6PVPARQvYiEckP9BeL2LO
pQQ9I+aszk+kJdtVjcz3D3n51WgL/EGryhC/y2CwJoHAx0pVyA+F1aygLNs1nDhMZBjiDh8Hf0FF
WAR5C3SR+VrIPli2B+hKKCTkFos1wEy2ZbU8xOCwyDONH54ryuan/FVHaAZyvUT70k+1hRiRGIKo
OmCnm3MGYpw5TBCE3PR2WVQNrUZ1mPKL54xMDGzAPnwC1tvQaZyZWS4crx3SC/uraWaUs7+WJWB1
UNZY9O4T08J447cxxR3EC4LMvKW/ICD7XOcslJZ+Ktd95iB2kVFdM8uuXhQ1oCbTcfR2iSE0U5vP
hkpjvGX7Bn1j4VvrdUvIH9xMzJBBYP2z7xEckv0wjwSDmOkIei7wWueIiFqIKCIe2aeu8w3/mTOm
a8HmMC83S0ekAk5E4me2pah/85YLXl2lFo0MrpwFNXk7IiQGryXWrx6IGYTMcwUcODtjqNAPqMwS
s5pE7mERww2f6L/9yGXVSBj6CSeDRBGEbDMqn2V6FN86J1xMS2EZIuU/7M9fYeMpPlGUixPsRWq0
oaJ4YyizrtLF0XWLnWUUYlWqAFSP2wmdhK/PsSM+IV2KvSNHHAxFE2C6/ScfGydp7vhWdSg4us0a
D+Kd4p7U9S2hlZ6KlCxXIW+aCFBINvDYANnvkXbe9ZUaF9QrU3+/WOARgf/5G7JdKAL6rFfOnnRo
h++ITtVxVLiwi1mXCitqIMZrtAHXMxEOvWYp8zFO3lUNLBNOe476wVperiyxzFzlwFgl0KDWT+/n
2qxEYl9bXrX6qgpbXEgv1Kj33B/N4gbyQyI1C+IL2GPjfh4gWOWSVfjuOQSF8jXp+Dds19iTP0NC
BwjSy3mzXXmOXAXAOVjgTXlNBwdSaePqK6mDn4PuaQAzbQmAEDXZQJmeRHx2J/cJhYmriZpZKR1I
2am1hnXeRLFQXRib+HmijJGc7QhriFSt+T9QYOku1eF2ApXtQg0zfGEp1d4DJmIUs91gj94CgUSv
jFYCwpY/Sypb0mh2HdRbVUq/D5v713sZsMNrsiYjn8xGXXWHNDPed9aa0oz/1Eh1B3T2BAFDpxDC
+JQxhOsMuVs+C/iAeIl/BaX+ztnHlGkrJNJh20AO6Gsm5ci7ZSHkhfccZb81lxgFm6/BHPlhiR0b
CdyRfCtvtSuI8Hu4UL16MqbwPIkELR3JN3jBfWWz3mfXkHv0u73MB+kZAmFchGxCa1F7iTXX5xD0
oPRHxYJf1IaHhQPu0Jzd/ibMs+knycuNLOccgoZcNdiQOayEhe7xTXdGH3Ne2m54yCzB08+174bJ
GOtm5s66jtAgeQlXpHsX5+6sXdZxqBs9xGHRD6tTmjmU60B41Tptdx4ARst7QpRtHR1hVnQr77qH
KKGrq3qrOiX5u5dBJsjNGUO/Zmaldjfaevi2uRItxYKBl0I5EqC22Z+KQM/PNcnMtVMXn1eRTNu3
Q8eTZm8TC0yzUjf6Cb4LwchGDsPMhBg37arv0HECce63fNhfPZRIndSFdOCOiMUBNGtIQxzWjFFJ
HgNNmROOy+6dycYATcUHFrm5vZHgaGEwxnHbmpDOoZ/k4qSQvtAOekMU94ZCWrh+pB1oZE+2kR4h
CdZ7SGJNM28hd8NapVVYHZoSur93TJSQny4L7PaJnBESyIhgvElNDsJvKiZIduScGhQXEVJRx9b9
ByoWKfKBza4jZSGSIVGHjp4kHTkHaCgznLEknjq6w9I3RsSJVsVNpY1l5Udkx9oQgLK1mizmo1Tv
ybvXvrwvQ2xOrKmG6AhiKxTec9Dw3BqvVsvRqu/Rg82/I5dJ7UXJxLyslfDkTXdebvo5lSO++k4a
Umte5Aee8nau8vmBILGAu26+1k8miw3LT6pfol9B6Bk9klVe6oAZcjcicOxlu0owA0um8syNzz5e
/1RLc30ofVoJ7jQhIa32hZjee7gO5xHTNoYVORC1neSFskn1o2VxKlXqpHX8tMx4oKUyRUbzAzB4
CWDXOUZitlz5yYDtVNyyjqKUcw/Ewx++p6+aOureByPtxxzBuPq+mj//2c2fWYNxzDxDcnpnNtbr
NblCm6wgHDh1kk3oU3nfyIUJbG6bDBb7iOAsBfBCU5lfTsYcAk9zCM9gpotceYBWhIYCyJEvOWu9
cmwQ4M9hfo7SsZTFDRbTPRh7KPYk+0n9NQyH76fJMKnXbt/IITEMCdkLmrlNT3niKtvM8SemCKja
fkdihEUAtpDXzsAbrYoQclYnICMcvrd98DWy4iI7naeenQ15+PwaDnAscBzkSqJkXJWE6Xn3Hfdf
m3kTJ2kC1F/3v6o0LpL0R5+xm/UQf7VHktemOvSGpnCPIwdAxMEgs1xRvT5gCziysxJjHE8tqaNW
lc3gp4UFqbhEyocgx/hqFX7zG2VcAspULj5JXmwH7zDJoRaNg1HIcq9Jj/fj5qvCzz9Zn/5fbbll
wZDHhTVo1RpOz+RAnUUk/4PAX3Xg96uX3NmVA7TFeUVA6skns6dtP8Diu5BxSkKAcD5YJ5A/zVBJ
Aef9m5mK/QgLnZjbjxYcgNcTQbjT8vKpdTezwbcsOs+q647PzKcf6DHfB+vhgZ5zNFwanVFkRH6x
ae7NrSWlkqyn4wA39oN1zGJpbTb59HY+zU7tov0JAUAfQhqwKmPgaAmQoLYg3UtVK5SM8obLMd53
4mC3QOFrM5O9A/PASKB42FQGF1pYYcUoKkYSAEvTyqWan+5nwEp8VEAMRndn4W9zW3MIMl78tDDg
FIqpsjcOe48oucwwxq+BEkJbmnGgNfiz/We0ldYlv5d7ubngtjFm7jhn+jTN3/+pj+yiDtSTisiO
6WRIYgHTuLUJQ8JxJ4Mevm8PeGwdu/zAS1reO5PT8SM1O17sSNbpd8J2WWgLYwV6Mnjnw66uCfoS
Xt6+nlUKN9tVKf8KV3bk1WWIDk4gJc2Ce1cbggRygJUJ39RuHrmod63mJoBVYEK/Jcsf6QntevbE
3GWzsHnERxCDqIExCH1dNY11/yaoLU7fdUYA8aCEU4/6eIBXvvz5g4XAegC/SOw8nyNVbrLUMl/N
c444C8dB/YL0T1yUPZjW0YMIhnKpptk3TZIfVmvSutzdHpeNKzsQGsSCGABPgqpWT854EjSt8nba
SLDoZO1OhQkUwrU4/iMOLG31iUzD+ukdYHGw+vyhG3DkC8ia4YeqqQLXhhDn6H0/GhYOhP1LW/N5
Lu23NM6Qy8tqmr/hTy6sm+fL+iqZqSlDYzyPR84szwv1Yj2YshtTo9NJE1iV5zzWAN2QTNt7cQ3J
w/KOjL49RFmcHbrOwpQilbP06Y/1H2WKxwKWSQ6hYHxzhEgyeAqZ8/ZWJg7K75QE2bvNSgyG/dPr
+3IxE9otSBlkkzFoZXYaEtZ4lCwcFV/7Zesdo6izLTfMP7aIDcxlm277HRLmyh1xIP259ZHS66tl
WtHqsTSfYsc4/ogbdWGqTkPICogVVu9fFLMIr2PP+lxkLLT8/VNez4LAp3o2Vh1fHaVVMXokalZj
a9uIXc7NAEFI6NK/gCjASF2/ayBt3LiUpHLWLyl/gq5mYIFb7Z+UfpHJI9y9OkGVlsQO8nqgDNPt
IeiruE/zhYIXC13loVzWWmKwOrHzBX7u7oSsugGT/lndjyo1psghuVl/f8CapY+E85Dw9ZZbySMv
8IFjV6dguWtlY/B/0gKoGd+CgLeJ8jiZ+/ICxTLZb79Ch8NL8UyuCEDVbxjapU3znae3Q8owZz6P
mErYvNlh45pugk0K4QG5dZm5smcojN/0ojxvvJDnVC6ZG5aOh1vf+lF3gVYnQxbDYtpXC2p03Prp
7p82JFidqm+x6c+dAGFuGkm8QYUNvY5mX0ZWk6nlDFjL0a6SQRS4S0LEkrx5nB9CH0SDYLKYYV3d
C/LFeLGIdYDPug0wW8dlfqj/lpq7uQUnxD0TWzelD8DXzYgCBiuP3JYL/z890d35KQkcQQt4K4r0
Uv1WBm8Xmj+2Nrcj44zvKgVbq+JwmjFH3NhpwAFimDx5cazKKrQViDV+59rX0pVaXQ0rdpOZVFj9
sbeydGfC4/IJHvK/e5SHsWMZuDKYuRIJwkRF3MhxxLwg0CiG7AssIec3eUaD5WqyZrEWlLBrMkXi
q7ge4sNhT08d0RDsuFdm4w6+KpbvfCgG7OidUresVZNzOQ0fCACT3i2fhlq1OKT/Pz7UFPrfk4Nj
bw5pOY19o4DD+NdP+CdYqs0BR/QAqYIXcaUte1bCTqzn45bQztKY+m1F1VEjNwoBJBgFWBZpkBjW
ONnqGL+J2jAKz96pgVuIxjPuTsl5bjuTvFnVnAbRx1rKpJkAFpITNldRpMsO65eY8Qd183ci47Sd
FwdOBFrJOGSAJDsFOV6opA3XAKA1pDCwLdUIcDBmVyFfRrz97p37uHOyJTn8t7i8xhjfB8svPSEC
NJSQR+Eo783D8ZlsPIug376G10YgPwir1cR+LCg3UZNxxfIsh6785BdosJYWq5QphOC/6x826w7G
Og4/VAURWSxbxdh7N57fbVvwr7wgZFjS73JgaWSVFgkxkg1pYPnTQea/fwMY5+D9ynrBgR4tXXR8
etWeyt1iGJ5mdDzDarXiFk3BfRaSPH+Xkxkm0iOKS3WxyT10Gvg6VyONQXsPeXF+q0hLd1P/I0Hp
M920Q7axUNXZh/mnl1IVQKGAvGOVqlKVkPS3opT3uFU/l2vRU1MR+5sxGjgyIqGEbmez3Aw2e2Vy
HTZkOusXXNd4sc9ReCYlxYOb0E0DOk6EjQlbAvEUKejOd1edq6ut6aucRJKvE19p5cY3ERRXPBK4
9pwEgjTt24GrSra+Zya8fTn4FBL8Ra90qr0WPxNu2Li7hW4oQZ37uroj4UD13RBjpSAa7s10Edhc
di69JTTBhTTf6TBwkh8k+3CqgOzXaUteTD2iBhIJ9b3Y7c5huzxsAtJW8b98xmUkssHcyXBDD6ij
w3lXWxmnwwysfTT0Pt8axegHt15thj3ThvzwGHtCbwv6tIVkwkX3NmewHA+ty90x3p/AC5YyOGzi
j4A/Y0q0aD2qJhf8G7ZiI1k5tnBZsoYyza5qNvBumqyYZ53p9J0O4xXmnXJoCi4gp/wt+ulf9k8b
Rq9XGZSsUX0aRXOBFlB/t+wT6dbkEKi2yA+YmzfJTGEZ4Wl7oFuB+JUKzHil5tUW2MD8OVf9DGEC
lzJ1Cz5CBzlzSZA8HiC4Symh4HUAwVvgRa47iY/d7BVQ8cN2i9t8qTe0asc992NF+MX1CWcOtnZX
KUoMMk/wxbY8HDwQoLbdPhjWRI2FLNJF5ih2RqB9uQbZdb73X1u/VoQitBnJczhvQ0i6qo7vZQWZ
oOswonKkxG82HDdt2OollOfJf32jYvZA7tY/FEYgIQyZ1mZ3ombIs6BDgyvsyFhIQGtImOKm6Ro4
8TY9pTLx9M/fLptjnijTsmJQBYAFjpmEuUm0YasuQqNvQzN5PgTiW90CgeASktwG4yI8fTemu1cx
3Nm3r2M1AbJ3oA7uHAbn14+jSy3ZQAYz+ETXS8RrJI02S7A1TUjEzTV0dKpRrEVWCU52K47BG4Pw
zziaMgGOMXiVhHg+xQP6YRC1ImNBz44L18FSRxQyuPZmCqx9OHPRpKZ8ZR2jj4ouiNReKu4vAxil
rtPw08V7zd9wu5Vs8/vOBStpW1y5JhHmIX4qRXtjjvmY4/i2z8hxAf8GWNYM2B4bhFi5ZlcvkEMd
8MdCBxdWKmZkj+uvwsuMQrcSCVS6hO11ZWkphlx7v0+rIgrC2YeRZ+F9MDq5iYLd9KAVESqjU8F8
Gos5xbKHkHxnWvoL3gRVFIhrH/OfGNHz8FARzkFUsVwy8D6QjYLWKdI6bkMC7NH+Yqfz2iJd+DxE
PfP6ntl4TFnrDuWG54HbiWU3PXhTVQcWJr3FtyxZjfVoEp5NLrUTMYDHUO/D4tWiWvDLWNcelUO8
HSxZFZ3oIwHdOoM5MVzN6Qgc6f4b4+/RRbjnOTi1axGCsk12g6Wlg0l5LR8MXE2K13sgjp2PsP67
kZkMNozRRZMVhjwF74ZwneZocLo/sfnccTL/Z5D5YaiwDoDZH0bN/KUl/2+Lqfcb+CF+Yq+wDaqz
WBoj2z8KAeiavlkzjNn/0zpsS973s/quTkIzZuTIYRYuqf3UDd07KJaTUy8F0jm9u+7IfhVg9fJU
1gJdoaeji+aEEclPgi3aE93ANsIJC4bVXuAbUJs4W8bK9lO210fjlhMxAuPLBSvJSn8TA1AldXgF
JcHwaVgWCydSpyY00kJ81XepbFP4nFxxTGWVW9vn7Wylh4cwdPT9w4slbC3TG5PLrUypiq6oPjLs
Tmfj9xVttY5YSaWGxI0yIPx25N1keNKKJDeB4he66wkKMsOOfWWCf/QbiFPBv/kgbaAx/Z+/ye9w
QOIe5E+pYc1V1/6XTBdFvflrlAkM6jDwMS50atu6AbalHgKTP/6B8sXSQpBfQTTi/kjxIeeEEtKM
AcZEM51GAFvs9jxtkSxAWqjL3BLS2WezqPyGyHPArwJ26NZ+ta4/gyOcJUyfToksE+ds6BVFf9BN
CcDHTQ0XmG8qwAruEDmlazNpYkivr/gWF/eVd7QG3ozZ7jH/xrj0i7VAplKUWCqgZ1zPCkSEPhTg
E8j1OQWqycN0gROmfjf5njVxuurCxaaiCa5WNX3U7mGnX8VXFWuAXmfIgTo4GZ3wueNCraWbKpF2
IYa7NnZ4+X/hDG+ugUDJjUxtc8tjn75eb/s2YDuELkmSyS1qRSbTIAYT0M0WoCjpXc544drhalOT
enO7eANbmjrG3dsie5hj32eQHvT3oLgmn9AEln14sydJXi4zdco0Wq3aDNMb3GhnnmKQxV+ifJ7D
kIuuTCVuOao4n5203ZcwFtEVcCCl3drd8hcdJYtToyxwir+mNj9iqZs9WXFFEy9Kx1azanC0PVv0
XsTClBTwZlCFRzyNnjCJntPbpdxUxEASoyXQG52ObgtcQrova8qVVHLv2KzgrRdeEwKmNt6A3U1K
6fLsut3dgN3TzEqlfgtSqeGmQycYAKJiocDgJU/BhHsb06hFnG6XCdNWtPYgkjsGxTg+g+Sc38wi
7/+NPWr9dOxjrb2/L0gHEbmXtyx/ZfAnSRgYXcKFFjTYpm6FovyzvsHaomNGopFjfzAyYdJHFxJa
aGG/cmXX35lhdXQoiA6zlwboz23LJ6k4QhLYYtBuESwQpC+yvH6yxbwTuYtzrOEiD9C4egXoUnZY
C7CSLLQa57bn0LLf88B4AEMCYI5V1GvUmaJ7VZJEeo+4qikAm29lop3xY/UGEdBjjUN41LpZw3HJ
I2bb7+QU7rDaw10DE3LQ8ImhL4GXphBNIEIhDOu5mcdeB+Zp4Yblja33+Pd7dEr//UUKBv597h49
Jxj+hNKXZEuGw1b1UapSfCZzLAgznoYVfVsyQmUt02cyRmDqXDyQ7vec86GiOJ8nlCshqwZbcNP4
752fUvVIcMXqEZujHJ3sXMKjYEzeJ+HRio1n0rrK0qk5UVAhFWO9MgsgVuRvVuDz0GCBU1juTxdg
+ipcHqMpRVRZP540zEyp6egCphD0W1OH7pkeLLp8YjeLwAngHKSANH4OAzpH0os9RaJWIG/VOkhn
INyov8EKHSRYjKGVGEQQhrIxycx23/w47qcXI0mV/7qLTxOOx6BfKVqdV5D8ZxUC4mMkaXssBHmB
QQTNsK2SuBaCr/YJOunSe1xcVzaBy2ATu7yO7piqVisA3JazTEDFpN2KFMHtKYS9pLySinHijnYz
ryLdKfpCbaoWgRutC3zrfA73Y80i9yaQliZZft2vOJtLqdBMVwN7f16oSgzdrUAU7tU6eFlBkypg
djlKDXRQWfMFJ3pYsoLYyr2+c0rrf0AG0gLxrjyxBAaKrcvIPFXwoZjQq6XLuvPtEv7Fl5zNbBJM
Bp+YHKXAcZTdetsMycVhBGLB8C2nXe5GrdyEQtUMs+uRGkrRRvcJnAtaApT3Acx8DVs6o8JapzWk
fmTEf+9vBPFUkZY92nP5JMnuBZ6DAN9FgW8BbS/VBm5VMmzZboNDOp+ZcsszufJKMwLF8bxgyIyJ
PeLPexw0N7WKgCMsRSx08eW3VgARUb2VGxDJH6YzCQ9+ZgAvxRHkK5ZU3I/rjXWH4TYfipYzmxMo
daXvVOj3X2qglPg0+QtrCw8xJxjTNXk4DLs6Eq788HUFzdJ0HIulKOfmt2c+/Qh7VnRI6CNNc0BJ
LJGZevdZ/RdGOFHW/1sTT7MXZfTF5Hqf74KRSoKZq4Uqf0kfhImCwsn2Yr2e2/CeHQaiQDzCwQFI
rEetwunIwVnt2neg/Hs6Ww1+ARDXY8ItmCwLDvGHEYu+okLQ4VSwlQ5ZP4VWLmkx5kA9DMOQlToT
GJJaTviHUoT8hGuuSfuoyf3wJDNp+sAxBlrgY/Xy7UBcpPdcMFJ2aT2ClqEfEs4fPxY7KE04hsdu
JUbRwWf17E5okI7iqt4ahYpab7mK1tOmNj7QAHkwLzOku0C5J2GZ6HO24L11YWk49Qd4TBJZ6dX3
47NL4IGL+9TRaJALiHoyv8CfY3T7RxT4JNm/36PN+BNrSgBBfet2W+/dGTumEJmP+ht32w1CcJ5y
+2dOHSLPX2nvqCpHE1VHxMQjkr2Vxq2dn/uNyRPdN/Z3aUOcN0nSSKPfNWH78EHx58k7YznHscYe
mBj6hMPiFErPlh6FnDTd7Nwhwt/XiINKSn2OlavhXpepfnipmtXKdJtqsQ/akU/LOxjMkG09hhG1
WwIKt3dAG1a1Auk4vggYKKAZrL2yxVNjrxE5D+SiyJ/AQwJZDFs9heja99ja6xZQnup3ueF5MWVS
dWWZQComnRYitHg7EsVe1+oe9kIshszanr6uQMDxPuf5UTvYZP1gOId4BZ/Qm1+zRFUARl00TVhp
j1TwLNXfssqj9xjP3bUY3pnwJRNFJYeni5OWUV2XRKlCQSUQgiR8OlA0iB/801ACLOZh8VUxRjLn
s24tdlI9yVFz9rMEaX6wNbEEblHJaOLRFPCNB8GvYT8EhQig821McOisRHTJLJWETPUE+nMPThS2
vdA+uSi2KjAFvZ1AKV3x3/wBXsEQqQKqMUWroMnCL5rkosOjhpaeZva30gprOW4zH84j4mRbYGEp
p1YmBOkmWI4e+/ZvtS0+V6b8wJidSQi2GoOPe1rHPfpl3wF8pyzbVPqs8zABVj/aEq7TYgsyiTlI
AywgjUFJjNDY4RiQMbVuKHuJYDmhvagIeJM6yMS8zA3UmVW1K1QnzrjAK3q7GhIjckdQ+tAre/hr
LiqJmh8ECzhtGcdPZ1FCEwEsQlSapTnnPZf13o9wOX7wCdNFUKuCCONhjOS+cS2gYvlUw9JSHeyX
OA9r1ipAS2Vg19bBy2rVvcIFwmxt1fh7Tm1760+w/f1vCIy33qsnew2rbVntfBIeejuz9Jf0vAZm
0e/APL3bSBG0KZrhfa+9LjxiaoHxtRJc4rk1yoGBmHOI3T0EynscYaMzJTpei7BRp2/mDPma95E8
LSOsciMxr4mGAiIHJc/lVwas4woE0Ww8bqPz8Q7kEXN0VzTdJTBD7+eAhUJzO0EY2EI8jRWuRDvD
rVqYdkkxRLnw8i3g3WEpxDrhg4clzS6eWLFGdH18dfyNFqVIT+akp49hp7njlc1B6jbKWDv741Qv
409NyCAWATHvvJ6D+kajuh7djiBREiAxrelHt1aupLB1tmlO4NnVkxDZYUXsH/DTUWn5ROOeVp6x
wJ5eLgYdSbKG7bq5qiVmmqpYaqgEQhOuGLgFP+WjRKSgZdNmXoUWEbMnprlmI2j4xVl3jB5lS102
PALF8p9i5LtZSfrv+MZhLevhEtFgrilRj8F9pgTYnuByOzt9EFPBP+v7LJ/1MUcbGDDzoEOnSFCz
MtsIKS5PnKFt1KkfXeF60oFJm59yRzyWzLkYOzooicPRZMd/y7iGOBtVy84r+W2RnN/PSPFPJPWi
DUEv0t9+gIClhtGsVlg7T7k5Wqq6iAuLZMRc/EZHHUtnCGeksSsvp/xUoqGX6WI/nDGUTkXmt3da
Wp9MllEFeXBm6vfgClNN4MnL/Fu2D1zhj6vGe6cylTkQKjMcWUqQ4Gh51WJiaXwUhGWT6kkySDu0
BibLwqOsoO5VqnyCQoEispqL/VHda5WfaV+dvr+ulghzPRGmL9JyuJwzsK4NB3cuL1EkecjxWML3
cZnyyRT1WBTO0QxFJO+Fr8lGZ628d/ikQr+FXkKLa1AiqES0JKZ7TOy/25U6JNDtxxFuSX3p71/8
FLEJZKyzeFdq/OuQUXoQYFzfBKcDmWfGzjb3p0ZYdru62fb1ZoxJjX9jvI/p3ldnc2X1YmrFar04
jnmsZOZpss+vaB6x/BsFOGPK9aeyjWYd8RI7r9nc3+Sz6VDgsx2pZ9Rn0mb67nwebE5GfXXu6sRN
4TczspvwrLvV1k24jJbL2aXYzKpPwVkRvCfsZ4zHn/JxupPJKFblK8nmnA4lHtdjRtx5AwgObyOt
iJcKiJYeoVtZ4MKSbdeTNkrt+vUfw3XQK+Id402+cs7yBb3dVvFuyiJt6ivxHpQyYoQesuCxyaDk
FLpcNj0Q3OyGAC0d1SK3LlsFGibDrUTpFojQq4I67XVcTmc4Zsbs3zeKuy+mxQGhf2IgaSFgQME1
Y3oN7aGPY8z0PBaIA8YjaVe8lf9dJEx32kIWRN43pMUVqB2TypaKqxOp6cBam9HtoFS6SYZPSUGC
Yg5qgPJflgyReFGONwVdWp5ycvLcIk/MC1FeCHvo2p0Ei7InG0gPNPSs/dC97MNiK8nBfUIxcEZg
DudqGVb8XRNGgXqKHyrnSWq0bH3cRP+EorIjgs3n6aTx8gql+ZYgHbAVEEUWwznw0ahXYSRSUYni
3IsgfT2wscYX/+84A0rcfILlColaAUV40OTaxWiYdaM87+FFMOwxZ+8D2lD9ME2Dybi33/SIQf7k
X49+BTfAOZjAPc+BJcKWWgzgrR4Cs3cBKss4mILEHRH5jOPwRzxxHjbtv6QUjr7n5S2Tn2cIcNxR
bG6nvBuHcmp7FyVdBtJBaG+1eUHk5xV2koyqHsUpCEHEeumrnlWS1mG+HxM5bjcqIMbl/H9ZCrg0
6H3sWwVJHnDMjLmlMg5Pwww5VQ9khM94c/4dIEv5ghj2lqPHGiegHkgehnX4huMqvMlqDDpuBxYa
1sc0EfkZ2AGZ4x9ZKYwA/v3MDgwWuD7bxCrg/rFgAh9mzZnYXaEZ7iFhB4feFNau1vqZ6ZlrTni/
hFZfCbWyq4TuyFGvcQBMz9ntjCul7uf2v9Ew+3k4JpqyU+A3uoTe8Ld5s3wQy3tk4bVuQUczz6jp
rimfJhtjKQx6d8N14yV1LbOazvSYumxNgyZyqo/qW3NyiMjeesqnQIZB9f85BA2tK9QndzgnvgfA
SbNwcMpLaVKfGzbe/7HAj5BDM7hPJ3zE2Gvh9DjNO10bfglSqiPaLMBA9yTVwQDv1xMCAZzys8r4
EtJ1WD7wReVLaY9C1I3e+GdWcpxOf+Oyxshl6adWZh2zMfHACNxds2A9naGowPvH+hmHrNSBp0Kt
vyDH88G9vEuHR8Rj7P0iCSHtD5EgX0NAk29WZ3FXFMwY2901syUV9fMAfee8NcM0qjBTlZfPO6dH
droEdp/s3IjNIY03Qo6FtVnr2vHzTuMbZOCJcrCCP0gi41bJbf0HNBLDk1HDA4PZfuEPQC0JYwuv
2lPMYQlfnesOcVWnh4CZovw7KV1KP1Ccu6/TJ3xYh7i9D48RR/tM686X8NUbalBpahgarDR+Xhsg
pfbxNc9SISn/LQJE2so4jBX+C8rsCF2m6u2vMNUkkvk5/Wsv/HS2CS3RWswzvOibsQ0GwB7fKW9U
8ay+rksYiZdjfBZG/ywsBN6//J/qpUmCERbQI84Wu/RMcJMtng6vykkPNpRrewEwPc09OsSdByeT
KJhCLgv9Ydu97ifowdDxmy/U2KsOmV941pqIRT6An/NsirUfn3tnJX2REhfRAtqyYmXnwAOZWKn+
Yx9Vdgxvu8UAxtXVLPIcqKLAd+P+FekyTJIynWhJ43rtwFx5zlSmPUlbOYD8A/vWygmCzXJqGX/z
8+7BiIH1JQgfHmR8ylIDds1UzsQLIuLZTvptRUSkMtXShwm3ZJNQm8sz1bOWn0AwwoDw2/w6iAOu
NXdY0qIRZvJMpDPCTHCWsBzcuVpcJI02giO+MszCxj+sdryObCVFxb4XFmZXnWuvhqZ+YJif+HgE
KaRqaz4miVHrY0bixmWvO/Ulbw+ZEEQ3TKsfxYbX5MibllFGBLWmzvMQyhR+UHX2PepL0Fe6RBkf
mRplcOnDYopIiOGwq9sMZQsrJy7sClfncLTrGL2czkirq01P88FEtqyv1Ro/PXxTbbPqooiXiS5A
8tTnqYxaXTYS6WFl16/jM2ECAXT4m8d+qIbbDyJutcMyvk8RlSUPXyewvT8Fh08l2agIc0CjKfGJ
yTTeDsaRpg2i0DndHcxtTL6zBS3dPWwPYtP+CDCkcL7isDaxmtSNylKTeChBPLu6lT9Kn414HSuu
cjwATQjdQjdqvV4hPHA9icpiWWGgYhS+Wl2ShOzFt00v2NHFAuJTDsAlmn7THL0Po8djwbMyc5ay
T6aBAqKmIsTY3SHf4QfFgFEc6ViXnQXQWJtCjLB/0Pu3XgFHaO0g5NYH3M8oYto02O3eW8sXgQxZ
JstdvdZtYwoJf4xLUUxDGqHQW4hcMnq0gMY79CZG1R91aq2Ua/IUcfaO00BSMOlde5loS8NRJ7IL
buoJSYi+TZjbLgwonehLvCQWrpshaNRRLhSrRlByYX1FvtRJ68x4Qm7GXIGAw2oL0PrDL9dz8gYH
+A0+AgflvrYo88abXZFnXmrmAy2L9QKW8wHb1uYwe26UFKMBP+FZCvYrGIHoH6IK3Qsk5VSlw2IP
YFnVlw0Xv2Z+v/QWJQJDI+OocMmpptTsILa8sru5oxiY45KzIoptOsdY8wUFhZ3cO1gklkU2mQcW
SOTn5hJZ2/hpCNgOL0jjBI6ULV5hkT5KGND9GVLmOzCIgyOy1S9yDJMG19m7KUeOtohEjyf8BbJm
4O7RCezVUWb5VpjbLQf3//HELnmDo/NV4cUsddRgTDw+gGYvCo3rJPqgV0bunQMSLRPE2Qr0nbZW
X4Ke811rCzjgQKoaX1XlKvg09usyBS6Hd3/s85I25+Q2azRzuSEgKmqBR8xd6/eEg50/aaSvXOm1
p2tyRPKYbEDg69Z09VbtBKw2f2x2RVnL5RLLpq65MnkFr+QZex/H5xVHC2zBXs15tzWIxk2xMaIw
ceTrEMPn6PfZa9YXFQFDKJh4jF4KApm5+o1AzML3XVJaFwvzyT4sKBZDz9SYn6SBdB4fHl9ndGca
t1LT+MPj9EIpjRTcBApBfXKF+GBwMkCgxmiq4400NEoI5fChTz5xypdDY090p7Kzwh7wX7t5PzLK
xoLufnw6L4guR0pZcJCYuqBWJOfgtyJfMEecGsuf7B7hNsgIFu2gQUfL+vqFNcFPnV31Dw6dhYGG
lFX32ZSGzqXLieZ/MPbMijmu42AxYZaGhutJdyCk6XWtKad4QJufxgiSnCYHOiQPoQVGXglmls5T
V4uJaYJ3NISbXM4bJhP4y2HVfwZ+JTaSycE5JrIoTv/HQtwcMpCoUr6D8x/0KJZZPq3zodt8TO/w
IdRwP4nSRX0ulhB4fXDQ52oyiOeToLdO55ZNXLjBIGgfpttzIhpBfIykz9+jkvGsR1q/KV5aDTOB
1TAHQ9/nDu7NQRSL5lT0cFsDoKw6j4t5n3aGt8wtNhydtGfpSH8VC+JBgDwFNHQj/uvxHO7EqBR8
TB/U6eRBxzHkw7/r8DCHmSjemfBLlxognBh3nEb5Ki/TbB8+QU/cZ+92UrfLtdkjaxuOGD9/4T/b
uud9fAXboCjDt1F9RL7A2p7eCvwCoqTYJFktZHtFzZlVdVc1lW9G64qxPkEWE9gZthZvVyFLLFIH
MbIfm33r5Ij7A0YzSZ4An2vMT7AFHyhyYkhWDd0qxdrEG5TD5eF+8a6RVG5dd+zJ3zQO9nwAKQ5H
fAfZbSMcg0ZkAiB2Lgls6QtKD4hrTOKQShdtEMxGNaXT0sAItzTrY0Rx9bpqZ9oNHP+iHUfMR3ld
0DA9cTjHMk7sjEtzOuQ30H53sNnAhKITT3RhwdOGSuZ8rly81NZnR/Hy3Xz1hYwTcGoN/wdrf9I/
lcpXdmPw2pQbKo1ApUFQpf2vXm525g14amuvCoByKbnuhZvJ9ldDATllo3uFcZKUon/w37hxQhNn
Vf6t5lp3ajwNWh24eHlVXCUKYL44qcTPAFtdtJ4uTGqxV9086T6+/BvVH4kzkzBXan3PBxGFg0Mv
2LxgVFZMYCa/1QuH7SaYC4Opdzu/KZYCfOiYLxvYDO4UBvRxDGv+rji1S5X3mLqFUOUJLCKH6h1c
zNkws3K6fV3+q3jruzLkOwJGwZb2jzgSSS0xz6BSVpwnhqhrqORykPf9530nqqcdDtYRKLSekXFY
ted7sm5LiEMpBH6cbQe27Wd+47JnXJebsJFpUQ6G0srMLerYLUaKzRBT/CdmPCopKIjhowffjTfQ
RGBfAqBG17ZDe2dJu7DGiMhJjC/k/LZlwNrfP/1IgT6/ZdUJSPpavfAMBE8wTWf8mDHjhVR6xVs8
qpJpjrIMfvPdnhEIwuj3LuylQtP6aHuvbrqVnSGHWFzJoOd/lP3Me3wAmQUxdkGwfuXadAQC0J94
LJVRBgbILw5qFurE6rXBwd3giROKOgu1mG9XfjB3BkAldcakeRcEcp23Xz/63Cg76z/9NqKPpkya
mdLyBo+UrHd58jQJySkb+OOTv7QqYs1mlP2p5ql+2DGbWlnrxIx0SusE94NJNQU0RjN0Dq1dKEkG
8cOHFihQN/Q9pkUm11hS3GDpwC1qmQAn+yTrScKBMxqUm1u7XEPDLcaLTTibA03/MMnyPXaHftqc
/biyeHRX2YyR10pDp0E5pDEimf+s7W4w5YCIzZ34wVui0eBqqVVsyweh5qd+j+KZMfYelj1+CxGE
2OfU3J1/yIknCYM2gEwZTCti3f8O2215qaD/hGbt0WELUbVYDlrdkFBfYADVgmX4rmkJso9iKzty
VhLbZcQI7uouGG4q754CxMqGpfsVzvK1/DfJOS4B2hJUdkecO54hV750DcCyepKty6yWCTTGGSah
csK/41Uv+Z9uhUz4iuUaGYuzGgedwFsQ2roge8w8kXXiPtrO9laLWCDeGkcjA92cpIAUReKUO+A6
N9jTx2aEe1Drsc8KVH6yQQQ8uduN+0aUjF/a6CTlXBJlTgfn0uJoolJ+GuESEcTT751mkaNWQGZ7
+tdZQ6ByTmxUKKBLtF4M+dak9g2zN7R9SuOq8W6KCywLbj0NLeoMi0P8bd0KLfAoFWw2pq2QN5eN
GfNV4rri+83tWtwIloUkDM+HJ2+wqRaCZahX1OTmBir2K/HhqDhOYVnhB9jrzoo6wuEKLty5ZqDt
lRurgMCHVXt8xH/2+82GOnkIZs84Y5AiminqrJSdhkzsysKrkFOPGeeJznxQhEDNllWC0R4rFwiI
PzSxNN3vueMEfdu/vF21FZ3CaXmJ3lIZhvT3GgU31AvEHfxrWrj/1+kp5GB+pnzD0Cy0uESXn+2P
wMkHVEoyhJ9hU+DrDLKzOtTZzZKc1LhHMl+LTHLCAGpo+TZUdw45wGdEOboxEkU9gxw5zrLzqmYK
rOoH0ta9iAy9AvOCGJ0+wDXSFpX83nXYQ5trQncgFTfctMyHCLMnLG612YAe4sSmueQYVuumE7Js
eoBgK1DdCbcaFJ+Cl+7B/nzjkO18qOwSg71EBIBw9RGp3agS5X2CEC+aodXt6eOex7Cfn0DQqI+L
PFTYiE2qalui/jyuyrRMqP5PVLAjpMoDe2xE17iC/zOAjz+TFDsbT0ixusfEv4NfhBgn46/1OMP2
LBhSKd0mMUXsMJzTxZjB3bPGqD0iNcTgdB4bCzxxn7vh9TzhX4hY/FxOE5vwDOsxljqdbC5PwTKf
3junnCGIiafqVhJnl4BGBjKGOMjO+Is0eQ/HJQjd+EUwCq387N/G3qNI+1hllGurwWcPLERu3uHA
BReaGGSrYdmZfhcWByqGKc3XEGaULF38avWwa6pJLMP6rMzrPTs4HpSNH4IQRSRgRLtPI6TTZHK0
wv9muVjWN116jsy+ImUCHOf4oN/TL+T2MZh4AsfGZGvcihZBMGUjr4gaRuZOxQyXkuv5fFe448u5
m4PRKe5zkct1KI6lo7JpvBGLRepEZu3cyLsfXcmi7rH8pP3LtfVU9svwKZfbxWDzTQ6FzIDduV6x
sjld4d+uRdKLbSqTjhXFPGfTj5HILhAiCTmLDcyqgo6fcNXU0MCsXRraKv7neUFF/5EfaN8xWu5h
fPb9MvfAZhmlN5ty/psqHgc6CUD5sI/i8N1rLgMuue3D/pSSEsRCpyR/0j/tA6i9iKopd/hXxSX+
e1cISePErYV6Kdx3Uc7MCyWLutxwi8xLNIMnBBmEPJZjVuf8nfxyVAUhuuglbCQP06X3AuI64w9m
pU1b3KByNpf0X0+sw4jl4yWkZv+zUpYRGK+cGagvS/SVu80rBhvlnVNW2IVbBOqIM4UizXQ7+CAO
2o414/0KUs5rXb53iV+QyCi7WUX/OyOjma6kAs1Xd8WhT8dE6aq8w6ETfycW1r32YhzcT22CeKH6
06jWa97pC5Fz+uErrX3zOadVC96/qATrApWj4Ws2R6U31VIUmy+8pQB2fm1u5u/mMWmQ4bcGiY4W
8x4bn5VSAf+84pZmrC0PvNVMyPijxfGjJXVW9HgseK0d3nRI/6EDoOQrJn0SD2Zzh1Dhs9TZCH0V
si2ShKdLXLrEOJAShWoq4oYJYD4pw+8lXd+MoA3CxxOXdMzbuziPC9/E4xzBX5/M3TUpCGRv0ZmC
uErjeHjrYYgM++iQJH2FGGnnEgZxvqbn3pKAptCyZrrEllx5Ahtn1wE6rpopoNKAgM0XgOCtCEHD
OPuDelLYHm46JXksza2cmE7CznhH998mWFVxGG+jFP4ri7nESsIpwCf4LuVCGvPEVVdPOuSU4LBs
Gtvbom6Hq/n/YSfcWLz9uRQFf08bmPlb3KwDD91242wpbXd++yW8fRriai6FcWDuUkztpTdkuSus
NCBEsJNANPvfyqvyMAl3ut7GJjdmQkjyy1eB40PRqBYe5phHNhWLYuG8p8X3v2S8c2EnNRBINHy1
X20Jueo3NJMYJv8BhcqC9uZ6X/Eps7UjLWczoXorAypkMtR/qQCKyuCt2qIXh/pJrynrtwdJ3Cw/
IvpjEWp/viMp2xt1nZtXbNJ/zSt4PD8orWRogmq3gpY2sOqUQi+WMkeWgL0Dth1oBhFu/OAshofY
6UcemwOy/rAxlDvCwOY9c8P30kFNbsST+/Oo2L/QOr8c7zuiKP4P2Zbv0Y54lmbljPgYuaycIO9T
NJkaGSPyLQQs10n1JEluQ2i+opE9qbiAsxwQox2iBzkwvTINFTmzgA1Wspnp5DoWZQ/OgDjzaVzN
MKIR4Q10BRcpMrHedukFn0+ZiVQeZq/U5PaOYLnukTOVJUXMPWgRU9ugd8TmX4QghgV2Vbv+6HCj
cRlrg4WAYHNugVQNLg6dqJcKomLfesf/jjRFwgf9mjecOr4k4PEBdhBpjpj37I2XnTAPrSQYOPpN
IYs8Mvg1o6HwwcTvKjbbL72pqNXjyWnEiA5nqKLn64Xm+eWM1JojX9t+teoQkgHnz5/lYeVub/HI
5ONmJZTvGaCvVfT255vMXGVtwxrSeNqo21bTe48N93kiqBAms5tmh1ldb7QTX6m4jVCEPaIKjTYu
oRnlnpTrtHgMWB0WAl5xcznTiwztoEmTbgcPYJHbdGecw1GDzu66FU2CDpgYoSvkXwOUk1A8OdcR
y6OiTONeoAVKhXwvRM5lj4JGYxIZkzwo9VEwzmjq6LJD2UxvMOOHGoL1yKjoM+/UsKEn7szI4L2M
xigdKrypny2jbBPayz1zqAap0dR8x7gEesKUiWlEj598nXIRka1RlXXiQW7laNlIGbxUOHUZgtzH
L4zZHr8pNhb3ZTHRrf4y9wkVOeIahT2lsYZlbIoLILZ1m+fT4f0Lt1KB3r2QsGd1lloE+MQNVWaC
r6LtJs3St8TXL7Cpg8ayWgUC4uL/lbfhW+aovfdRrevBkTeOy5+S+K5Wj439tWBTfrBoOgaH85q8
oyxuRzo5Y5oBsCD4Eu80vSEBko/GTF4qE55SDP58ymX+XpsIGHr/gcTIHVrSlNpcQSZDPF00/gp8
ncOQ78+ZClG9FOBjc5IIwA70NFjd7pDZh6gD8+LBwbltCuUY8qVjTvPQkZ+B2RXoVi7SHRxzi7Gj
1lejxrgowj+Dof2/Kn2PyS53i29VrKQB4dfKJ9tLWkcIOZQ2IEf0Wzf5fHnSPJyo0C87n+hqmHlS
hHerdgayBWkuHBul4ss3tztL4hV7WMQXg1rMfGy8hBuJaxmCHdIy651Z3qdaKvBeyT9yuJNsreAP
eihssthosq6KjzWaa6aMvQ3BLMZ7zC1JxUd4JJ1MVmBPmHWYUr43P9ryllE8WgrRXHM4ZawW12sG
oGKkAhDxZFUN4gKw2LBBvr8wQQk7mUvwrtJhKmwWdOM1yDYHcdWkhxhHTfALtOIOjuVmXlAF4wyZ
1NUFPHW5h52Iv2yItKqjHSaUw4MB4WzTYz9//a1zoUNvgHq+JHweodNE6MJNaFdbeLghSt4lxtKw
APeW7K5NlGeuNSqLdH0MF1NHPatNNg/9bzgnl4dt0pbmVw4zuC4JVOOLI5erEYa7VljR3gaAO7m2
2NnYFtKBRXjI4QFF3EgSVKHmheWvkpeJPkws3b7jDo96rShL+Ng0CEP+l/Z0MOhepZVmA81qQgaf
2usij7UDmStU4bQBVn7RK4I6CfK3Xuhm/XkJspw9uo3QzVFFKRdLqd98G43CMiiy+rBy4WC8Z6rV
L+39bpgNM8WpbiEHUYfSg0h8lDotwJVrGxRIvEhyutTPwM9DsmW1jHRzcV/FrT6YNEbZUgld6NXJ
nqKcInj4mm857cL0VUopgX5edX2z8wo1lrt6OZDDSYb5HXsYNl1TNh3ecvof+0Tz39TjoA6m/N6Z
O6H+bZtwNHHOU650+0AYqOm+W3NptlEAMqQt8rPm/sssROQyuhiAFP2+1dOVt4jm7PaJDjRSduJ/
4IEyOm9LK3s4vewJPgaQwX2dmlpQTY1ABqUdz6UHDONYmY/mnu5Bew0NJzyBfKkyIodK5+eslkWz
BA3qldCd59Ol0xzOYFkmDacxFna6WcVlj/3Sd6YglD5IBIlNPs3mtZn96ReyUVPB9vpltyGDia8/
6qS8blxBGl4DyHMrVbHBebu9+uZjANnUnb157aI99smX8p6Jk8RmKaN+HKewkyqfkt+d9OnbRHQn
ANq0e0YwWwlnZQndybRYBne8nYpumCL6aXj7/VfVBuY5ndLXy/dr70WDHbBOxrstYh8atlHRx6dd
k1eMOoTQwvJBW+1TJN2MkiaI6s/FBImkvFdXJBhvD3K5CwuJpimsd9Z3B4DGlyFgEbV0OREYQoNn
NIKBS3jFIDmG1ucpY6koAIEEWzxZ9gd7qHBJaMlbgnlSOLdAehVHqxXTszuoYkip8olH6DAlQLe8
woLQDIwXlSeiU2HYD2+ZSqeI/O6C1KULYxW2ulKwheW1VDCG29eIDV4NbOvcPOrIVEPjee/mDxOK
qN2jD/l7XwubUO0JvyHc/7s0o5hxASLk0CH+/9HDNFdu+Fwp4hx8sHdwWpEmi8Q40ZL6yzdWxw6K
1Xc+cJuMjzo20W2zKgSPg3EBSg7VlfUATjGFl+DTVa7SjXg7kbeAsAxSSnC/tFPMFpUAT5oAOuYe
KT4KjPfnmu0RrId9uD7/dMaqa48DzEp5p8DTIfk2scW0nTCTRg+Qf0tmw7tYo7HGKlbkmnbrCQQ8
pc8GoF4gqWEXtHVlH8Dca9MnQbEu8+Vyxn+wiBJLcE/8fT4XRuV0WTLuh3FPVWB71HioBVUSA+7o
CJc3X7SqCzQKEUuv3C1Ov6DjhT+dHnlSjQrixeNX97qIl2kqt//dVjowsk20L5UZ8hzEZ8/y/X2S
zm20EXKTuqoTKABPBw1CPgw7yCgYpHLudJ/5IvKZERxpd/AcTuEY1W2UR/qPU3VkWOUC+a3UpZZJ
Ni41XbgdPBz2IuqL1Wb96nq9JWScBDprs8ZlTSmZFzrAnS+AMlG9RK8sDh1ViKzvJ+Hv3lLDKxVg
UOnMET3tCBwt75OO2RL4Ls4xYxnbnUe/q7UC+BzJ4R9m3o9WMB3Atl/4C9yEH/SfYSUyvK0DevpI
hlpBQ4umZv2TTaKmmhkVzm5kzUXCG2vHuGR/lckNJi2pn+r8el6lICkx1WJIVPC/QXZMNqro9UAe
LypZCNg90ty19Q6qb7Hz1mNifhIwip3f3G8jbV9FYllNRUuHc8FKwbe55eET6CIfYmXCy9ih1dz9
gxLKjhEFHfxdeA+3W6nbYigCLiERpwL/FrxrnPBt7qEj2K4buYzAhyBOE9tBUWHl8FH6TmwXhZOh
ykqOdDIGwgE/UzfuCnkDjmq9rK9MnyXtQcYC8rlaVZzgkhZMJG3qn/O6BFlPSPUk+I/W2re01h+6
i5SCQtYorFVTbmoQPO65YNKnFBcq8zjxjKFiOZV5Yq3x1nmKbLV7PRKrXwEqQcHecgStes7TTsyJ
Jj7nXt/Ddp0ndgSo6y9+kpxuZVlopC3K2rjbkIo0twhxYbM2+PiVlwU/ssJhf+AuxY27s4DG/j4j
YGjRCq9ZI2LLKNZhMEVkMlwshiNpmM082BbriHNqRtrb33mInu2xXgskI6mU6zTKRAxG9GnQNtoC
0QXSb0nuTyK9mAP/fKxjt1DILsA0XGeMPjFBLL6/kyvuUwBP7WDxm4YJyy+51rait3vGyIJlgyP9
o7L12TiriUtY3tIq+jWUf8z/HC3vVftuskuQg544lkyFkXT9xDj5XM4taEpOqB0LMStaasCwkRh1
EnHxducZDqeQ28SW0Jx6JMXQh+wSK+mDFa6RBXFm2qNW6bbPw2/P+U8Hiw5q0QPnNfTzp6gw5Ph3
GZI9wZk+6+t6mUl9ISJLMgJTJcRHNNQ0fCP36ZGCpV3CSx1bmu1lqKJEk1XEtxwK/qGD71pIcBu0
tE7AMmbQZ5mDc/Q05mhOFq3kBLnn+97/ZEvuf4mMOviQlTt6ZtlLX+nj1xy41Xx3p7lnRV4UtBrQ
lH7kzm66BBk2i/2ClNf4qG6yvUFpCcdfPioi8KK3tpaCqY5qGlvdNUH4WHp2rp+7SyYWGrIkYN1y
NJPy/odI6De07X/mPX0jfM0XeeUjtBPLBuP/ZBfeKvCkR7kDY3g242NxOAwprdXWJM9nCf8DyQ6s
CKvNcfdL4zvAHfUGIy4vJQZaRbTki26sBK7jmF0H699u3ms1NSYDBavLEK42vIdyINxgA6iLRl05
ACSYpATPOO8Guxwojw9Z6HIS7RfP+MpgxRgIfB1VEechEn2FD72Jz5KGtsXyw0mQd9nzWGxYQt2y
M825NEO8ksTS7yhLh4TLcI+RdsjSG/nAPJ3URwfI9TJWZ5Ed1qQbkHWCPgUoNNET5hVQf9N5+8Cm
u76XBDsliI/hFMOYD6siVlDxloJ7/rHMtsybQ7Y1rmRDJPuW7OAXJlQCPVQVQa+/5cQXVayMOuJF
vKvXsBxLC5v/luXoOb0f+JuFVcDwwBJn81O2p8LW0cv1DslCki3SPaWEcXqI5prW9BfpjgofU8HD
OMzdZ8zK8ZFoOe7n31KjNrQu3sVW2KZe/cXVQrK7go5PA8JkTkWsYCM1dO5oYISw++J/lWGpFWAp
uIRKdA2FVOH1K1VyAM51naXzSCL7320JZK6MhSff9R9x1Pt+UoyxOY5Z0tE+Q+Up0INaLP8nxgk4
Hq9fDjVpnjpXfLeweygT4rUueA7k+uQVR/1HuJqcXtZOf9aWMLAm/zO2+F/JfpayYx6R8GerdZF3
E/1XMbyMvfSKXffIRyN94UTuoVvK+qXG4ztb/PbVNKOiBfD0fWorMumLO6FCKUmNM69WlYn4iDgV
GE2g3WlLboJ/nv5Fvyg+AugLOLasx9AS+/FuJnk0By8i0tZ7TbUt/zPYi49beqIn8/vk4iwEY+Ls
ouGH++a45NlbW2x5FN1qbu0Ntd7lHaB5BNIon6GjVVa3A2e85N1ro2bI+d4BKYkjBuOnAQ1Yy+rz
cvXu39JDcCvp+7tVvbvvcmsaKK4ZD/qF83GG3RPyP/drsDbR8QTagqd+nD5AkTSiX5CyYgfojKAO
UnBEtsEAJ8zC//Gt6MdjQqmHva8f/KDbCb05VP56ApdU7fkJR/D17pOJ1xCmVFEsvJs3HnScbkZH
0h7yeGjk02FJbJ2D4atuPAYK2x/U9I4HKt2pacJyF4+CRzbzxiuGvo4mehNT4cgk7fQ4Z4DzeyM7
PAGXHy6+Sh/w5Yha1LnrgFy0NLpw48LzeIHMxYEN+FyFMY3moVlO9kLC5V5etn8dm7nyMzT1mfrj
1HhQkbXzWuV4C/7DM1on50i8EquosraEdhdjQ0nL+yw0DJ6JJY8BJmBHRSPwbSYT1Z5zoVhS0rrx
k6WFSws5Md+5b6GVHa5QIN9QPMCTRV7OTrfupGCuSm8IbQM7LR3Xw67JSg07o7PNsXByRq/7Xfsx
X/d1io+ZbCI/HBUZFvYzHUxbIQdYrD/XZcpduJYsEQY2Uj36fRHZ0l4+S+yoNTLfB32v7qHHEGHN
ktA4JcK0bDhMUyFN9iDnNOPbaoesYrkEeKrcijZKu7Qrk/HkcZl8JXaTpyzYptxepbOlf9zSoPQQ
pdBRsaolc1DERjs0vixK0wepXAFjU8JY2pF9fPwtugvFBsbXqm9FhOCZyfmylBF6iyHKnQLhPfeT
Drv+Ter7rcHd8wqfmO2hI+UPBBRGYKiKcbF6tYNtjRowhcnSXKbUNXDf1ouQb6YVVJdMDE5P98yy
p4VExwcPNtE/xdhkxFimH/9aCQqalvqnXOdeAxpgwqXUhEnyd2QRObgpK5M9dGK1BfZS8qWzkaZ2
VBaPeJrxpr2+MgS9LW8TvuxR/J5TaPj2dHCWXdqlN/imxq3mzTWYDaG6y5vUe5rckfz+ybp3A9S5
S1myQ/gr9xtxd+KeYAJlN5q/1Rc6bGDEc/B+89kA4ItcEzyvAx8WpyQEBQoRvTRMFS73IkFAC/zj
eTQvEO+Qb5+39Ti5/kQh4VG/Ol0TbkEyPO5GlozqS4PtQt3b0NIlWs+huzoqWgXLAyKWo5GaBSlZ
UQQassgd9uS4tpeEj9a8GLxVu+q3SuN1a42tA4mtVYLxC3DB4WYfdmfjn7hex00LfZR9BYZeCXoo
TQV7XBfqZQOEzN+3zM0gM3JuIUSN+nw0knvjoOWTL9K1tKE4/0Uw3p3a1e7XUDfOkkgV+Nd/OJ45
lvlA6svMoyKE3i7lAIrmpHOrUV7hW3CZrdFF/G+s+rOGpFDdwgzERENRoTsd6tt9G59yHKP/bV0Q
BcFmi+pzra5rPNzMCp7sJKB8/KVEKV1yfg15cJB57SInhjJSO/TyicHOChvGFme5+p/ifxf3I6XF
m8d6WYwcmt9njgxun1G9IUND1hZ/r/av4jKA/HJL3B1JMCPD0FZs2j+Byw21vWtVO7VEkbpzWeRK
3tZnHrF0bwaXkcC7+d1/7zebwPg7sFS1LsukGxkYLePDRb7IdhKh9XypL7pZqKWALVHN6mQbHRM0
DOtvxCzV6SmvoPGKce13QwBqABuLATPsXgzJHtHBjggKq16cHN2exnEi9uAsNvZvLOjyFee+I7Lx
tA7SrA65/Phf6bPgTXsA/QWPLJYvI153my/0DVhL8HH8alOfpCGNgjdyaVjwVePeFTsvWQyYb12x
Pfu+jLh1LhH4+rjnmH3tDJ0TLFbTI+s6+EsiDdDOjHlGrkQ8EGf2PKhJH+oH7AubBOp+SitPBWQt
XActKJRWTfwUcsiYG8C4TkOPN8SFiRCGMfkvrrJCw7BRj0fhA+4JtPZqszj0ymh02lYfJmtGOtEP
ixwVq/UE2UDwu9jUKYuK1kcsCulhm6HGBLojLPVGWwBrQx8VN1lue9haU+Y45wh2U484B92xAXXc
KT3PB1/bRnAAS7g78uVbx1JQEZDuu43yoj5MYsbt6bVwqDHGTw1GN4qiqkTAiqTd1S+37DJH/bNP
Of/SyFOVgwfrG6Efrlhd2+/ms2qgGGT74QO8r0Zm0ZQQRqeF2JZtuKF3tXRucHBeMfQQmHraXPAb
3Uf/KH6gUqRTHSnPAbM3srVNDTLQOEh3oxIQpWjrOUjAKYpt4mj7MG6rZFY7Px7LjAZl1OsFqj3t
Q4p3qgQS0MuHUWykB2m8bAFIpY4IwP0p9Ifg/U3JPeF0eiPbm1wr/YmMpIPFnuyM2ii5XGFqqcxB
ejs6ncoiPSfx2xBEpTSSEGeQzy7/vx0dhPl97G+WwuE+S35MzD6+6mmvibslX9y3gpYfNpXAJY2b
/5/jx//Eu2bqcLHl9f+OMMwQ6pFBd4Atuj2AiBU8t/NYZjKNhrotBzA0FZHECET6hYJrAz4CsPM5
UQ/t0T+RnWbdHA/e/hCMAOyJtBleOOrrINfFae9JSgPaS5XgK8E5CAifDUj2kcXQS92j9bwdyZP4
9TJs8RaP99PZnTTg1KNISO5Fa+wh4/3uXeW8mkRk/9EnZ9SgZCwk1vejDcEWkJXypLCxWB/FPehQ
hLh+H5z8ytBabmV55kzMPoXfB52Vl/BYQSZsVPR4nnzYYJTjlYybuuhDG/raKmTlemujGNZUPyad
yUjcIxojFVP7WnyylMhIjtNK09Tskkv1W6FC1tR9cojZ7uEEQhTdEWquDzKhcPES6vvM09X9T8R9
/KQxjVUBuXUU+eR0Zlz8PITufjvW2bAhBW6C5BZSPp6LuDUQMTmLWOV5yRh7DM8IdOu/ehw527dH
IaRm7w17m+sPedFArRR7v/VqJc0s7gOhZB96swLWX09GSh52D92sCjeESJ/1dI4gZlGBsSN42fPV
liRo6wNWbakgeD2OKeW9aFXy2xZWqY5JHzDxbEnYcGy6wVb8gS4FkImX1r/mO15Fdt9pVYV3Ungu
6WG3BWUwf0iSWg08Aoo2joy6Yjxx/RGUJQWRDdvdOikPPN2GIIc5fRptAJhKyM7m3rykwqRO446N
FeHhgYa25EUFTYuuYxf2y+REvz3yCtjAOxHshWOfxrtA+ConXcYu+Rwl7Sw+Ay+mgU3HJU9fqgvk
HPeJochL1XD59IBjBFgimXIuSeuAEueKtBKD9YDmLbakMDm5PJzeR5/krCY0yFa1dXKGbvSpYe8X
bXQdyitwqN+cJsf6u9JKt+l7vl1IyHL4s9+LIB9A7aUMtZfwZUgSgWUqoaLuxMXZj3JlarOxDOsD
7kWs/1k31oo2mbnQqP0ss2U+Ne/FYMzrLjN6dW+22RCNy9iSHHsxHqXEPup4b0wOvSfxYS3yUshV
jbkpa5qRTb+l2LQfPXjATlxYTz+UjEEzkTqGWVEjmDXBlc5IdrGo2NBkVJjwQM1uac0OkNKXjhxG
0xoDJiFNAX+zVeGLOXhM3MstWtms0hQ8fkzqFcXCsZkGITuBT+EC+V0aodswS0qTpjba7PV64Vl0
R/y+Sho+5mEvnzJN4+WxjxiTLFYO1UBShFaHf2k9H3XFVbQg7KCsuecsuqo5SWSaLF6ysMWuAzfb
URU7+fGeyrC7xcQxi23QWTVg/Ykoo3Od37CEjwXKtfJGqvGUNX5dk7Hg5jvVTllEqzhDfEfACwsS
nNa0W9ZRhMWvrdy3K9sAvghTR2+JBbyuUSiqsiab7rkjlPyL0ijqCel0Emxtu3aK9+rurW8jOE/a
DOR3fjWMNHbZ7aM/4ME+504o/QKyHFbIJ0qGizn5EsVR4coOkniO68INrtJhb68nDk0cCfem12IS
D6xcRgmudQqnN2B21zOj9CKsotN30dDVUXehK3rkfJz3HRdcM5GlFAzcXmlJJQvRO+y9FhTyzaZV
0pQwhwev6b+g9o2pBrdMmQ2ewgOhX+ivKkFIGK4YIGtAzPsbxMhrM329DilLZfaXLdH/uXFy6xs5
5PpjQGKLakXva80jvKXZIHHxGO2h/lD7NBbwy/HR7AWdbLH86YcKRpB7dq862mEXX8Mzxgmd3T9j
e/aVTSoX1Uu2O6hTOZOfZqw6SVrzP3j8Mn/iIjCAB7kOG3a93rGSicaulSYZ+JYXXBQDpjkQRYym
oQi3YodUJYY0CRuMFsXgY0s6lbSAg8wo8hHrCmGMHtHARJstVWBGqVbNfmBLkhHN4jtAB0Nlc5E4
+xXmElFaAx5GR9yANohV+I+XMdYcYLfhLDLmHKMd5KPMfGgBQQ1k2vCgER4kHCwE4r5bNiJsBAEQ
HySq8xwM7hoKhGyqXiYiLhVaiwGRimXrv1uwNoJznn3mBY0v1OIG9uMYW3j4ZVhiYEv4uKMMp1jo
vzgt6gK2vu6Y1hRnD4iJn/ufK/Cko3xVWd61Howwujy2bwJGQ2Hapc4XBPEOxSYhpGDwCwssJUaF
fEfhtSKZRre5yrf6/R2Oha+1yoVh2sZKtPADGKLXCIxXV43FlbJBWiXobUrJQ8FyLs7gUsABtC2t
uoGbezCOVK1IvwJMPqGXCmuNkLrkPdnZ82RdDLcKrtqldVTLEA1Zw/d9xx61KIohH8L0rg2tThib
t5eUexIFt/acK3LXjeiNwDoo8iwsWPc7BpRkaVFBIoDa+aC27AStrkvySgHLugeFT5aEl5TmkNGi
6aluyMJrqNorcRdIIFvtvR89nEVyk9XArRJPN5DODvGWqJ9pgknq3ZRDFAptPM0mHlPF43nXnoCT
1mo4UlEdm06OXu/HHyWT22c92YRasGDzRgNHcUjNQIKo4Af93fn/Kh7bw9LLJJtVvgkJYXOsvCO6
LMNPKeD6mP4jYkVllTqmCZ5jKOT4KHDSuIFnIHl+qNA7NPWveN4b6Elmofrv3Rqjm16SdhMQk77q
9/A3w0YMnAJSDFm8IKftJtYdSKJm6svSJJ0MY5K8hH2wflDL3+nKfbSBz10fED8g+Ew49BNTqYmO
INOviRn4GXYBt4FeNrgcI5u5XzvTqmjs3IyGWOn6C7fOg4v+6HA9mKOvQOWvU8McEowc76hHK2JG
EijdAZt/qQEuf7zmhkWqI3H3eXT/0NruxzU8imx+1yvHsRbmZ8WCwhjVghFnFROfh5G7ftEQBOTf
neuxZchAPf2gp8eaEJi+tXaX+utEbUMnizTjUVTiqJ7D/BXiDF+Erwx8p1T43qXJAPtCfNry9gpg
5fcEmwxbYdJDrBin5hthT+Q2LTGKElGUb2ymAgYigt+uCTP5KLWgq/LRJZ1kmbuivWS5twkdFfKs
dzoBNqgZBCTK8OV2LfEeOqDpW5JyNFtVB583p6he/PPMFper705P9vkCdp2+uZ5hzLWuj1e9rzdA
7xVcJ/0pygqT5xkgzO1cTnDcY5EzZKDnrpDoHUhJLLE8kX/uUUZsWIgo12VBpoH2U8ce/NVOjdSL
AiL+td21Suk6FOv8RM9B4U9gAdB9bhhrV639PhMTMDluJPBQheGKfxFnUJhapWAJpq18yiNjChui
EUJINTwWs2ZTQqMYxCOwAlqpGvEavmSiJmIfax7Z9OyWfvJ12v0jfLCx2eXueYpodJfzd0sxR7Rx
WLDNgKJAbf8eLMt+/jlA4zh3HCr4bDJns0MOO0dbXvLX8hQanDKS3gxMLe3gSkFL9K6xn6N3koF5
C3LbC1Gcqm0Pd24CtL1Q2VicUDmLlZDcZFnKL8SuP/pdKYrJeqLn3pZcYIXhAAcqLLZNBZcHw5AW
IRhHIMSqIUXww6ywX9FGkCkErX+vory2WHgQ0+vaOm04RBA4vPksb6kea4ptzsjJ2I7DuSIEO8rB
wKPi3o4RX3/rgaaX2wVDIJpfP4ytdbgqNT2royxfqJPRE8EAjjhDNaBqq31Pw59FkO0xStIdTTB2
stMt3e+HNLPeR1CupBEkLeush7bHrHy5of36yCkiE3ws/VAmqgS+Us6D5AaC0pmA4LRNe2bZG4Bj
ZtjBs8T+Db9t9l5fvChRpyS2aZMsbLgcajkqRpo7B4XZMVWDzUWrAuqPJ53Ysg58BvLKBaPXXQKH
of3NJvZzbLT7TToAv1jjK2+SQG3vTvWBLPWRoMC2fZ2EoA40M8uWuWe4BrGeJFBz8pscY4q7r3sM
TsYBzEz40jYo7CpbhqaiirC9qmly/kiHMF9F2tTJHLuuvEGwQTaU8EM4unkAxuAJ/BuurZCc0grD
mBS/euQ1IPxpZopZtAcuoCgiip8RO/F2sJBfzdMSNgNJAPzCi6nLEACMJ4/rwr4VSDKTveyJ7QJr
b0b5wFMuoPC1N9EbqFclgYCZ+mN9nv2hOxUjJLF0z16NgultTbIzZmBW3Gn1sge1q9mcAUR5BqqS
SvMPayiiZwwAqAdRnHJxoaXFhowd/mRgQ5mihK+Rgsjt5h2rZ0e4eBOCF5KdbAk0PSVtd4W6LFv5
FZ4Mr8MniAaROY5B4JPNufONsYDp+08rH9RHszareUNNmyKEbhhmF2tuHdFix0Pr+t3YkbSbt2D5
VDQ+MTpRggX8PuxRjUlIhyH0GxfHRO/85EsJ29HUIQcWvboaR4UcBZ4dgh6P+awJWPM8ZQtOr9O3
t6J09lFvPk89IoGGpwSFXU4wCrnrA/wCE7GHuLtrBXoDAUBYYegncdVv982gUncMaN2tKU9RJ4Xp
w8K5wv104YkaZPGIKVbZ1bNgK7fdRs/grt1k3122pAqZCGrCtYzJ1asOgLINeF+6uOum9iER4h+2
n1ybcRzF7oFW0AU68KrWFWJ0oOvKB9OhscGX7VwmBECbRFmCR92NcYHd013hvcbHKr5jkwaKqDtC
tPkDKniKSJawZtWCGlyq+OjgI/dbZKO0hfi4FswfUHZ0BhA+PhsHmRtmpKsWrTSTXOOAlwqFJ5Ph
kiNwwqxtiGZtU4jtg+SIeWAzzqrliX+Cr9rZ7D9MKMlhF3OuIIw3nHOhznjFVASbo8W0QV6RMi87
qMOxxwlUQaG9W2MRZ/by0GRjGkKHAbXXhJegEWNgBmPx2izXFCtuPNb7Bz3pduUb8AlLg23hP7gV
5dsCucFhW2uLTahPsRg+Y+5cxKnCVrxsLS15m6+XRtRO1YYMzEeSdvqbTSJdBFAeDfHIa/u0QaLS
Lk8txyw0ZuVAS8K4cK8kdm9qOf9i4COYeOvrhnpdi0nIY3L/qCU3mfPCytBlXs8ptLgfDI/xubDT
LZmKjWrnmoI+s1AV4z05EVktduyapYyVGYMnZlF+Ubk7Ymjk3evPygc2hMazyXU/bkrEh7ieh24i
jv4a/brGro7fXwLY+LCmjIy83gK1Q6839Du4z1FGIL2yeU0Ms87W7AR4zKdwBvf4j0kWwDqVSLbm
ck0apt3IINDByjCPul20QLMxs46+1TPhobtoVSdEWfjRCyhV4Cp+BQt2YkcaYtglqkCt7z/nsqoT
rgUWVGFIJSGXWFC90/x2DxUXz9sWSqJPOZFo5et+NXgPOY3xJHMBJS3zb2/H3G4CDO54jgCt7X1h
yYD04S428molGlbRkOTcWpYgofvtp2waEIIDcX1j4/14ZeBHgd2KIBRg1N4R3dPxSsIv8WdKlfmC
JhIP5Wr/wd7FnKSA6pM6nva0vkAj+QfMSI40nws0tPfll5eMTOOvBItvMLTK8agCa1Ik6yZH/ABm
0Av0rfdjzHkW3OmDaJpdg5p+uhI2qBymSB9jp99uId+i/dIhAjn1U/AJp7xCBu9j1JIsSGNWeh5V
xYKS7TIlFkTSEQ+mXlTAZhNjf5vG2zOcD1MJPKHQ2cBJbwrUdpIFoji76DGVFG9VfgebesHnANbZ
2sXv3t72w2Qt25W6l3FDJ1dViYKeRl8HDvkNhUkmV35xV7POzLhAiN/v2RZuaqoHa4sw/TFBRA7L
myAdDjJLn95gMDGRHPXX2twsJAeGex6XG4gWlrWSNzIrx93Cu5JGZg6uYE3FouOIheEkKKAPQ8dC
FTqwdYXRFuwz65Thu94Xu0e2gHu1TLy0eB94NKnINdCBiCqRzJrB5Frelq/NdrVYL6+sDlral7LP
Tde4ak3rciJ6ehY2IXUhD74lxqVprB4j+DwpY3qI/a/umE+08NEtuYUWgm1y3pQLkW1xco+I3CXC
bw7QBu3RrygC+iYD5cm9QIer412zfdihn/j0/8EUQEbjfQXklyR1g6gprinJds34UFonexjzVtVO
BSWMwo1ur08W0ry3MLd5L81+NnVlWDD7TBq0ojVrFPzcBj5IYkZXMdnOh+nSSyRUo19w7M+aU53p
A6bI6MsqQVy9ZLwwu/hinDYH2Vs9Rujn/sR0g71sW8jB+bDoAHPjkww0oeQpA0pY5F0ifXYA0XsQ
lAGv2YdELZ1yzsnCu4Uoa8bYraBEieDjcUNUTxFWvFJCHWfS61xoY0pCu8kBYwVWIgn2FvL96qYI
7jziC0kVj4YKm40UPtGrPTF5p09TAuFfA8Ebz/lo7V6EYaUuqNeosiS7zJ1860kj2q4ETqYNGEPS
y4kNcv0WncIiVXeNzAi4olAJGoK7Dh1K1RXLvB47BjsqUIAhQ0y0+78AyYAm8vcOw3Ot3EXRx96C
9S2Ez37jUYa9w/fCU6P8rvm0nqnV97sVIFwqXwlFiFNJ71HoerjXmnIMyVgFEMyOBYojpb7juPpX
IxreK391MF8oiQ19kKqFj0QGZSzwHoMnJtR8KRuWwRqnDZ2s60aF9gxI3Lc3L6bw+6qIKHFnOemf
kN+hmBkxtKCQ6eTlLJRZ9EKQR5T7Y0GCcxHi1gZ0NiP4O4nN6Z/csxmhqUIbn5e8AVIwtnjB4nDO
fx4kwCz+gh0QZsWwhMI0XDNnqVgJxJrWJDXlYk05lGm+mZSWWMegUGT1lxKH30s7wUA0Te1ycDoE
ia3CpklAqU4c76cOI8RCoezaKStMklqbYvf3no7N8yK6JmcolACz4XRZI42xojmjvDuvdDTSn0GR
j4/JYI7Qdp6vooL+Q62OZbe8C186nZJNoL2nN06Jujjm+Dpl5rX00gzEVC4C/B8qOdaftdYVcE6L
jl4giqxgmtYi8/sHuymI6Y5E9Ik5rYeC4OcGwBk3tEKg3p480Gie1Lm2BxSYDyamwScni1lwdnZT
xo037ZgK7o/98APRBZcEzO7QyehTDa6MuWxUNQMOk3iqpuWX0Su3gEqm+eSNeSBTSphOJX3Y2u0V
r0XVJAZvPtoyBEy0c9BAkq5pE6Dxc2/+oGXHMh6gbA4D0ozdYIg9eo1MqVpboorqz++2NaszCdMs
Br6NelrbHl93LVPBKOnZeey0o60ajMbTT5KsGgWKfxEiqLxp3CwnV/2xN49YyzqAyQd2/cK0oYeF
tvY2BStGM/iziRZJDdVuQOyvtuSsGToOz8vGNYbtWnuLBRFgS4kldpt0SZ+ld6plXHjGnmBWUjRi
PJMbzEa9R9pMw8fvTY7Hi3t8mlUMt9YaSJHErmHf+9nIs83DixeXBhKmIXC44Xdi8vJB8yGOa8B6
uBROT2JyFM/sM4EP90G7xQn1mBblz16WUymYqlM/C9ni8Q+DwFRlr+zKGylJMPe9Nb5LyfglB1J7
KVE//FJu7cH0YFYBHO7Tm2ouldPhjbsWWCFoBLAXI3ehn1UcOKUhe4ZM+Oc+LQkphNRMZBpcds+b
2Wd/8YTt8OT9BpMQV6Pw/Z2qO7Irfhil5qOXZy9sPSRWlZXc0tZW0hxLzT7lDdQtajty39RouEr1
cQIIqZbX7FxLzZDTMPiH4D41MEtQM2l/PLmz4kjjjztKDghsQUdaFIh1GxsCRtejxC4d71ONOcCM
tpQpCcT9oBWbnDG9x8A/ukQg4eKpuTKtn6vIoWdhSOwkx8nIvHIouTAwe7B1UTg/NmsTcJjgUZWk
v5+/lFtCFvNnmhcTyfGEcGWYP1AHGUhxSGt8kwJu8qAukNoJuXCyHhgdsUCe48rc4UeLeckPIGQT
OFCEyPcpi96g9qKzSR46af8zFS4VH8/AORcyq5CJAleuI748Xkg5F26//rDuq9Y4R4sNjEIB9z6c
BNcIXBPTE5hPP/nQ864oQksakTrq/6PE3HcAgwzJmZlV9lK06R7uy59uHY0ETSrsZNBQSRP2Oqdq
Cbnq8SrSU4QZg74o+JNzxIK+adh4FUdARUhQN21QwaiYlM800hf8RCmr6zOLga2xOg3izDYNVEyM
oCoGw5EF++31aQWLkUJsI1Qc0Q5/+y/lj0W/cJ9cOXT8g/en9MzI/9a7b7oibNAjF2TzoWuSsB5q
m9C5s5mtiOJyQ08jKzKoraY34N15pz5SjVj009uXVkn18OA77+dUVg+NakdfVHoLtULpLikVWKlt
BECTRcgfvTGs9zQr/7dWMKXOrnP2P+FHv/NKKvi4BDzI7Mw5dSPhcISChMB9S+ejjgAu9JWdvDa2
T2MVamTWBOdD9Nt0nClSwp3MI5xZQe8qqSbwWOy8N7bIEg5n3AjytwzIS9IaDyj0FBE5fmexUZ/7
84unTr1qduEOaZ+J36mzeKIbqnFBMUY/E386GSMJtaN1tuIP1/Ka8g4gXU9vh4RIZdXI3qRLWNaw
l1gkrvb5r/7lw3CtPFFPKi68fJfs+/N8HjlKPlf8sls2Y/SSFdw+ud8rsPlINTdBPbKuT8d09WsO
vl2ouc5Eq6F9fyP+HY6E/lMxS6Fij8rKr+KNks5w4cb+zEnF3OcU8ZqzOjHDF7ROw76EThqmpMoq
2zGcEPsVZY08zK3QPRgyxsZxD+pzdaeZv44uEfcvzJvG0uM9K2/aSUWn6NgbH1KQWJ1MwKX6UU0z
aQxirZ3ypul9WuOl83AG2lTylXQae4ns0MvQc0RKZB/L02llEqrbKqvArZpYpSNlpEZyJwmwS1Yg
/sVbF6UL2WRCt9ZYw7CEFwmy1AHTNoOtmDGQIU0PK8M9y3ZPCC0WjWIeRhZ36HLSmI+sWW6T+Bha
9Eg4I5QIW3egndQgbTxavvCaUvHz8wCVm2oC0l6VPcrGWuercuIVHwMlQP+3BKUIgboAHVH/wIrh
zCMeWAU/qzpD6EvNyXbUGlBIfIOoTNLV2Sr4ppMR6CDpGftdXQ8k2jqTEqLzxxEmsdI1ATN9TTB7
9JwiA6+n07KdsNHCLDKhlyycahqigjpTfzCSwobfrfeMOMjCBN1rjBysgimKatudFXZ0af9vo48r
LiVIDVx6xFggIKANSlqCw8Kawvz+b41LxzS+b+xgQTkD0P/ad7w/LytwFoGcZvYgxJzJJJNXFxGx
9dy3J2joDQT4GusyTxAKBtCJn41+JUKHdksiW/bg/b54NDRlilqxYhAWHwj3HZRtB/7tAxJF9Em+
yizBlSKJz+6KLWau7/dFOewf7AJtifuWIbVgjPOGxFQhvuwptVbqG6Kx15EEEPDOWxZ7SKiaNInt
suuLKFG5IMQQyyoYiVL+Lf6kJh2zB8ohw2kSh/xsKRPaEUSF7T5dxC7U21RNpnSwfQcGOUqM4AcF
8itXZ8WKObDjc6dH2kRv+PZK1+fALPQYF3JkC2EE1ugeSz4OFYOI8cZF9BqxlXc8YPVeckDkuXqR
Qft8r0ieDUlXhGuIs3H95u6cLJslGOw7PF4S0u37LbYXCSH/0VHC9g60YKtR2Aycv9y86DLvNzgh
UZGJWgc8mgvE0cNmmAUnRQ/dX+u2TtzXx35TISlIgbWT4yHe3YGsArQr+YQIok5koKCf4S5+aeS4
782wy3M4Q4Y+OaOUEUUWYlEhhJmG32Hy+hRtTAr4ICnuGibHAVSjBP9ag/GQMz2RW0j9D2zgs04V
+sVxU6JWQ8uoZXDDdtVA3r/LMO8V8RPZbipixQmPvjFEWM2yI+CDWVgFQlDFMb9sJ33WfRvPWh5H
Ds5QgXcz1oNIQqfrq1nj1cX/h3xgs24O8dAZ/AxBnfywjtPcIXTwEzF/y9dwNNERj5jIAG094Cny
JRkNUw49TPeuIrMHx77Msjj1mrd5+4OzBQXh1zoX48hDr45yHsddQop3svpoJrRWL2kLAomJyEaM
ByeAGnMpM2OLQHDZoNJM00Zw5ZdOjEuLyCN9UKH0c5g71AHU+pi0jOquMSvxBAZ+nGgkX/Yfz+4c
nWzMiBvckHDTAi1tbDgLnL06/XOYxZT1bgkvWTlwIDKXeoQ/1pgzVqnAfwxzsdphMK0rs+4WeoL+
LyJxYRUcYFVDDPr6LWQL8qf6/hwlECk76dfu3V7lL2dLVYUjeLzLszHx+KAqjYzW1BK2kQ1aXZYH
n3kOmxM803xfVW4uzvccyzbkBChKCAtO6Z8VmNGTou1YhMdGYp0lGw8/UKBBTwyBUZZKEwtX/rJ5
A8iLsSXMWb1irmzdwFXuqq+qe00Z8vW2bJvQhtN1o8pmIFNi9P2P/1Xy2WYUdEQtDtRR7yXyRt3P
QWkLaUQv6ej9HqFU86LJ+sTV2oqKfK8fW6vdKDbHywS8rS2AyShgPrscTTWFOutRuMkIC1LUySij
n8U5h3tbs+WDLLrypPPm5BowtmPgixj7+e1ih3RDTNUZPGX537wBBw6XTQVLyTLJUqBD8KOYLfIt
Aizz6j+pm+jZ1C5RjT4ju+5CsMZUdAa/U7XxKkQ01O4OEqNtrwXLBqdShdvHVmF55GWNcFcmeRZw
WqJ4e0w7ym4OmOb7GQfBnFubek5/MfkTvSQ8dAfqzjd1ZXGUeNFvST+srUIaOACWIBwMdXEQLHHf
oTgKOisgvjAvSMQ50J7/OUVG38AKEfBgD8QudOywZZyC8h/v3Z3dDs6lCwPRFurm+icx9ydJrUta
blWwsNG1P1i19RtFfKlGGCnk+RFCTLmpIE8FBNx+vTTDjLjcnX6q0mfVP8yALJpyxNWBZ3C3cKDN
sbIObLc5YTkCTPdb1RTnLTzBFN1yXUb+Q4CHYJH/4rPBJLF+SpUcG2jWlL17fPSXX+hbyKAU+vgE
UF3TrTVlcxv+CPUZDrTUZA1R75AUeKSRQJpUOxrCH/nxp9k4aWjDW9ceWykyGNsGbPkjE8gX64eg
8GZLRNDN2Xp/dhPHJVoJpymJNtm8AsBZGIAOIp0BLdaxorXP1vGtB+nKZUe/brGQURmbdsy3BdkO
6P49IBb1NhIpWBNbUIT4iFyuVvmIz4kGkB2jDFUY89lTqNBwDtH2AW/Hd2Lzw/1yQN+qJnXku3CW
7dbkB2BBy1falD/mri0KyOPN8GfZXTkh7MJ57zX8F4HyngXtY+cuiNjDFmVNXOgcPoRdxXE3VAGT
tAlraG0cvPjzpB5orCM3NdD2jQEJdKhg54B+hxWodjZtd9AzA6vKmRU3lEuoODhM43leOqJsChhk
zIG/vzM4bFEJQMVUAanpxB/kBuqRTU0Cm588tZ24LTbpqctU6mE6CN+G1zP+37AJwCu9uc+GV7+C
L35BUarE7xXixZgtufnqliuF7BhceJJg0NiGeGGpB1F3GHvvoZqRmURr+/x7iH4ljs2ZBmkiCwzS
/WfijfZRNh1GUDcWlKxa7DkPXMK4F/dutmfmfJlFbP66h5/3PoPdYgBd4B1QiM5c7p46IJ9rcffA
YsiSUPRMXQlRm2iJ4zE8NCItU0l5ZRfgfvkDpZW8q/gMXux0ulHRksIrcOFemvek+s8hPdfK5QGx
FF51rvxxQjPzOmiyEot4r9P6eLk+b3r5qhugJAAeQoEZVFZPm6oGTHSb6+sn2AL3zl7b+YnvwJN4
jsYWUxkEaR5tXeH5rdkQhkM0z0AVqAEJyEOZkg6DbTElycUfawHk0OemFVWZt0zSn+sPAi8f2O5N
lxjNhhWEVauutlfzxSzuHsgCrtRzt5NL/E7L24+KVN957AA8knAYZn2dp/nkF/JY7qZDDaoUHUHl
pPNuI0OkZGfRCYK6gJBcWVl+YDZ85yzHK+HYpaPFNuCBuaKyaPUEuQM4dx/JnkOW7gdkpMNJbRyh
1g7W054qqkPyNC4tGVLpNKPWtdMzL3c0m85IcJq5Y4y74cyl5aOsH1vH7HR7fiNxreWYdjFKrKAw
JgF7XJWkBFQuJQDwKFRsr1tcCOaoexTJJAw+JrBHxzJCW8X8P9h9YsFGCMRlFSaGqWHLjg1aWPNI
4UGxZbA9se7fLWpFK2KwhqohGMnEjqyCwOvF1tp86KQ4BQdPBSmnCX26nxU0w9Y5HX2xaQywOF81
CCU+Lpn5nz+Lj0YxoOW1cvFl68TFjISH7BN2Q/O7GfMM92+Rm7ZHBrQfl/tm7GoJStECsronNjUz
uUBmpqiFbn7HTjwD+4uvZYBsUDmZQD28fdlfA7aKU2vD52dSSgsKURxmxh0Zn9kO/hdcIY7CQTFC
dzne7bI7IeMv8jPR+dz512+t+BZ5ZpHz1YXd8KsCzRtDuzxz3yOu5JLzsbuuC8wk7hLKqljaWRoW
CzOWr90QaVtHrJcZgt/jhx5jekZDeUSW6lpyU9HKJRxn7oucXbpkqqLkNgaWEeRRlNvk4KtH8kNp
4IylxTfr450lePVae9eEAPdNdw93UkEZghgsakU8/QpDThqyDnH9bnU4f6lrxlDtob2b1OaXg5Qa
bEWXmj1zufAsvrJLu/mwol7PArPuYfgkk1d3YF7el1gqn1KmFsLRopdjACZnQp6zC4QyGVjy6nxf
GxwKKqRct4YE2bY5FYTYAowxDhqPUN6XSVboLe2YMNAG2vbhaI3vBm5JkDQrP9YnufPLcDBgD1y7
tYMEB3bCDmhZ3ddqFx57eaOV3WkCCiyy5A0jRxeNi3P0nyjbo+XWv/VqJLjppR3XJCdMab+48iWF
fdKCCC47KoXPc3E+Sfg5wsg0skCP65esR3sBXG5kJet5hedGZiuhhpTB3c11enoCVkZcmuF2VJFX
2eC1iCvsaY5s+xHuDwL3Bti14gfjYwZTGY/1hK1uCd8gm8V63ElwEkQtcyw68az0jqeBdq9LbGr0
jg4CKb38ZM880vl0vqJ+jBPAZDVIa7uWRHRbLaziHbde8/H1XEm4DuVLvYmy4UNAe0+L9Jui435K
T1EpvZIr5ImDFzWlkfC2/qwHOsqsQ+Y+qYx4mfwA/rhFIhT+CzoLLI+C8WQpcyDbq/tU+Ps/Y6vf
lJr1d2CCtyM53zblk1Ga6H64rbysfgaqXCIbcg2GP35wvJ2KbLN7OoREJdnJbVppf+/qOwGl1Oe0
/nKiNUX/crq3kVZH2V6PhonPr3nsM3bj3G34XtVtZFc4iNZU9EZ+lUTkH6KAIe1IwnVnMxPAzExx
sjj8Qnyn+6QDPsLEh6krZ7IWy+c0FIVFf59NnXFNL+6jC29lg0ZfCH/bYhQN+7aqzmlu8he8NB9M
TYBnIcpt2m4uF+owNqhD9ZPn8orO0RY2nATX52qJayH86SoPJfbNiPcBC08n7dx/GGVs01Qd52zj
NPPN2i7cDuFlVSCKHt10vIIH2BGuwYZ+0UACcWKT3mTUsW6sI1Vf5AXiOTk9UJDo06DJ+wJHRu+Z
43GjEFH9o+9kCwLFa/8RnWNq98fjDYPpOjZ3foO9iZH1L7pz8qzkvAjmQS7BBGR6L9Km7r6/b8xY
6tDz1aeGlpyiY0+eg0zS1orA4dKPTpBIdVBmJfh1weSkAT5ACeuQqcyOPIVxV/g7+vdcbX7Mh4p/
38XzdVKFLiPSjrlyz6iPhp+1MsuGB1VCzefAq5tm/Sh98qNBgyfjxFsZ4oVCF6YIS1ZAbk93Fs8t
E//Ku3vhAUTGs8atLe3fsPVBOifJq9XF6V1CfwGlfE6YxR64uwusmfzlS+SSsSZIm+oTNsMuUzIC
j/zBfV85v1NAp2ZvI8f+EDqOn/xYswyzZCva4yMkWOoZbE6cjjh6CS2WmYRsPcQbH6Fp9ksPLf16
p7dmU+BbHa2amMkMyBuLjt4sTmCCPG9RIJP5jnv5MytjL/ntV+k8+7PxkHQz/kTrRjWC6wPJCZ6V
L8MZjxdotRcKDnBVpRbL2SxT7rCru0X14Xd4UMh12E/sNGSk13MZJMMP5Ae6LhZ8eJN5/1MNKMP/
hYqZ3CYWaXjxQao4Tm5mPxc5qbWdvShY9TJJKVehdCOJKwLqnIY9eZGe6rfeIhRcGItb0CbXf9/e
WvfywWxHtkdYFXVujJlWV9n9lMHQKys7L1oonqoTGdCksMSGlicr2neNQQMg+iB9kO/xZtyzW3QU
DaK1Gs5akdZKonlK6AuNTHTRBBNRV25TZvYWX2XcVpmQ50BDndp+G7DQjvW4UcWNRzkFMSvqAzKW
YtRUyhhqfeQtc+9TBn9mV37C4q8eFxru+gCAtL7+ZEsbrI2SwGnzAw9sX67ebhFh5ju/YUK9PsjL
k5cpWzOMmFig8DAJBXEgUmK4A/U4OSJ958EXpcUav5wodZWk6x8jntLartoLvey2LD7mkS8Ru/TD
4pRG/cnpeRvwpEG/L3PLnVEbgFGecOOpXMFF39e1z3rfJ+RCCBvh/r+VMutr9KNpMdTF5BYNvaOE
Ps2kMh1IXZs7o8xatQSRZ0N9O3uCW5DoqoMaQSzZF9w76NwCl8OcS29Uu7tu7QJIsB+19Ke7IKSt
2QGOc5/GMUV94uNaMSibBqRRJEr8nbcwPIxLnFY/Z6NWaU4ewcypBr3K7p+Zmq9UhGbcvSsBBc28
HoRL30PzWNisPotQnmUpwsQv2IDeCgp5fa8/g070A7SOYM/pynyVlKkaa8o7oEOR3WFJY5n3tqry
3SfR1EpK/aRLukHcaBk/sVjX8QO6g0g+XevJ5VxDiaaf/kvqItlraL9KSGZaRjf969qIQa3CbBzP
yJyN71g98cvV7A76m1pwDvqaE7xHR0R1KgAx1YATwbv+CH39hpfCrb6H80wJJSI3jyIQqd2Ti8cm
OHAGxxJwfdACCU0FArgBHApk10el5hNMnX8iBbJIBT8aCcjhoW5UoRI8ZBwIryK3fJ0gcqaYH/m3
JE95wkRbfPwszpwnPyHYXWYohWp+jDRuHSM9wfZzrFf4GiqVBGUYf2qYavmEcYp5g0JRyQhQawgg
ieUNzhfSWpPwPs8WFyDyuaOuTlKM+s8GdSeDAmomUQt48vFpKC5BGczcPYJvQMEpVJSdqZYiEj/9
afR2ZV3Qqvr2hvlcEd0fVC3V0Re48lKxXYj3+XqRZeqMnyvuo+hIQwqm6nXh7r4epTFqIKKprmHw
Bp6/gxF9RVjxM1/07X+etNBeOvPLWMLaIXXXX8NN5f6/gBZ0i/ynSM31nkU7/x9b+5zqpEtNShNh
ytX2XO0GLtaGQvzq4sD3P0/d8lD6cUNS5Zb3x886tM2lQZTqzYiIWmA2FPot6+HL86MoPoyeIvHd
fwcB4QwHRrn+DsmBssFKEw8d2mQUu5Wkh6YZCqIMXAGA1lPfMLyfxPYFSGHjRPX+s17kI3sFY4vN
ej86G9hUiMKC8GgMGZM+pEY6VxibSld4944KQW48fCIG70bdWCF7KuxuTaI23fFO5tqcS8EkxYSj
0/KqLpgedXIyBUKAYoCiMkncdxrA63sYcJXcDANX4xZ3mSpvFHD7ZaEVj8nparKgknQneb3U8qJi
RzWR6rZgtwjJNqxRxtL1sTU+Uzsj5oqCokd2UNSYSTgpRI14DMs75ockpNyp+r2IW9MJw9zXxZjD
V6fvmXKKcOdCpJCXhB/LU5G1hinJm3F8q4Y/iw5MfwUzoA9aJnRz/+LB04wYQY1BRE15kmxde868
WV167U9Ex+wVEZpdmaazH7NUh4z3ntTOv3UIx8R6+Vxki/V9fheyw50IShiBMGZpL6Jz8R0ehP01
TfPmGrJzsi0vLip5r/k8LEm1/PXUPv5RRIW41XXLhmxwiRJerzGxz4u9R+IEZ6z3qGmlvkua4NLr
kpb6MN0/jWI5sut3FytAhOalCRS5RISS5VRfSF0/IwEOaEm8xUQJY8Q93Yp4lLKEaOs1VjN0ImAZ
CHgZJsdoaVqSEN0m0F6lfbXTlEf4SfwxjYFKFSNaxw3AtXLpOBiLJj8BE19C8SpMcr9XanrByNzF
rMUvMSNef9uoyYQI90MQ7b2EPtexIXOwN7LqbfUVJ4tDdCIaX0kNP0bHkcxXIashBHoCHxCI9hjj
hLEf1OzxHb+DwsB9hMz8/igCw3pHJlrpwxtIBX+EM2ljgzzELAdypGg7SVFFT7ytzSrJ05rpoTlh
Ns7TmAz9J03F3vQ73iT3S1XMvMX3l3S2OzHMPFxz2ATvw2D7s5YFLUnOyDrHtTn2c96dgkvTELLv
iaiN9j6Wullq8Zpkse7eTbKOPFXsuva404oZn4epQz2qAsqUcVet2NPbnR00Nz4yLbPJoaUa5dHZ
WiAbeufOdpIWTojmzHvhH5Gg4k4dFEecVvRIiDqmmHgIVRT/VNKXSCEqrIqHqGxom+M42c0qBnKP
1lJP/KMdfj6hucomHTyukcSmSqLIiLQMsYvIDwpFI2E+dk0UmlDnm3p8R1gjNEi2VmVWpUXqT+wH
Ql/IujMxDdZsJ0XOkmcHojkjpTRsZt1N9uECHeioKHA5s+hA573MjXKNTs2dPov2qBllGcZm0evf
V3+c0QOWzCG/wFT1FHEZqtO5K35VHVXd5vduefJ/GVSC/coJjtS8RqZFp1+tGPU+/frfmJCWnCXE
pmu3hNAHPK8tNv6Wdopd1oHw3r4D8Bj01wECYY/Dbmqwiw+q8Y3w+tHLDBGt3AEPedriEBkQ0hv/
mnH7XMP8TEYXlr6i1J6SUES3xhqkqyq+YqE7KN2/krC/1xRwvkZMWaIFyjbHB/Y1U0Ujqp+g5dzy
9ZpvEaf/5bjbxD5bf7gnRuK3jc6caI2N/y4hlK6Mn+aq8sxt+re1XKDYMki4bpSj81siWc7Zjy1T
O3H5X/d/o3dscmio5VkSEV0lyNukzxo5ERHJr3rZphvnI8vHA/P11TuFlW3XR/KI4EM0s5KLE3hp
EBpcW7MeI7DIKLMLBPv9k6vsynque0sq8+9Z4kZo7smY3s2qMw0Aba9wxNZPY/XnOjz+ERVfeDrD
NiQaZPDaqZ0pA25vuELPaGHQD7FlTMukxL9wvfikbrIbGwXEKCy4YmbBe8Re2CPh8T59/ozdN67N
BWHcxCpVMMtPSMxaExEI8B6Zv7HJdSUPrGlBbzbuWRwt9n4i4ie/Fb38ExYcbzFszTIC4TDYNnDw
d5rYWcpsdKRi6xJTq9TUSE+eqCIK8g94f2+vykR/KXyCnF5fowPrwneJanQNqjgCyjbCRiM7tuep
E26kge9aUoD16fgMZLoc1a/FEbcR1u7LXwZrSLRf/HfD1ppPjRH4oIsw8BDq2HPlW9i3UdSlJ9P4
m0k44XkV9Lc0IjeDsnexNYLKKGT47FnDFDwrIvhH8fTtyr0STTw3z3b5p1s20scUIz/I/Wb1mdVs
kXBhUuEkhyCvIMBgCszCNPc6WMBlEIRF0XfYe9VdMxudwR20IngN7tAZvgAL3JFJ4qbghtgXVyGY
3MK4bvAhXrLu0iMxGcJjbfTCfJqxh8Gj8EsHbCPRBjBXBUhETaKXgUgR8IgDFMZNl52XyXUd5WEa
hMXe8KyBWNzbGYHk7KvHty1fRYS74osC1Po3OG+uE/uqTjaRAmGoADsVIlFfTxFcEfVMHTPf6rcy
Jw66hOETzI+bSb6+pRtnT6ZajvbIGp9Jb7B/He9CduGBZEy2/SdoN4NfXrl4ssV0Y/4Ell2yBWov
5mJDllvolsGqHaU78am5r25RNmdCbtrI6/kSfuE0IUwZHMUFS3v+uIUD8tVsv8ADnlqaFqEwx9Cb
G57g5i9q46MmMRDW2/bvh0+Mhc2eB7sQS8S/yZU+hEG2Wwc8Ac8pgoUEm6JpXLR+u67V14fErGdg
H+RTIuq5i6B+wuqIThqJG6MxLfkkt99ZdwzDY9KbOMxcAxjw79UMuodd2Xw6tLUPUbe1TzVItyTW
R6sYtDhQg3kWvDBYrZiCNrx9h9ZXqE6ywYnGwUOzE+5y1nZf2N/9KkPKiuWCTef1r0BmIGCNtZgb
onlAD0dMKQnUOS/E1pZGi5eIf3IukEFnALUMNJD9Hc8yFfapbFouqXYVdBBxW5rcKns9ExxyQJoE
DvEIGyfqkLBGugceA63xbbwzNHPyHw0MwCi7RGtWeRtu45ap5rMXUpCKuKmC+mPpL6UxA/xsUo0U
MALFFGM7SfIQs43H9p2dDfsC670FWeFZDKIHBvO3tLQ/YDq6o6z9WEIYx2SspZR8S3XnF9nzrqDv
V6dmey7p9unShSd5FMgqyBVZDhMadt3y4XKAzKoNcNJQBjUXz9XuDHtnjayLrYQkswMNWpbkXy/N
mlCZ/exiTXkhOKk5kX9SnhXH4EEkvntOgiNGyzGVON3sxha+3Bwe5JOfGncRhAyBZVtKIv8zbHOP
6Hsh1Gl7WSD2ZhD3Sh/v3mfwTDT4dI10fcygsb4Y9zvGHEIvLi0KqXAso7gK2QKGKXmg4Xnla4vb
oz2Nu4bRX80mMnQw0lKROIkxaWJHXLRmsA9zSPETL47yw1ffQ34VTCo+3PdrP5OLhQmS3OLMMKTX
S+UsU9wFetjwgw+kehpe1oBiimf+VZxS5aQagQbGVYu6tLV3eNZo8t2ZnNxeCaRkmNsROV6I+4ZT
AiBuEDcZwjmpESIfn3ycIhGwIQ9VUarOK7UoSEvBIld8xcJ1bjz75ctRCi9mQnrAoCs56r11S7eY
17Wmi75+Ak/eivbiofknQejL5skxYa2MAgAY3gQRjtTqQEH3PNyXRYWP8GeBExc+5ezGDhBMi9E6
IU9w7NF8+KfSNhDqWxz/U3+BnABABJmmYG/c/R0lBHkhGD353ojNecJK6iFtfPQGeEbovFJrnVuj
kNZaidT3UoMjD3VfDZ3YtEibrDTcpQJPZlKWY2i7ifwip0qsOEIXCKpOMkxqBHRGfPkkA6fNyAi+
KMpgWdbs0d3RxjK7WChTFLVKf0NjBOXRnFtInExYlc5ml3qLDZN7BN42BD1Vhv0c9+rAIRnK9vvK
DBZFbKKCCBVmuFuSBsyQC3Ru7I/4SokFyxGqBoqinoNiiX06tzfZntUstkgPMhUC9Fv1aVuIlxW/
f2f67TNwGqd6JZb8qUGeYZ7oDScIGjx82ZlX4O8ghwfs/lUPTqOsR2M2qicYVvUJAQM+XeiMS+Es
QwYhP+XamhE+bcVdzbC66oU3nqBxStbNZvMd7D4h8duZWBJ7v96duo+CCuyFxnJilbI0xYUHZY7Y
ISPuf/tTy1dPI39PEaUBLOPTHwIlctvsRr1w8NwRYBxuQHm84nZNvOoWu5Om4YWo0TLjrE/s593M
Pq4MqwMkuX//cT8C+09W10yGc6Y4ARZ6QYuJnvgxbRSv8LwFIy/3dhEd8Z7xglRlDpnQed4DjzGV
DX3cqzfI5XDpQowRAITz57jq5oO5/ThEgs6hCdKQERjemfhnBDgsRTqhm9AFGhuRsYzmB4py1Mkq
NteKliry2hKIhxQ0pBawpVqfzSPJdi5w8IYixUkTHr7v7uCb9kf08Y/2lA5zB54c5gGyvDQ7oUUz
/bjMe8gREFhD2UI6vLj1kokAs+/8X553tgaZbwk+6XvqFcNW9CgLGaciv+DGD4Td57juFt+HQuGC
SI/4OJoYbmwJwfuqBV09NYTzt/Dnh+ppbZWZ+puinR9sFYBe3rPNvm1izO3KYxmjyrz5seg0Q501
x+hauJD45XsR7z2yuJRUZ2vcIc5rjH757pXtSFvWFm53d6ptvZicFE+9CgUVWshEnBVgMy3NvMcq
j9iWEycKhtzG5rbNJNSck/ZtGbboCEuKb96T50Usytf6EV0KlsnoLY4YNODReHqTW3Mjl2Qo2sXx
t6zvacrrsPi8AaFeBT4SGrqRzEXCMfnBIqDfdNJuUJ9nbCmKRKitqwXVWGiF2Xqur9lTNHmNRXNE
6mSlyiQ4jiPctRtuXYqQ5lbqlrjJiLXPVKfLP0B3mpM84Qlb0ukhI8PXwjAAfq2oKOJ6lP51OVQ9
XunykiFS1G7Pg0II4Xswjl0fJhTeG65gG9sknJzjcQaR2fuFJTfNypCXQweH+3CDwqeC9hnhVfVl
u8lpAx62i3i7VdE/hLSChfANwEtZhmFMHf+2e9kBgkdmlmyPz/5kDoSGEUGkbhnhkwdPBWcWbFJB
ZqqPJtkvFD/uUS2amVwM4reaAGApoTkTfDw4/wSJ1LakDwv0gSVZQdore8LPZYuA2rTfs57v9YHM
6Hig0nNsSYTPqNnTeRUqNuOkv0gZf4zvqlZqp5mDP1h0F7MDa6S4WI/wQzrK+/XI5n5nbZ8U/XQG
gxGKeuE8HbP1KXyfsACsrh0aKyuukHtR6Qitd51+to03lFZZ3Efg82Th5xgOtJJ4laoS5hnQ5gqq
H6s9lnX+lZcBtBpVGTlEUF3uYRXa1/KmF2erWdx3WeqaXDulJrFVTMNEB8KR8ynWqoLLFBeqjYLm
wYBy2dZH9J60TuVfayeXXx5tTYwTEHupqMGDcDfTFPc3mITsDlxIMqEB4MX4IHe4gM2yHkF4DOtu
BXaSPFpiqSlRMDz2a9KonQ1Yo8vuxUwDJK3/vhExV5qNP/f8DT03fln1lU6nOUkou9NwJkD80rxo
MFa3uQLBEdZAPgo3REkuOFhfU8kpKPBENnjs/LIpho6LiM50AWPH7lroSJPwOSjzCimZISR3Jjd3
qCqOcDCSD3SOVNtD8iZtmjosTyZAKB19l7ps0HUZxLCzfW/BvGZCb7Qq6MmxB32wubitGPgwUg5p
UfKivpr8gyXHbzhVrCrovy5sGFkMBIgovqsUqJMS2z63n+TzNWo0gS2YgOP+JF8NWLFdj04tS2Xg
FK67pDH7HV75ZmLzR0f0qMlmcmcDYfk2JofRjwfRem7/neYHnL7Q/AKMM9BTO005yWvravWFmyd0
9pByXBA5AqJYZOBvcVK6Xo3kWZYrHKoNnNB5iCk2U5Xs6752MNPVaWbHji0hVKcuLdfA0r+2WN4a
wyGApIfPOCjRuKf3rou0/ptFZA6Ou1V+7jV4Ly2TVotgP5cOZ1jl4yZYyGDBL7bhX5BtvPh75ZEF
ba6hFNVDecV80SzWobLXyzbi5MPlzIVAV8+jPT4BzeXB4x/j0q4+fjSZ2pCf7oyX689jPa2S/Ggl
2R0d1TnQueSgmKeQFIvpPVpfxSbAYs5W6gYF7xlpXsh9TW7yyqIR0ykLtziV9eIxR78VqraYLYOk
OaysGh7KjsKWXmkphkOccJIfhtXTi5+ROGm2KjwyQ73WTd+ot/mOG52lmP7YmJL64jpm9doJkq3G
E1Inh/8Lt2v/A9taVKO9+0QI7hgQgDJd6xLM/npQwYN1AwgZQKr1IH4zg7IMERCkOIYaSdc6315M
CWXsaLg22QBScSJgmbv82TwBNpiqT4czu+Ezf5aoickpa2pNprVGQhTf3x7bu/ACCFAIJu7pOegF
1oKqb0vlujGqiFGT/5mPS9R3+OXCFJCnrgbDVbq3myfVNbG8PeFqSxU0iYzmN0QMuhFN6K0/wLB8
bQQ9yPdbHYlozW5U8iPRpQ2JpU4U5jC3kPOCBDykhSeB2diCAXGyiJK7m9zBSLCidqci7IrjskeU
lyzZ//iAr9YlCcqeF/AVjm1ZdCP2EANEP2+q4JQWEYMsMQIorH/Oz9KmIBSGtASg9cxEilsFi11e
AxjUuonM3YqxUJp+X5xGeUDsYNrvPtUo31JnLJQeoHLrh+2ihNpPEeMpLhUxtq3RETS+l6Rc66++
rbge0hodtgNG1w+kduKx5T0PC6QadXHOduHfjr0F2yO/y7Yqk+7wXFM0YqirNmim4x9vWaFixGcl
Ldx0wX7PACgOH5p7zVVdk2JqMNejbnRjk7fZb0BS27s1ZPHj8vEKdsXx7hfCkvGKmPLGy3cnCdhU
Gqd1McOmabyaN2IPbpWDTO0Ep7a5ubudUeZdwyb7iGYQr1qqxrns8q6Glqpqe8LO15Uqd+Q6xVpq
8F0y0zRQAYRNzLU0zIdeWjlUmueTZtDGCwUax7jbDWG8Fq3Zdq6MxQqJqBlSFfRS2SG2zQMMsfYN
j7vucaIMU7xPpozXTkUijQ6uRxnRXTl860kCBJ/Xz2AYJbKWgTpjp7fxJ6/4gL81aFUqExG3yDLi
HeL0rRXvwAZvbOnncnSp3YBbMAYYpDtZjAaoUtfrrC/ZdLBG3Vck7TSx6URZ6BrpXJkFHaqQ1ZAD
8zDi1UZNmHyZNwCh8HjvEW9GPNHwnD4NE4+RSYUGoKcKdEPmbfOayxo51fTpvKuJOp/SyQi0gfhT
wqwj7RwnsumbZicZSxCN98nbIvIpZgZHGzPlEqaq0VzD+DUKAevt4cyRZRngGDDqqZR2kFyls10v
Z937n9F+abdfxWkrypnZm0hyIlAiUjvDogZ6pBF3XTWpYWYwOpmaeXFWEvXP3squq6poQ7bX0YGv
NvF3+g3Yswig5imy6vIF/OkpHd0uAyTl8smaAOCKZ+gECJC8LbGBjruD1WWsI4zhq57eNtRokJ1b
2u9OeglDarAft8nAqdfbjHod0n3dBNAtdlnPTyUTsInPZZmFVbVe0DPIY3RWWSkP4pDnA4z+7BpY
rkEcpyuLaM+t9vw4N5XIRd+A3kPmOH4AA7EvQ0JCUaNA3pKUDtznJ1dpPkbhneIUv1KCUtZzfHap
viP02ACG0KFeUANHukfP8y63TQihD6xxM1wArK+ez4jUaUzrkvGRiXjQcizkN/emRgCTmSzJyOM1
5N+lGr0OgY6QvzwfYRi+HEHPAhyQvI8vNKxVUMzgpvRUm8Mpd5UxrS0UbZSiJCLdfG5RUr5g65wU
LGkbe80OwlkRaRyl3HejJPTaFIxLjlawnptrBC7fCioFM2dZ2Z4GgJRw1GJDeMYaT+9qet0INtof
63sHwywvXVlwuiBX0OEWjwB2VLXW4ugfTUf+IN6Tc7R2pSmW+PXbL6fjZZUA+hRcDzDQBvM2hAUH
9XuqnEoz9uXgkll4D7N82RLdJp9K9dmA77X20NKXxiYXaltWjz/1PKNAMd0XwLFj/QHMjJWxNSXu
HmgwKmRV7QkzCyeVnqpk/bdEen5smGQowzy2xy8KvOWx6wRrNsUpx+tFKxKVH3HIY0mZOwaH0tlq
j73MjAPqnoay5M6I4hA+yeKA8V0IqBvFlWr08Olvkyv+xc6Bo5cR4Wr0D/FJF6cgl58a0tM1R5X3
p34dFbc66dtXJe/1xvBBbNI+TZT6Wso4bnMjhZN/lwP4uk7LKAsFD8mIcP2s9guMu4jzJjsMiKJi
3TL5TV27KFC7NjJBAFGjVOwIH9uKFu4ucPmifFofqGK9P525Gwjv2s9MjK6JFwUIa3aqXzfy+S1E
1V7sE7yeOOI6QQc/DOHC0mgLZWGp4afuchaDxxJns85IaBjNyBEwMMMzP6KbKi8AYR0EpxwxR8Cb
0zEdLfaaSXVDAHiJWtBozLucvmwbul7OSzFR/AsqyIKfM8XmJkVxIoRhc75ogMg/NfEwzSx7AZCi
GOmcuJ/bF04ZNPoaRW1GLYtos0uL96PT6iU8Qoo76FZ5j4fwDEoxtfWOPfZ67nROlhIXYBaUquKF
C+rINZ3uzQ+BpVd9xpOsbYa4h/z6hjyUS0J33uta0fno21nLPbysT72tO0gg5RK/jRVUWNY8rBL5
rUdEbg/3gchu27x77UFKoxdAHmCGltQcEZs0apYwuspxDm20pcXclSU+XsWAzAFj7cAIpwH7F5sV
8MX4/PNR1NvdRxzG+Yxzzzuw1URrhf1S+kCghgui2epy2SnfQPz50E2i4LP0saNMLRRqWi3MtPAO
e1JNmz9YqfTER2PG6SPmSgq3nyGzcNOzI6icbOmDaHlrXh3Is5Hjjo88vlsyglGjOPjcfoi5uqNk
SDfkAc/T7T52y5B5DydvnUem+DO4n99isoNwb2HzDoF0l8NGWM813ovqEEJyAoyE7G9EaplpQtgJ
BLLCATSUGVTa6Ib7XbXWYz8nYh3UxKUN7TumRfczYy501pQOzF4Pwu81796sApO03MB/i4JekNHl
vGN7BzKUhGJACA/f71jrBRMOiLtPRUR2GJAWpLEgTW0ktfTWHbJDM0g1K6WlGVq4GVYlGHVLj5qV
AHlDJlLNl9nrSN+XIWncd6TdzGKfyMHM+lYZEj49CEyWYuGS9aY9Zqwxr0wzaBpgxA5Qlex1AZQy
5hjCjoZzGY3MWY4iNSRjyOcpIJKDIeptieESKOt8drRjlUACWoCw7/dlzqzvFy3Bq3wBPMysaxfT
PMBU19xDgOY56BhRjidw44fJvyxJjCav/Sl6uhwWUmHAyA1dSlaEnqG90i+am01brkYHYR8BbROc
yINeg1J/OWtsKa9GyFxDvPUUGz3nijK/zq4wnXWJ0a8QQfF6e+kG2TaVDo0K9MaIcAbWQQeQIeJC
qRySbMgr1yOKIHva3SOj4nqm74yMApmEOZEtnNSbr4oiwVrxKtiZUBXZ4Nm859rpC8mOQs6LWZUc
/pKnzLmEuoHtSKZVFW2m9y2tgg1SAv8kHJt/drGiYE+3V5UD4d4zM6+xv2E7XpxxRlFJ3RDjZgjf
jRJo7tj1IK6HXJ+Er5Jd1F5OWiz/wiT5FN+qN6ixea7VzWH7VLIVJSsUyuWbZ4gXpUmPXCEhz42X
eiw/i0zbGjkJtyLg02NF+s8V+FxoD/VXwccZ/uq4zf7v0okOFQh1hRIphplUOzTuZAFu0DGwBIRU
dr3gExVSapHN67i+eAkqSo4XfXtR1OPTRhTcwbsimdsJRodLwgFIJjFGm4vT47uJXpJEsl2Rqvwi
IYg4a2VcRCNnvfCsgnMOO+2J9c+lxdkSJookkU7zUSZ4Zojx1spT2D9x2reHj0C9LhMHN8I0tTJr
CtADw3il6yGe5AJCTh0pU8JY8z7RVzc+gIdzdjoSrVD9VRrrBIsMwqWmjxQDS9l/HUwwPMOn6LAm
cm0Ml70sD8QKzrKawpFaaq58+3XCGnXxCuMx6dOZ15SJe9m3JXMxWlHLMUfjpo0WjgfT2V9aB682
9p2UuZUjiU2SlwiQCMQ/9GQlfKIjj8ahUdyD9lrSxpczXIWGfBGeNDmrPnKr5/Z0EOKvnCz/lYBu
jJA86VQG1eon37yjCSf5yC0YFekronrWrIsqBTgWIyjxYc7GMvq9uvUgqRG7muVHWtD7MmlMWWPd
Ax04BNJ6ZCA0XEg9wM1/cEgeNcskrbVNe8ylVAogqf+FnmsLih9SwZh22SyVmRotwKhxQQMntygn
qYUz8++TG3iF+LilGCEOkzLtmLXp5aWFHZVLbWPRuXO0TaUDmiNdxyuqZkfwHe1ZxF2FAotWVpaH
73Q2kPPZVhVeYwMVGsJIScqpQ0M8cVUBgsV7D9gRZRtFf5vfmOfAn7ZoBYioCRjeQvthTJug6q/N
CQ45wUBreFPLI1zsSgGAl3aXNTrx2q9ko4Cl+/GGD2+u1CIXSRZB+aGKvdhxOW4dTxpg8971oKTE
ywe7RYYYsk0haA9HWnDLd8TsAHz4h7KQi2EK8hGcf11xPzsS51lWwofHeRZwaD8uyht9CckSHQn1
b/oka4BrAUEw3C5b9F2zpuGILNrUMj7kV10TWiVRZ9gSo1qRHAZpl5z30t5/fvqxth0KZQXDVTQD
afAEqV9oygvxR0glzYy3bB6bxV8jEw7yaYeOcjZbsuob2CENayrRrkNCtaLCRHVOZK4gBEqU0LPK
7TG08Wp40/9PcSHDo9FWNkaBtcrblBB2gszdXDFCNp5RUoCmyY8uKg215sWw91xM92oAnmhrdfMn
Xlh+cFjV5PEVRNdnoEOsJv31T9INPqt18W7DNKBCmPEnhOY2mG3VhSeto/U/Q1Hs8M6uKM3ZcS6t
s1vbZolumxOuOP8K1pzcDJDbth2uxb0E2cKmzqbyfpBgwLtABfX7hnCuLXpGjAI9r6yE8MByCW1D
VzsrZAQ/aZ6VxBsKP/g5kZ3+Eti6RRLrl9UiEulEGkxOAGuAsa7o6nPb4onpo/V5VslxF3KACG0B
7suiWxfcAb49s+iglgO8wgeayo0j7kWq2sWLSYhE0KgKeQKNOJPr2rE/oTJsNnK16d+/cmC0k1iU
L2+CGaAishDlV/DJ2/UVU6NghuAsFT7PcCpe4GIc3PR+Le6TAw3zQSr/sacERm5XiksX4L6H/9ah
2vONfkuGZqWmttwDr76+QvfbmzoxPKwvPXOpPgTrgMHlow5cRclpY4cDdIdZkMfvNn91BhZ7ElDw
zuf1th0gjZwUaaKyu0EOnUdIcPxhw4tESEP9i5mFNnbNbk4wI1/TzpcYgBDAHbAQ/u0dGhYDvhXI
dUXEJHQ5UmhGof2fhSrJLswIMxRQJ0MU3eLpEqEKyOgfRN1fr827JL3sPBOvCCAQAH4ewhKl6HG9
T/OL0cLvDOnvf6w6+iBcVkWaT57VsRO4ba3d721S1VBFg4XLdeZyDkJrcPrbNyrVxKfzIXlCSKrT
pWlDlXpBxn6lPy1sHm9W4QXvqTux9GEE7Nk+vCG6jgXAxFjc7hRzw4SyUCua4JMu3tEBYdnGJDx6
X4jSAKB9DKcc3sb7Kp56zhCiIuLVnvStvDAeQNemUuWIqWw9awPx6rci/L32MQwpEUQZgAh8nYr2
HtjMf27PGcFabjLb9AtWdXmiQSt3pu796NQF9I0vDzMrMqSXQHsLIt37wZupgyeJOnzpn6Ew2kRK
qh5kNGpaNL8pOMZMG99hEbnjRVFDpA+8EmMNGp4SsLhkvhxHuHt+hvneTZzICOJeCNjMwb3qiJ5v
RD46XbT5AHV1uZf0bAAkeIUmf0Lu3mq6CN9V70+JO7DjsIaiM1VuOQT3M65k0Wo7JgnOerThDSxQ
rZ67VqUs7mxFollaBQ+aN9SjGQFZ52AVXdJVgHLoKx3q1GiH4Mc/PFgGt9H5HUkHBV+EusmvDsCb
mWQFT4aQ0/mn1iK8vsK9jF+ZaQ3tAAxeJm8daXnhmYIgzACUZY66lKOSjRimDJ3PgCbQ5ut7B5o+
9jqAXddSeRJq5rkxIppVXcBZM0TiOlyZNqjmMkJEPeYVG869kzz4pcvxgOmQuFjOxfQNBdMO9fNu
19nAjl/LrkHvJWXi9KWFqpoX+u377YjHKE/u6sm1F/3uytLeyNBkD7tXT/Brs4+zYWr/ZyD/4HAP
ReEn6yOVOg8Zmc6Zj1Y9w+2YErRKf6qTPRaFfkZQphxc1sdr0Bdk7Uju2CgEW7f+vDv42myDMzl8
p1B0AceyC/FqGUCfYZBVDUK+uRHqvtbvZkNYUpN+LnV9jdMjWbNI8UikIDrjRHh6qvXiUB2pb68+
FZcSKmLorzFn3deU0FjpWW7tgyfOG79hpfWWmsJvysUZ2aK+rBHmvZROU/OCPvkISbGcoq5ogs0b
KVWHPXeFHIxysYr22sr0zxrDnFGD14k9gDU+XjnTY70FItAe6mn7RY0enUIpazKI6/URp5I8ujZ3
qyytDYTzOwlAC+tpRAyubpevlJV3bosxyN9ZSkQmiW4r1P2oQn+/2QT+bx9TXioz73/4I1at8wW7
KL8pKBQcAKIrVNXOKM940PUh3EjA7E6tlz5OJuJRSt15eKxFFrz1LHgCPR81RSUAPhu/XFRw91JL
ctK+/mWHMqWs7JTVlbZ3cgtnKR3YpfDDWlsxz/hSnf41+KShSjp4xewrnK8IMJasKjJOPeBGK6UY
v4R4Z2uLIPhwQ41qVbf9idP/UeQAMTOfzgC9kVWRwKzHc0mPeDnRQwhUFXQevRPOeB4WTlRP1oWK
PHD+cXVaEbDEOL1m33+9Ybszqt0p8MEGh1ZBYesBYFmO3DYnSkJn4KgMiKfhM3tAZg1zoYycjEee
Tn7kpEySWVvdInYwdJ45xU1Ewtb7oPZO9Kr5qJBkSihgcQy3M0ZQNpHDPWLvH/nUtuMmluJKN6gE
k0UVjQYFr2EivFDSuGgdoLHgBN66BHxuP8lq1qtWBZt3pSIm1eGfQRM21BmXqXDd05pT6lPshEsD
QIeiwMst/ihMhB9mISWz/uqTzmA7UBCfAeF1xn1hvamqcq34Xn3pSJYVcq8N0norRVhhq765QNDR
9uvoTfxMCTuAeRvlWA9CmQyvuNypWagn3xnJ8M2AVSdHzb+vm5zixV1NznDlbyufuvEzyDRrHnCf
yOpYVJy5l9o1KWQhg6UmKUXfE/Zqp0IWQYI8nXDeq8Hp8BcfFYVjK5IxGDSvPyxU4sClVWJn22x6
D88f8TIPZ4sdcVPED8Dm2KA6YsoO0LXY/N7hshiMOXy8WFxA6eNw3BB5J9Egs0y6S95/EBGjGxrf
vw5HhQzJIxSGgDTsVD4+ShNkDhde/QG7Z7wv3ucAfaKlAhp93LPTIRsybFFetnp7JiejIF69ymHi
vUuMROxBiua0SUE6MPcV43aAlvK3yEgC04mELVhDzWB6AALa0XdpwSFjNLfOEvHtxQqimZXLQhXO
IXd9lipqm8W/RSBKEoA1rS+6qeZ7ZV89mbDAh2cPpPaSrjV2bhWcVISGzMD2mw/4iHojL4Z7BlJz
sOoq62Es8yX3kLUIrNuazPV/kc2M+eVliIgOHwkVhWtjiaczzmUUf9xWLhtNCCx2kNPP85YDTJ0D
DHfiPXGK6I9G22Cb3XRKPWJ5ffi9OLAc5vQl3Rk4+QefYWSIJjiYlIuAzJ0ZmLS9UaW3OAmxPVs2
xy8bZzGdG/nu5kh8iX+5rtDHG6VsrpU5GzHG+h6+v5msP+YDPz5gCAOF0dd1hMI2dwIz24BpJo/c
JL37182O9HcNwysDqA+YGf0kTlYD2qAIVnomDsom4XhfzrywA6wzumy0YOoI3TBRdMNLBrYQky0/
Ds0+4hYM1Y31R5up/AElQJs6xZLexubrtxTmIWW8usGgLRAfLsRSjzv8DeIc4Rgo2lJUdbedmA1c
2hiKFqkmtvN7+Y/hvt/IqViiiXTirbm5MRLwyIM73ZLmeMrtmltlBIuF+t9mlMCXdPpGqdf7xiWv
bt4nvt4TXZShJR73ESJLiUobTU8uyTecMIyDwMxAidFzUYT9bwB3yYaJe6890cFOQ083W+QWrQK0
WDTv+8ptgMmJUg/Phxo5GJrXHixwuvVMqzM6qGPVnLHGOL5TdLn5WIMO+Xq7MOuN0/+989OcB2RL
RZMulTakGrsTL3TclMPDjlxefFsmAlmDOVKt2/6hm3hI2zEmz3GU5JW0qzK10YO8W9PYeA1l0it2
SzT7DidDt/ztsDEo5LmtnZ9nuKoOGiOOPitAMqd5ANR/R7wXUAaghwriLKYNgNfiKih7eaq09LLv
Oy9ZiodcUXgEY7is5Ff6dq9y5M9z4WGIRhtnwGnXWvo14NWVFEUBq1eqReyW93rn3GWsFQREk8hB
cBqGnPag00D1p40p79PUyk8jb05TM2lmMSkdbJDBOG4dRn23BmfeNm3agqeBJ1s+eafYsb67diwN
s2C5+WDMPNEOpfm1A/XUzXoCNBdPfxCdKkBNry6cQnm15hftGUEe9bAadzxLLoLGC917ZjejoGCO
t0Ig8CF1iL8O9/HzZH5t6RJcPqy9asTO/2HSusJ7m77i3rdS/y1eSK95axI3kC/q5C07XhpV/FZr
AyoZWfaiAbB4ZSqyBkshT9UKI3bXWAehbcgvt+wlQk4H38IJMkZxXcQ5mBKma1NzWQRM2WT+TK96
bEBEfM9EVdwmd4rX4UkcjJvl8qq4hHMLXNQuAvRHfU30iOqvNZXWK95eAsfC7w4OabkpeldzBjSF
ChpDoIR3QQ/OwH4XZdARp4ICUF/RLGuNPKF5WfN9LxAsc7p+QcVvaKxe4WIkp4f/BFq1hUarpL4U
/ufC3bOyUYrEBobrINNbjeI1fhtSdPTnnYVAAiYZLU6lVyv1WFTKxhs4BPMlWlZSZ9WLs323QYw7
kNb4jesB8JITmAl7+SFVcAWqwTDx6DpcQMMr0Vqr1CJ4aqjKMtAZtJzr0LWP+Nyu4CpjdY6FwtFx
XlEJyKAagC8of8XzOD9GorcPeuaUa1k/jkVvTgbRimqcT271FnnqMy8Ug8rL2HQV8nJQLxYKoY90
xj5iKacBa6XEO0FF2An1bcELtxlJB+STmsYkijJ/Fcv5LJDUz9gQ9Nj2rg1WCVfg/bTihJZvV2zB
YLv4hV9zR2nYSsORBk+Tb7EtgsNfaMc/Wzg5KzvJliVL0UaoAO8sXRkQiCJPzGLwh8MVhFikpOz1
X8ixvmAt/jiCMFaV+i0CGFomcdtLNhe5vKYrCkZ7guICBIrpHjt87LlNuIHH/2mG5Ly/RtqERNCo
pXIc1yzn2l/geNGYUZtlb6yqvlT2/+uEZfdjZMyZ9CEPvdsyUhltoNtD1/O1qaOPsrxjROFNisQn
lVNuLr2qOI0fyVpgUWJ7uon2MwH5bzs+HcJzUbpvyrvg2L95uLYadghQL11/MdAfy2oIl6pmqWJt
K9i5BU/Ay4funAwfHPU4k6ha1idIjf4PFAD2QqwrMLL/ikDgvjkz2ZKx7hPxEikYCz9MfZdI3h9o
rgPYtGjjizi+ViSkjeiyqiu0W/CYDZqHg9JRupCC+yhk1Oj2Qr2iiVtaJBNEBSduR7aezBpYYNZZ
f/wQcu2n7GfyXPmMSqGer8nZTO+ZapGHe73VoprqU1Y9UF2XLhpCPNgBzGmI/oq3ZpNSiA48maV4
o63OpLKWmDX/G7tMvLBE/OrbTHiQPU6N9nklpkFUm/dijl/14baRM7wP+bG4IHjHf/rJeazLwyUg
jwjuIYUbwK7/wm7Mno4IWi27hByXNXtU777TZsSEPGCTRaBR/pF9i9V/QdCX4/KrWMWLPMxrTabD
PAFO/LEFRmBkL7oFCdqQaa/h7T3mhYdtvfFlHOgbrlpPrcrvSSMseUfEiODMWY/t+/grqlHbWqcn
AatxDIkR/K/+ASldL/9CBbknUHL1iFOno3RGNWoPDFJcOOoBxBAmuno9dQ0Dlj8jeeT8jQx2tns5
FJbMpibWdQ43amOz04QU+LJ67B7hoPCrMO+OQU+IKw39T7vAZPbTJ4wElX1lnMTkoE+9MvLiUGkw
j+E/pQfzuxs2IuWckQK4tc5vYgHuo2a37SOeDXtu09kAg3SIYE9TlpsnBcfXQxE7EhBTkfAubtpp
tkIqJBwDiO8qZBKePFBV0S6j621mynsMom0av3T6SgQbGGsFzjWx9Xg/qnifGdwXoH1vAzFG9psM
t3gsRSUSR5aFnySnJe3L+mHQjXTx7gc3V1F1i/A0779nmKu3yrnX+ObwP5MePP6X1bGZJtgh0cyg
xJzdUOiyj4XCQ6TD0KsxkNPOcLbOj4l9wWEW18XkfyTH5UHR0aT9fOtrIkLKCO5i8MXQi1j/dagF
nQgNRN0NTMnTF3UAflQv6Lqkr+vT1R0U2Gp1/s4RsoRoTEPP42VjHMUATI96Q3s6pATV0RBzfGfx
X1jQlftjTXTGwZnZphjngNz2eep20Xf6bXBU2Nr/72L5F7gcEJD6AzesNKg2tJkVQByrs3uhK2LJ
u4OCfERzuBvJ6fZEw+3EM/EVmeOIUYAUxPZCJNzIxY/pgTSqzUurw6uZcPdbyeVqM9FAeL0F2LaN
SXZ2LPd3NwkdwCzfxgU1xQC67gARG7QJ2K1ybNxMrfhdDdT/v+q01vHyXDEm4cr33sU+W4NS4Vna
oJzJ1l98vJatD7emFHVk4TNmYmAiRKrLFdkrG1jT00Z8k+KASyoRD4u7gGk+mPkUTGZS2UhW6gN/
/G7hWEfjZVkGUpiCOCb07FP75TphqtSva8oDANH4wZRACTY1bPRpdy4hfOjo05M7INW5IHnE4uGt
eDWjgNzQTw8N3aJ1j9j+IrbJfX8KfeAhYOAAV70wFwwejGFAqFbN7EheYqzucMBPPIqdoKfFeqUd
3MI5JtLTZSrO18fYPY3cJWv3o7npEl3/G4OK6akEnYuWfnPyArLN/zTG//RR3J5WIwExTpRxLdBK
n3RxZDT9lGfJ7r2wAU0XYxzg1MbFFPWwYzQMwLnLjJ2LLmw0cnCAsL2U5IlXAVtW59xO1pn4exFE
3uShQ6IuLf7kxQPq0L3is/cqoszdHZr0MafP3s3qKzNTXYyHiQUERwEy+NewuRU/xQUccKh94YxQ
p6NI12+syijEWPcd3RVR0cHvPy2UKL3HgfP5t8bvIo8j9oN8YKdeCGWm2WLqqyyiAeROJb8QcrC7
24izf8A4zc5A8znwL2BiCuzInjl4ItAyqqtM3kxT4hj9dbvLYrtNwrmae7GkKJC7e1BINHBCyQfF
VPuMVLl1WxLbujMn90nS96opR25vmENbScXr7u2nqZS6A239jurg4vllW2uvMGefi4tG2apPcHgL
NevYpCdGouiJi/DyZOGRk8Rf5dYF8hgMqLFnGSPC7pTlUFCnuegzjpTmh2VfziR9AoeRHc+Z9Li+
8jkYF+qJm+adrQdxgu5bs3tHEProtnzGIjTiuxknjTIfoXwuS3BdeIDYIntdsEMS4uv7iQlq7TW4
qWr2fjAcfbHOjoCyyv5ouWAax1nNx4TKKPJlpBj/xj6b5tE+36ozr3KQljduEXDXimuXNTSnGuxr
bRBpJ/jtK9Jg10CsVGzAYh01rT5UAnINE/6H1xxLA4QCjb6AXjxyP0SaU5MJ0yNPn1bvGPLq2dRk
8jV68cuIwcZhdSjr+MpdfcPXlITI1zRo97bK2TPJ3tMWT1yMeRjRd2o64YjkViy3T0W8LZNYPrpT
SsVqJ13dD0m9LYLlyKMB0INKLmz5zzOCUZ/nWRu9jzuHyMcG2whQ0zYOl3zKF53c2S1yprS2zwWU
NhZePFSw+qDAH9zRuZAJaLp9P17BmqkBcvRG0AIoilA2CSI9u5szemiWQaOAN6z8sYfZ5FJ33hXB
U56jU+VFHZxpwqnzYUWN27eptMwoC0qUy2SkmO1wYl0cUZuHcNa2kjXdfmxUxU54hYK17rUEBkwt
6kKkQ6wGcYbnYZ9loDbd6/264Cl1ClPPI8slDnVpbkm28Ha7va64thDRQXKZt8eZAOdZCFYm1rDO
qrCgCYBd2eZzzH7iqGYMKeaNRnRceO23LAX/jbxTcjMJVfSYlV7k2sw/7dsoPmPC0PdS0YKeyKKV
RQQB8HwrMmFM9sJNg2iqNbcMQ5gTYIGbbNTNykNqECmBoER2s2lh9P7yLikEei2neu9B32lyqH9H
E28parXPHiXF76mjzbg9kGmKpkP3cNmfF2Op+jLFg/RZepncM/0iO9b+zsMWj8oBHm+CwavlGIKI
C1ZFrzO84sHsRcJrs2igr3DkNodPre5vkdJzUklQkfWU5CB0nRqnlI+1Kl+y03S7ckO/usCPgEI2
Uo4nsKCrFh0HrjKn5itEfoW2jHZbGxgGtNupK+g6omGSMS+YOET9eLY+FwwVNnG40aMWtw4cRkIi
saOAPyudo3ayBMjGSME40fI7N6nF3rXoTMIhZS3p+sh9L460336Xh/QmDl+/0gNRwjDFNei8IV05
G2tgzNC5gwlMkY6RR7KkoxBDlyLI498fu2+zKkTZwx/2MkURvFsmS532pqGrOmmjLB9D9dD2vDea
2AJ8lBH+4bRcjlKeSgVwIJO0Pz/0ClsxfBI09TXLP4GffRN87baMmeTGdIzDHiV6DoVWjBZySAtd
GZZmT0Z/n/4xlCqWVZaONRGDG+LIuOahlUoZ9pu3MLNQ26p8cR5i5vm+HhzifcGj5zsaeMdqP/0Y
h7/dNV+KvqGO/klwrdHaBZ08W1TkKFvlLlp33Vqs76Zj5rNDFAh/dggWCh2yvPW+n+gfnsB/A+Dd
cFjWFu39zYJ49OTFs9LI+65v5A9oNxz8rJk1FYhr2ytchynFnYTHRlWPA45iKoow/5lr8HObeJIW
DRFgjkMem5YZr9ivlvrNGy+iXSRLaE629YEl8MXfl47mucpeEqUEY1Y5X6gsJJQJk8yl035X3LXw
pCXpPsnMswNEHFOW85OZEbjSsh4Q6VtQa5hNZPc+Yu3iwCwqwsVnrjnUxP2MUCG3K60S6OGWePEL
2TXyTwL+ZL9kjqWn3oy6QUhe5b0KKtg5Ik+2BMvPT0fEsS4RDDReFbTvZOZcH58SjkuPR3MptBnc
gKyLY1/wpoI/7ZJjqYF1PUmImOhS+TEyzRVgR8KNmEV17UvjYSsp2Bt/CLcMAdZK5C5pgSA57WsT
rxrTwAnTiP9DktYwqNRqslD+40V08OKjfMBOXlX/sbnoDqVqa/kp03jmli/eB+6ukj0q+mhAxMyH
81dHKhrvEBJloNFCXcM575Rky8yajwSPhPSX28x/uNDGsW/FXDg7oyAy/7+QKK+W1ZLPuNkC5sBM
+zMJrtQw43Qo0o8SQEfJ957cptDreLIhsA09Yla2rXiPzL5otItL6xolLEE2JVZvdWax93eFltNR
poemr4CArBe2k5UlTY3Vxtx1LdrfKFtaMqcSFSYd021hlpmQPB9ud0g6iPGl+P2e7jGc6R3QlDN9
phg7XqfGC+V4mFIaeEzV3zpq+CE+FRxxGC/Uy5bkpcJJkfPT+JHgjvRxi71ZcQYURbjicBNlDUjO
RDG75bL/KbckWmNz/7aTjCCjBydCmjDhn+o0p20lrAh6KsoRpA78t6txkM0CUGD6eUR59DBlqgQf
2AHyXXFFwu9n9zphMhGFtUlzWCoeHnlcgROH1oZpBFB9r5JosB2H+ju3esMnvFWeFPOJvXREFm6B
SpDaJjeUr+SeCd63baxARvQZ7S1IkGHTwe8Lkn8f2vc2clXF+bcE/lIODt+J1GbALU9x9SKFaBKO
QkYy7Y0RE1MVbmLPWGbpV4A76Z35eWaLhruiuxeuXvbUT3iAELfy6uMkgsApS2XMYDxYgImmbom+
TWJU7p2tnM2/oDBNGY4kbbWqD6SpORcS26qSZ7Jf/tVJSIc2APiLpKYRFRow+guttz0mFKwb2RWn
Yvurvlbt7Pzt6adnWb6V2bTSrY2KdUjM4dDPJjPlg9VCD9+PjVmMTM+dAHm62K0uxRgQOoTptjCP
bFoOx1gwdG7204p15WjafP075YqMUAGhDH+ZqY3aV0BYe21CrmNB6autE8K1YiXMknnXrUgK0Bln
gZY67mCWeZ7YsohSwjGU8ax3TLQGgN4tfnyK2asARqeL6vGqLYnzSSV821fhKR/8GI7A/z7CvVXn
jRVvQNVmPm2QIBnM7j07rN0i2pGzwtRKZYqLLc1yTnSwolMpqgR1LrTn9zt64838MT3uHUwmy3rl
GsCH3F+rLUHSBgz2qEuedOwpZjm485YNqSGOQt4h2qaVl4w0kdIIUkMrw4psnBLSDZ1zZaP8ZhoW
PmhWX1jYHo4gKzRAOiDH9EjSs9nBd/ht/+8el0hVPkgMkG42JmlhlgjvgJr6QUH+L6piP7XHwQ2Z
k8LasC8y27Kbw007CjmHcObXebh9XBVS6m5GaFjUcWld+vIw5KUW+pkKnIVt7DJpi8n8RdwOOp9N
r8QM21zmhatecVD5nZIPBuQi4+o0XindGU4mg+eSBOr6A+hHo0O4YpmEtAsVAnRJC3jy5ClbXPW/
Q+geKxdjggYSXJNwZBcwOUUs07q4AgARk4R9KDp+JBTW9V6MkAx8oeWSPPmgso+1R8vM1i/01u22
RIZlU0TOxKCdH2OXhkT8/omY1xkRnfELfeEMD2dggrSdJ3XcskQvKIHaxQcxweD0/+/3wgge1e2y
ZasqXR1Xpx3gpTaIRA/2FGCkoCg8o5DcGeBS0r6AbyIcxXBL2GbMHHJe4XJG6Xwgt/P7EG1iEBcJ
NXQGe6maqDohK12YAIc8OaEuoSxjk4JZDFz1LqkGOvi92L+A3obrjC27OKB6BKLYKvejK36Qxr3E
1r2dih+aCkPODKsgI/y4evW9DpHXA0e2uuzb4Xdhj+KqQpF2TDbIqO/ut/ELvVcf6ajEClStjHNN
hYVXCbbYrDg08b5CeM5XRLm0Vr4r9nGgjP/6ad1LYOcH17qu6NHT02J0rLQ1vOWT+5EteOVbSCOO
vJ+kpicyB1l7iXNTDyymfnXc/rUxxXaIsghsJ8i8H51DSVmrIGDpgDq09tIbVIy3ssgVuC3V4D+z
3j+RLSxZ4Rp+sH8gWL4xKOLJf/cA4NRrAqqnuCblVPH3ZEHnkgwi5UlgUHDzMuxtQRA/yHeJXQy7
7cI1XMFHRm5NyNfbX9UtxzkaeAyameQ80lfAsrROARDLG1XwYCsIDqdNoUjAQKvhcECGD7aTIykp
tYKTO/vuYJcDIqtD8BNz/U4nTZWwGKBSAL6IrozMe3qHfTNZdN77eGAw6Nk2MyurNMmZAZDgEfIV
XLeE0J4uqjuwfxtLbKXsIhNUc/5S6G30SK2psAslO8Sw5VGdNqODqv5UIj3zYJ3yM002Kls3oOJK
sctISMfRqJr6xUiO7WqI+kSzt43rC9lAicQsXkBZC4ZSeoo0RJXlosXgxO+s/tojl9IeczGcAAb5
89ZdZ3xD9dFGTAPQqL12ZPuJ4VFiyttzfF85/ezDAnA8/KGXnMjbqRpGKT4Qt96eYxbqQd1zmSX+
TX98woLp4rL9i9zevOV39YjLI3zdcWShoXrE9jBPX8azIsOzacqxXziSYA4sBYZsw+7rRPuXFgQh
XgXlbJ3ro9RMMlFkYE332V3y1PBF95EM/wuo9DPuIlHWKKqAfrFNFYKbxzE6AeU5CDQs8h42K7PF
B3NMcjstQy+5jzqmixRStEQ/PvqeXZaigj51OGSk3VQkCXA4V6yVOeNIT56iA2eoeYPTyv8v743v
KPJ+Qvh5SW0NsgQZvr52Dn73qDR1rqhQj9TUWLqMAjGzTq37eWltfWdLW8rrAQSi44GNUyi/G3uT
IlZ+zCkUH8qBbGt/iJ1spFm1jVeOG+e7/hdaea+D3i4uICLMYDC4QJuzcNdyQzFuxWvg7HyHLFxn
OyRXg/yBdd5GMTNEUw+hbH8N4ihj56Ji4vsEPETBveFYRQTIiQV4JNvRLSvGw0qSgeDXmI4YtanT
8ydqUjUMGKHPooQ65q3mZnvdaROrdjKzIMeO7ePQFOzL0/CUW11YANbWTUeTVEW3SvFMG9dYEdf2
1DYLroQhdP8Fiu0fqq5bqpeLHGhfYN9o+HD+bTNJ+XJWPJNf6ykrvn6YyxKLHrGzyDOLgS5BlLdE
WfinLdTUzKqb6MsGBJTACcVf6KZOKlM7R5t5bvHMf4radoBpJqdK2+A9PHZSu76J7A5/JPyuP9OY
QHtIuAfnfn79lwvQj4TPXxNU0MWENEd4qGZM/5IAMQ5Vlj+8iQZ5qXTI1YlpCa6uRCmgUeow+5Ji
gMg92IL5p2jHW3Fwce053ma10rVbkEM7Tk0A+ZfWOFitddkX1zWgh/cA+hZkWx3edNoPKJKBYrD0
UlO/7Ne+Jn/nMVVzJOskKtYDgbPLKY83c3IcqkrutgZg8CA0ACsGOai1o9hf0bvnBL3Nd0DgwRau
3cKOMeAzAOKu6Y1pLLZFpNNGDe0pmzWy352SU5hw2pdOX2NbuGDh6GdzUQBE+aRCKQNjqdqz4TRo
Tnj5+VpWZbHhI+Kw+KNkcSXTkyBi8gjaUi4vcD6fBxAr9O/wLrG/2ZLwvr9NJp43t1d5+2XfErQb
8ENOedpXX9tV97eWHpExw/q0H0Y16OKJkCnIiNNJlj4NUWTq/ghyDkFmsf0FjLYvjBvcWLwPbWZQ
ZBuN4ejZarh0mG3CnaJt830YJOXB4hruDNXGIXmFN6R+HMY3sZ7t40Odf7Qns27WVTUXZbVofIY4
Fp6onfzQKo5JhBvjFj2ldmOzK6euc5A14REIy1y/JuQNIPYWy8I4ZucVj+hGb31lFpdBRuJmaYPa
XuCpcojT069yoF8PDKl8i3E+RIAyZYO/LZGcOi6OMoFscHgSGf4eIRFvC7C2kHX6BzO/Wb7aTbsY
vYZ1Unwcg6WRUZwt+QQPPRXC6xztK6I2nnsLF0anu2d1jyJ3NVwtpTXMpsagJRVR42YuIFIgvN1z
VNY7vZmMGGc1ohi2jWHS74+S8+nif8fA69nq3vl44fmguj2eWFkdQluoB54XkJLeMsvrlMV6ltWh
PGmkSTnTpNnIa2acSudWF45yYKPcTGpqVFQGsGmFDsvL/lqnBwAC7j+nDYXskll1G+J/jQZkzmzq
DenNpa1vOPqOXyKe0rBKQmGjrHEkxIfDAjwNEJp3uAt0S0cVUqbT295YCEyPYhd32xuBMOjtBKQf
+eVWDlr6SW9qDaguq4O+emzVZPPy2u7bFXpqjAWM+T0ZoLU1HUsvnVXgy0qtRCA6TNtwtiAvQ60l
HrgahkAUd0FBoeTJ/Mo/4N0kEd4jnNrP0IR2tGeDUSJzrvZgGaS/dSogqGycGX3n2yMFHMqQN6MS
PBOlxWtTkQlWFKUkI9FLV556PNrEFCMFdJ1IKRoGsz25+mx5QhHn4xfUAA7czKFmj3Ay/dZeZJpq
MzHmPW2tt3nZIThQ3QU6yRnWFOe08tcxbUA0ZYbxev7va9zjIf9DicNgdu1MTErgSyLpN4wDIAI9
nGR7fmOVNNQKGhdeUgs5Gm9SD9AunLfvMHR+EraHl8mSY9ySIeoLWvTDlOKpF2x9bJQPR+1e/fm+
99aIxVvS4QcONOE1ViKdwfkY5EPCBiDIcVUIe6gEcAbPxxTyySyvs8KrDSLKxIu19IaPRbA0lcXr
mSNff0fhiufGl0T5BOm3cqKZnb+dUk42sh0CXkkXzG3LLdhPCkuBmHTdJgOXxqY8maXauTjOd8f0
TTOvbks9DxbvPCWVgkGBkYK/PNWcOu+R/KxZOcS8tDxLOL2nI6TaL7el9EzDEHG9AFqsVv+8GiQ4
E3Lq2ujtzgyliLk7qrV+/I/rev2f1Arm1NI1dyfl9ez69pRcj31QZurJieQ3L9m68PFw6wnxRkVa
CkQNLegdpDkoXN0vHFsFQm4wnecuclW9T3D8IiwVBlBtF4OrzM3a0mJGiCw6IilVabwdsFL6Eowv
1SA0iGiuiKoSivsRETgoGSzoAv9bLPtUv+OC2xLMYRexqiPCtx+acLC/+pWJ+KpANope39JJOhTl
Jxfx7PMN7qvc3hnxFMDXmcHzosQsMbcRcqLN7QPYxL3sHRPf3EN3vPV8WpjwfhxalZALoo7CqyUs
JK7my7EdFjlbuAYMZQ8A+aA45XCH+cSLKb1dWJabjerUaWQWAshvb9V5gVmv9zY7pmi3uHK/IZxp
bmJy7V2wShkSG5mdo3NU8TyChf9JyX05j7l7nvtETP+4W7wszmXrkxPhcudaNdIfz/4S8uEyBAxU
27T5/n02DkiBnpNh1bjc6BiM/QUzi+1CHXFz749anWwvCVJYFINNycVHqZc8uzzpm8R4kvpeAm7j
pbBvr6qB17mmqjtrFC6UUJYuwwB8P6TBvnGdcm9SEzHCPO0C2n/iqWr22V/iLNOVZ7Fxzfp0irjX
8yMAjG4k2WqLzo20j9A2ejbCaIcwOZ7/wkNbZac3uCVkodcKZCxzWFt0hMo6nok74NGc9AxMj4Ft
Tt6n0mRJew1R6eV2R3eul6CScUVYFa3C+msn9OX6P1gidO/xg7o+TB47E125m5czOVxqTaLP4VvO
yLXZnf9JZLqEpAHZEGy+Z1FU7cey9Rm+3PJFKppoITph8nPO8E6mH0jdQbp/sOKahffLaxyB8vul
ZlrjWYMdIcrXeCDo6f0jUjIfc7g1YWwTIvxVDWxnCjCV5NAIp2uDHT41gJ0JXLpbTX7mxJ6PUxk+
QOvrU+vuW4ekY6KebO60Ok+mEcxjr3r4cW8g5cSdiurruNiPsgLq18sY5Mvkd08ebXkyOeBuh7wc
0biiW4gAm+gUd+8VKKOSoZnj4df0j4qtt4TLzSDod2HHbnDgzpWf3nBzv466dlH+FNH3Y9OClnHI
kgxyx8lfYHBQeER6q+b4J32uKkl/q4wJ44yyl+AIkeBpUAmh56g22FySN1pe6l9vPhQKMk4aQgFc
9eHkE4qRlEO81Nei+cX1lTKTGhdwNTYIibR9gAMQnxw5IbwuPn+GpJl12zjtfAHTGQzyWpalElKE
0GvNXOw4DKws4exPMcTi9kjYUcPkmDw7VwV0AGG1Aoed/ifeyqNbL6jG7PgEE84mD8sN5AYnPPcG
gne4+KkgUEEot4QJ6wIGgnuc867Ae/S9SkIk4YZbaGmVe+kBc4VMhqnL1XZOt7DkqU9wal0DoJNZ
fzcMX68Nlg9S6YJMZ0cgNVOt+BVKBOsOvOIvmYZGUS9VPLoiQoA3C+7b47DVRr81npO7jC+ce6bD
GpmG4BdhcO0zxpZ0wvonpDwFYOk0LHZkRpyrM76mIwBLiIOjDqcJSv73iWL9YLtehwQtN/3yk2t7
h5w1SGBpjdhsXhm6CvhfRrFAmnFb8O9c5iysXsFKLPEXcBD2yCj4jX6qjVKnFsVBy2ZiP3vf5Mog
iZH3dd2t0RRSPuHkJXjw9IwjB1Or7cG1w37JWNGQ0v1OUzFHhaOGgesoxs9TsM4ePev2Bjj7iCWs
xTmFhfaRNN7pZeQ0h2obe8WTJ14hoduAVFbp1BchDioIeDYwx7Ifm5k+0CziYqKRRWoY/YIXwjVe
lRNWgBBQx5lexpoAk3QJKoCxffUfYkMlNm659Emn74yWkrBpj4LtcZ6OeAAoSenIITp/dPazF7XK
fP/pc7QAsGgn1IamPLIjmAxh5j017MlzsSPTm1S3rY8yg4YgLgEDcGPJzExzo3T1AXvdybPaHoif
CPXYgl6iLzMy7kdKOVduDWa6RsaCOI4ioULcIOFNY4GL9saLlLGxS0qwaZhRjy8TU0V97ZtWWY7M
HkvIDc6SlMfb5z9FYMGy8YRgJj/ei/ao5CC3C39H6W7NbOBrAQWNTUhBWZkZPQ0JTG+oHKLa4yMY
dlzYJ8E9KALiTRh1Zj2ZUUOsBhIHX6hmOwaxMCJA7D3TVoQiscxZZVFrKw+Kz5IllbRqJAqZgK0N
GmjMpIq1maGpbfRgcjJV81jUNIZB+R+XGyMgHkrdub5DhvY5Y3syo102P6gtHLLLrAf9crFux8xb
Zj69n7uDinMui5myyvcuOjimaOxcdtNHRYTW+GAsE/2shF17SL2WEMLLey90a1eAs+kYqJsifrzf
/R2hUkb3Chvpmnrf5YE92PuVAEEuq1QEf8SWIQL/kKov2lMrxNptF5nvD5ALxHWGuPMOq5okuhow
mnAZcx5WLJG7cpFpRqMLefciCga+uNB2OtRORStEFYQi4tf3+VJeFAa1bBbDyz5Sg6NZdyamWxoc
pJOTlwt8uL1iscZCB4mx97g7iG/gwdg8A335tePtpkc9TeulCQeB6XLsTTEZ5z+adtmcWCPn/hxj
OnDWxnvl1uitSTGY6R0lktKrQMKXd2wVJqeQ7KW5TVMuQKJKKTauJhozVH5x9+v2g29X2By3kcN3
aXSWJwm6pkXl4QVBveQ+EEQ1AgPXCE7+cLNuXjo+fjstd5X1pYhM4RovGT0r7vB4AxkZOqicKrPD
HQ8haDprZW0YFEG46OGddHFHUEUdZjOXJVLFNBSZn8z8dmnFkFHXcGXGlB7IIFN8x+dQpqD+Erjy
hxzJ+9FexKlSKpBPimo5ilnd+VJwwaBB4bEl/zoQO52tKeqiTBIajRF5nSeRw/rIdIUSXK7YjjL5
3eSjmdV3PcXYCwRvW/qxnmb0gBaAlgIevRVpM7wqNPMVaatUm41kR2HaDR+rdWySEO/nljfD/RBK
Xci2kOehaIHAEK3mlRYJKR27jbb2Ljyp/MLZ0LaV8DD8VOE45KdpGYoL4J3uktjBG6h5duTh7p/w
ZZw7Fg6vClJ29p0cgPr+CbsiIO6atI7YOoQcxpimsRvcSoqEswA/6rqtyirHAq9KaXFw7oglGKDw
HphyRNIUTv1AkPqnN4LXlxO+TE9eF5Q8zNRcSQZgUrj5qInmnSreSYaJY/2hVeRkymmNZjds0ujf
INES/rQAoy5+oxz28wgxrH6Ejom06i0zQ86DFNTOmGzXm74yu3rfZx/C0sivZuz1q5dGDrBwu7sP
OLovmeIOuC64N/HzB4k5XP7aPU0UudL4Ig9fv84KabQ2v7JH96v6ggsyJCz/ZgLPXubuyI1KPhES
YKiZPx0C1ia9OSxSBX6I7xCRBFQQUt+WeNTY/Xiq++fJl/JJuZBUl8ZvzRoGpo+m1nN6FcqX4I1C
QOmM1P29Bbv7P0MT2TUFaAbEBdwLIP/eYR3jdDqfCENTDQVpAibUHFMO1hB3q9MblGBvn1Tju845
HNB4M56UOnthFACRahhwP8DlNhYU3n/BT9FNlORREIK3qZcyXlRkI70LXOPXuZGTkQi7IZ+0voB4
MfVwy04204t1HJ0lJgsBNBIElBIbqZSoE5/nr/3BJS49RfrG9IcPzM5ifNZxQ5dNejAWc49nB0uJ
D9UIIgW+56+zjoYrGmy8xbbVI7DFyw1+RCb4oGCg5feOC4hifg8x+u+JGpT1CkIwis8W4DnRnHwu
kgfwrYZpyIOXJ6LJyij1ahtn86HAsjeg4W0KJmgfkHn7q9FZKAdH3F8R4ANC1YbYadveKLnQFPWa
znJQ+WmjCMJZAI2tIuHlD5xP5NnVXURkWy7hI+Brz+6f+iyLLJ4YspCUfFxNwSJ+U+fzF95eJXD1
tYuVg6Dwenb47mH1GUCw9nO65o+EZEg69PrCry9DO116apJPN8OYhMVFN3ro0gil+40O/X+5XBoH
fawuCcWgSzk2Bkw/BSIFUIsZZcL5wkL3OF5SYc2lHRZp/RsSB3mBSca/EYvVE5bx8F4M5rWrI0DB
PuaNRXtRzUoYD4P5fWT8NW49ow35XiOw6DSXHSaQd08LZAM8C+co2Psj8aSHVuCVgRNeW8sY4S67
opD7MwXuKogd+gglu8VrIF+ls8LIdYdkKvNVimL7D59blYJeLKT0RrBt8v14vw0rrrNriYmJ24vv
OtdjNY/J8vphJmfRfpiL6IF5mu4WlL8TyaOBDpIhr8yekZXFxYROpl0F3COFH6ITOGfC5UXLTdrY
weRJT++72DZv8qQbaAGEDr844GfiPy96MSHbCVYe9ouF+rUyzX/C+klWUiQdwN02kBtkt0vltxRD
TY2/y5po8+qhMeMV54OE2Me1zrsCD8/kToeLzeIiqtg9+QWGzaX4oWa8zIltlagCoDSCCjPakV5G
IAbC+jSgbjCvQOFKCcIrJiWaFBs0pRtNjHdKYJHe6huRFWTV+g6kWti9D+ecQ60zElzzlZuE+DL/
pDH5UlQZ0xys9WCQUmRsTfzOO5DCRV41x21wfXw+PrIZpCafyzDll2qrcTlLnL1imFKzvLa24y39
mCJBSW0T1wWoa3WfD6DCchHUnpyt3eTqAr6Wd7kRkPz5f5BzMcl8fTLKl9TFo9kdiWfng6eAhETB
Ewh8H9LHZKe14VGSWAk1FP9oSjv91EwdwTV93emR8VLoDUrvUl9R5YZRXGAzsAIZE2jk6FEmI7T/
5PUFadTUkamiyaCiflojZPKHL1HnuEbV0M5vFyjbUTTdZxSwpZ/AZA64Y1zdKpfl8bR2hUgIDh81
EyGwSOTPJlYXF2y3UqIyJWhIxzzu4ivh+8uznBfaPBp12UQF/DNP+5z3gnRPtce8tmG6QPJPgcrk
Vdq++B+uilUgokRfXnN8oviRJvBB7Rv+N1WLeWqxhqLkGzRn1yYSh4MNRsZhb6JI7uIhhr0VWO9T
VaBRSkx2qTDIgWnjUF3rFNC6I3XYaa05s8BHtOjFs+kUnKfSDMWNmMvbJRLlJ24KyIPtjkdvSR50
6ruwWy+oqHOvJRj3UbdsVTnVYI1EdA6kaa++IyZOXGwAJbbZny8zP7rSnkyqR53VpDzTJKzq/x6n
i8ca49CIMM/kmtCwodb2RLBjr32SfhmxanZ2xQ8h3utw5j594HYIneLr5osoZJY8q9p2oa1y/gcG
b2JZuWMrQT2FB7/NrFfMXanBzXL6kMKrQiAhCThAJTxV264FVHKABZrs8fFlAaBr/4AuMjUSqVqy
9aJlLl7h6Qcu1eSKd1K3SvF4TmjrkA/xFBw7kGg6Y9i7UrZHhrqVQuV6aMcBY4ccabMGekg6r9v0
5KXREFWGLUaYF/f8DIsSxiUivVWrBHFdUhZs9vATXadfGTDhEYoVNa1qpjfHKDokcovRZCvwVVc7
2cyD2l89PMCV70kF97HWGiN+qlM5WfuqjEGxO/6ctbN7AgRdp0wefCnBRNLcOnJvu1S0+/8e3QoC
sU8zgpYI5oQhsnJdUUPlYb0jbh2iodsLol2X8+N/JogiHYt4+1eNQ4KEofAXIlXHBQfshb/wqUyp
1J9eyyWqHmNXyzQ7ldBHtRMXQ+Wk0KbA1f8COHgQb2pcRgpxV0niERDJ02u7E/X2rUVC1xZ1shLP
xUjVPMVgIpl7VSx0RW+QO4yOH+Z+PAQeQGDuMxrbOTuxfqTGnz5eC3K1dRG60RFJkAWY8UmG1OgJ
RYXmVXQUNCObl9l0GiyqIcVWPglltpG+x3c4UvEt5NEP147/bgn+rguMQMWSCj/FX87nbSqo6a5R
CwFJXSLHxwlbhQMKfYcOUq+8hZpfxoTb5cFLaK2BXeyju25VWum5+oHHlKLPD/7eg/pQaYZJBH3P
2U3CS/L0YKS8FnFrRLGxcezb57i7RwdCOKg/ChVsCPXSEgPbzAp1jOsAbCbHFJhgwTCJrMlE/Sqs
4WBwTfDXa0dnKEkZ+HYIVOqYg80ovkzvOc0w3dNK1sF17GVsErXQJUNT/G2l2aSROtVBIx6KzRsn
igrVyBw/Fujc7CILYCTmHgA5CuoTcZxvycXCHGp5l0E8ObMSQ9opYuBr6m+8krcfKbVj23D3uOv8
XSwZLcb8EwGa3hKAfQymIYlhkOEHqmnLxP3j1JvxNStD/NVqF0c7SlTOqZMsGQeur5CCaJsqQraY
egg2ndwolPtcmFp1CScnHNWuWjGwjRUEbdBoQF2layk4JAKv9pO7kGktYGsTzvunhBcl8JWWMiIw
doYgz/MDxD1i9oQ75a5+jB1yXHdGk/NYDK+0U8V31rvARPEQhFxEKsFiLuO10QJTxW720TrkUGqb
vNc2/8H/XGcREO01xgMnhb1HrvAdKvExoSDqKvddrdL4ag/2AjtcnNJWBkqBoTHbzkK7xs/Zzphb
lGxO22mpQiW+ZAkKRKI8gR6kQUpZa9lGTdqKZsjo2H6YaXYEDCPUNgYFNOT0pDW90T0Ep8dP9Swt
6A0+ZAfQLBqje3V9XEfT5912yIeEWJeIAYcBfDt3j0FRPvdO3gvN4BcICjhDzUtMxklTz0FZmb4A
fRz6h+s/y6ZPHei9OCZpNcFuZMw9B1hsheYxQ9dUMoWYWG216/UnLUMRRe27Z1dcvDS//MAspUVT
JpgFfixx1YnXe5spo8xJOWwm9mtqoFeBr0dG9fDjP0VRQWmcXZze+Tr6MQ2SFii6GoC1fWoAm+W1
FzPzUQQF4yRPsw7I2qTL5kAcB4N9CpunMQU2b0jt+ICP3ulF+wraJHB5udt6D4XUy0xc/xw6vHnO
A/UvcOxd3VmWwtn6Hj4qtocRLxpHlCxxTgqFz7Rw4iA0QcZUUh2bxa+GmdXM2u9eduKpDpBj26Fi
vP54nNef+7tVwYUt4WS/bYGaqdBYI3UoTnXxscJyBagYnaXNjEHb8CHIQslZmFkX68E8ji25Op+D
sZW6seFmg45tatjy7MoQEkJfuflWfJR0AeN+QpyJaOIfXIeNUKUa5MyJzP1ijB0t0t+gCdwXrX4w
Fpb1vPXZLZJ4pd/2+KLsHJV7opUB6UiTASyk7RVCJ73qrHc7MFF9m3lrsrsPn66XrGQzXLSSkvh8
ltgKWeRZ84Zb/ip0LyxiXhA9JnlrjkiUVb7RPCol1f/zeX5hrmpABOM75gWnFTIyeHMgeEOOwkUH
cGvd4fykurawBMYI5HCRQb/o5mEk0+78tgQIFzp+k9UTxIrnrHGBzwj4Q4VqBe7G/4DTTyvyCIc2
JQpY/XJJLjN4dCB0eztUAs1wpmNbW3BphEx85QIlb5RDuIXncAQ7uZ7qB6JFcSmshIQiYgYNHL4o
90RyaLgUjxerjeTkGUIgSSf/IsKibp/xCr29gu/+1g4tOh6w8YGU0CHpCNnXcdKZbjz3NPo8n5yb
HQwgWjY8r76cEyPIfovqFaevZPw0MpXL3N7rQUR/vrtBFf3pc2Ht/I2Ijj1x4IBHvVOfYRmNXUJK
JsC8n/7JsnD34QXQIvJp3ripiwZ562CNtpg/JYQsqzm4pVJgPplIhTG8+N4xV+gS/ac40brejmm1
gQl/KmRcVMOryRB2rVcnGqcs6SElfvXylNIBMZRpvxeRsztOE7nM3gc/aX/qON3r7jtM015rtiQO
cScNl9HbERYdUKE2Gfw9aDsIcW7DBukB+kSuglIQzkv5IjkCCSxXuK9t5TTIDe4KA71raaTRWMnp
oxd9TyVEOGP5ctKZgRCYPmh8dnvGxgQeOJpBx+L72FuBl6cCYJhap38IWPs878EXl8caX4VHwHJR
m3rUNSJEk4ZbxWwf3AXER+sdoI/dW/R+NNjOgW2fNF5mTRjskSJ8Tw/7892n+LAnM6hu71qyhq1a
sOjlpy4OhdCxbGl66+l27NXwZd6afa5ff6ghC60pc8kUCfgf7SXas7jFpOMzZYnQZWSUttDBDWd7
tjhnak9DCpAC1sz/AyBX5123f0taJbM0EU27Q7Lz9zqWGzBac0BsLnG8YmfN9GzZ0ZZyurnfeBJe
yrq+AXvtU+fdh7zkOvbxEBJigNlzrNbfV/Isd0ZOl3m5ISTYNqadU9wcQT51oQNZkCKr960YpUQ8
NTd2zFWYnmLQ0YhQ4S47vPW2XRvD9kdUzI/bdq9JY7ideQN48153p58yvsTR1sVU6BZ+o59puNUX
XOs1NXWr4eze2ZVJRlRDLWUH05ErIlEeBU+TIDyLru6OHlJHrxNoEHVztLXzrHyEMirfDsCKLv+1
NuSFD3Sq4szhOCxrMpV2Cnrold5aBHV5/TQNkbAsGxvWxoRDsJWRDrw16ewo6g9oUnSEXceyK+xo
HHYa2kE9Nlr2wEZ9hp0hNOU1GUvFtLHhKH8/RcNYSLuphcLK0jnZWJDwsPzF8PglHRm5VTGg09VB
oBI8dutSFE4nINqEa+FBlrsqvVILVeJu1y3jIOYIP6GTUGqPwGDfFfi+AlKsoD2pEEScWigkSlvz
9WpFGDQaYQQsv1KnjY1wC+Ud6LG+LRIM6fT3q3G0uzCjn0B3z7Z6ApCFwunKBcmkptr7W5we0w+c
3S6qXzsuobKVWc/3b14o7PnioTaxJyysEXS8mtW2+I0oYnBfIcvW9jyp3dUcgIMZIpVzDZySyOX5
vtx4hbrYxz4GmvqJINU+jg0zhvYyhcg+GNKauy0cb63RAsR6cYdUcGk6u1N8C7Y+BAPJkCDqG/6e
7Nbvr0bDp1WYApD5+ObFtPfclJbDubsupL0Msrh4Ft1V0Jo1+O3QHZVnJ6OuSkv/L2B8aptyHM32
Fi/vMgWcIqVlN6+Lvtuml4olpVA0AS2oMPTLsHxoQklDG1TWeSbwXqau8e6RXad5TljwLz+wd7a0
OSnbdqfeWLN9we1+sF5A5/k1oQ9j4qbMpD48gHwcTh8R7thvr/q0+7B45wT4gmFPBeYJoiOuU0ot
idgE9xqzCqQvZ1umlJD4R3uKJc6knfH/EBMAzlMyYEYBxnLRZWfA9KgVjwJ/WPv0/o68uY+eMoBN
s7zM8k4R/AW/kp9rifUJM5Vb8WXo4rQu9bWlQ4LfWb7C2rJ4iyCRs/E1T+UWC/FALmpf+CoNYRY3
Jo8VQ66hYwiRxkMSmxCj651E0weXci03DSTIFAB6RMxQn9/G36PAJcCYg7Re1cSvkKrJF5bU4gzw
I/zmGuWXseu3vv7gBr2NtwUmy5Rgo9kccUPwUfHZiUu5sgitVYDII9UkxtetGXElfecg9OJr5dn6
mREgOsl8mSXRVuCjENJdHJZQy3FDPC4Bz6/xGz1VPSFABSIIYjw9cxp0NqL0+7JPo7nLfNPOrYpM
6cQY9AAOltGrfIWLJnPCsp0P5DGKbkAb8ZoQcKpM7bLNCZitaDxEcohrUelPVI+xJUFmZvV9o707
MCH97uqhfl9uRNtzonFhd/TR6b5srCb60g4XTjQYKiLHKigOlVdgFB3mR5nqryLMo1uqzRH25KdU
it9f4fOsZ1QgBeFS/19T93usIQTBbfVQB3yB0dFngl+sFzTZAYXv8uKUn7/IMqikoK066wUbhpEV
SVHI0rmoenHAkyz1QMW3qIb0kGC3svALn/Bnxz33IW5n6hqF2kd9vDSXaEJMkFWGYlJB3+9zZEyG
4MH39d+6r24gfGn7hvm8AhGBJQpWSk60dLUlstKyV0dVc+47/EgCQBlkyHvYrOWJQge5b/Fue65a
nXkpxENCkXO3N0Ru8WKwTmjx4fcvD5X6M6qBCStl0864C7LLqfzU7W0Q05wOQ0bH3fLsDSi4EBG6
EFKrvsSrZbnFy3FCFVDxuBDC2//7RpdL7wF2VUjuDoGXiCKDwe9vYYvQZy7t0eLyW/dfRobXTSIG
zBCNOpNqAdg1CgE/1he+7ao2IZu6cjDSSJjBmyoj67IqJodPaT6T6CDHZZ3INTKDm6O6UCgVXdZq
zJ7Dd4rKh5S08805cgCRvM3TKxYfDpEOTEH7FPXrms34QZnj5hAs23i9UmTUk61WG/kBgY4UMrMu
VkLgvkTTlZ2DEfc9mN70iFMfm3jc2fzFj+0LT3vQN9fOrmJdEBzSJzkQhoRmbwKD7rRKmT348TfP
SJOBW+Hqi5wk2J9WmJqfauBbWRMhnPfJNsFfiY4vIsTisyx2YNpEYMe7n2ER7GQ9RhlN1qfDTf6R
+T6xnjmigIfk2jAo8AoxoVubH2X6Xf/VDH7AGF4eakgkTBm5b7eCRSJNqj1MHjJtOsiDbzsQ2fsu
kwA4FIPf2wG+Vz4htk1AWIF+qNV/LTmtDsanm2uTbIh2BXANQRh0TCKnXPoIcoGk8oC/KcmuE7xn
ZrtAALOiLs+qUkhSZlelQoO0IfSu0sTymqKyWgxTBsDaBkUcr3WUyFuV+oCpCeWTw+1x1sM9CyYZ
7j5Uxz7g4EY2GIU5dbwCz7pZBoEB64+N7CEjHEMvg17r4cGRvpUWXIQyW3TKBY6gyxo42O62JDUy
FMSRGnwNxx5ahOu6YRoIMhLRDYHL0iT/rzFFXlpI9fvyzq5L7LaLwp/yM9KTc/Y9EwwWksqMx4Wn
Nf9+B+18EWPg8Ocs9b/ZoStn/gDK5AHjjPlL0/al3TmAiuh9FtxEoeDSqXHGmCIGO85a6wzJH4vG
snjxbBcQqvgcfIPLqbnPFNWaXuQCwqZb+lfa8JjDekmsu4bpAAjT7ZPCOarYXBxh55mlMSu8ITdh
o9yrgfoQVOkPG5np9h1LXvYp7SyE5MdGOt3M7m0vr+PDWvrLbop8QAAPO2c6jRxugmcvZEjl+IZS
NVFaRKWVAZ8+uGNDUyj36XA/MKbHMc9LxbKRUrkuS8tpAPX2KBJbacwo3Tj1UE3LjZ11sghj624k
CTixw0QhY06LM5DodKwzuhYIMStH+XGpVgj/Kq3+GaIxnyYPE0v7aWmBFcoxX6ggf+7a5krnMIxb
GOSvfjGGh6oW1EuXPQpJm0Mup8h0NfF/utsmhogAM5KCoSoIGmMgG3Gudz+kCk4+6nzmdaJOhPYO
m3AlX2es/eQp8NJKeIjR0j0+coANJ29xm2xAt214z2c+iw1vGstjDm2w6pjtFzn5BdoHUDQb2N4D
o3D3g0g+N9KOPTIDAjYS9RFqrlGun+ewtiQbwgsFLTa9cTul0A3n2rPCxIHwN/P81CzjC8XzVUl1
muF7ktBPWjMVU1eO9FAmKzH1ufSIMkBmEJmgZs6zs02aXpmHfOfS6ebdEM34r+oF5fS67n6RPDrL
+AQL3wfDz72f7jLWfM9sli1XS27vg15vusiEx7+RoDLRJ5ZAZsgp412QV4pj5lvu2LKFBEOpeekg
520E2AGuSycrvrU+9ehatNLqAU8DTosFO6bXUlrMlzn3x95q/s+a4V/TDk1sU3VUC5NBuYugNAFy
3LUSEUVzZVPMJdK8p0ztd8G7mz4GdV7k9F8YZPZxH9ZQ7alfVcCFXqPy8NcL5bFwx1JcAP0CuxDk
i4vOOOJANuYM1luVnKYaDb0b3TZqLY+9kpGcioW5Si5VWETRuIPz2ZZoqNYmy/PbJDnWUc8bESbK
bamPf0MSXTto63/MhXWngO23Dunv1Ng35AEX99rGRf4pkPQkxFWygx4p9CjosuW7BF9Ut+cxVgBZ
WvnYr2kzYyGY7zj7y/vdlpd/iLWuGRdG9W5KA3uX11Tu2BfHf5VhNqUyTNFOXGnyWOT7qoRmcbsv
LRKjxHcIuIRAdjJT7TRjXhYnfAg0glLfnLjuxj0E8YyRDDp3JLlmFfUMwKe6/n0Ef2+Mcm6H2/Cv
9hn/Oweh55RonE2qnXG+EOM1IhuZBtRTtudHJX1/Ggz5dhr0M5ublhYrcz3lyVh0EhM3qCkUuaKb
Y5YhDm8HA1gTXWJr7IODHKLyfoBFv7o5K/e3idCWS75erJuYVGjaWk8x2vjxUIBwm2IlzBHQz91s
i3Wheb8u4XzfAwCZFxxPj19RV4X67t1Q8W6E2I61LC9PHNS8i6bg1KxuIyMD1H/2wXgS3xJvBvZS
5UBhmuBRqGumODnWSFtj8jk+EXLY9VGI6QeldeRiQ+5iu6jriR9cR05FvLhvzqDpc1TA3Pl6FNxA
WVx/AfPxmsFFFMhm8aXcnxL1jNvEfmS/XsIaXqMNVoPM3BrsQThQR4Mjz+k3OQtJfFLEvu23jmTV
vBxPH9Q8Wgj29jUxIoTaDKnul0fDHSjCiMEsW/VFbKPCaPVWrNHZWUe3NAhcUwehxe1krg97zKnI
+fw+m6cs65hke6YekX84xOeZ7PbWjjB7t3TNoqyg79+6Ml1lkMc8D1UL/J22AK1Ao5Ls0Lr5UCpG
ykDuAuODQxUAKM8eRSnDWUgnM4ZDm16pJCMYtN2B/ZW/zM5gxXdE7DIYlMHfUBRZ1xntGBy6sG/M
seB1dcEBX04U+aHMI6kywud7vyGnWfVd/lGSfO+a0TqkXRCcV/thppit/bfYpOunhIQXKeHqwkW4
kDo+4JaY26YB8p2zN6GW9J82kcHD7/z/PF0NbN1ErLciB7tfxh4c73pphDEni3DUEY+k4XQocInb
yXVA3Sx4hnJLE1crF1nUMyUqgGrCwo6GT+AVHJ2EXRhpXjG9VMUnuhnWrepK+byZrEGpQjjQ5Lad
OjyBwUu6xMOUDSEjDVA7fRS5d+p1ljEdBeFs/JlcO3mJ4OnRIc0PbmiNyuUbbWF8I5ohNSRhaLjP
T4zGbJpzLL1bysYpWa7nrtfzTV2Vl/Iw4dc05QbnhLJ4vTrGhAuc9e670PmYl0OsMTBZIZ/guuVr
Xe6UklbuGozBED9Sx5xuC/k6vEkMeb9KTOengLAmh1KikIHDULr2bkD3aY5QvR66f67nnG00z8ss
glB4n1wDbkJtqUXnMif5RP8kVKbQKsYdLSVI0xpKDL/yj7eakRtegjL6Vuv7ErsTCequvdDlSEpf
z4sPbDQXlFYR1bQRFqO8KqL4uZCLvhV615e8tmnPBRMeUW0A8PpXAJvhYSaLnBF69aGxNZI3P9Te
IRfuTwaKD07iN5E9m6rDvlaCRFzo9m5x2HguUYIkTwJLWo9+/EfIFNtixpHlOpAwWwoeWlknFfPZ
uxWFdTLtsQ1+q6Xp0HVha7iF1XDUwShofsKdWvuGvZFjls5AAs//CkxWaEMHCO8rTSi8ilGURBg8
9yXJJn7rUMW5cObp31kE1J5+3e205okBxRwyIluONfQv1rE1MjtWs+N8jZRLo9PoDLiP7JzK43cP
rMSrN6aJR1uEd1QK6XU2BDJyN9IRU1lDB06JWWOQOindR+o4ZgRgpRFho03CSScZrbJ7pDyGjjH9
MkPpIF2Z/aw2D/lboeOLBzQnAsADPVNSkYq+v5N2IJLQSG6uTqnB5QbvamzwXLhLBJn/kws/4JMp
gUVooxL50pVk0M7UXds+HsGeZCgQ+oBKPDWcw7wIpIsltBiOkH/G0KF0y/Mv1ntz3KiwErtd4HRq
b5vaQPjVCeTKhqpKZoLGJKv/NxPS/Dg4j4LRMmKrDm8EBv9ruzJLhlx8EsEOWKSXgyV0fxX9yAnk
oWNt/2q1I6vHvoS/aMSr7Ak3in0s717ZEGAKX9TPlrL/Cjz8Dusyo8B+Camcy+lYi6AewR0w6PV1
ZDEm5Vk5woNXctyOUohbunDNUsa/CQsdpH2efRfk/V2KTIGjBW+qE64CVlVWiRwr7I3DucQIiOCi
QMHC9oXJbXey7/AlqTO2l4DFzh87iwCsMYSgYjSZOAPyIAePRZIZV/YQJXhws6wUIVwQyUCPFej6
VMKz5b+jzYcLdY2UH1TT6pZzyH/fNWNjhp/wH4JIm6Hzdw+dYKYNa4KvY09s0kHvz2X5R/bD4qxD
/5ZO1Z9tw/2q/Hjw4sqYHRWNgBNTRlXVdsyxT8ZMz8CZNQOGSmFyoF7f+OFA4XC24wcDB1zV8lbO
MGjmEqZmvcXX8uhgHk89fSN/gLw+Y3nssZa+DEaaO5qdWpImGMWgJByUPkPIFNrMqesosWwmDCDD
VZb36I4edh9lriGG9zimXJJ9tNdngp9Ll2x05bJnE+FSkjU0F9qY87HCcwhqhdnmPPrlg8/j6XL/
behABitA1BdIXitrwei8dxiY4sIo3wnJR6gST/xTUtBD0kh0wisAg7eFovkJNYkHlOVqUY7ko4sv
8ElxlBUzMGgty9EPdCXP1uAhndT29KRD0D7p9BAsJxLYr9hC5+cm3FuC2UJZCviDuxl3uAc9/R9g
PU0EsVh05bPMUI63NzLlGY/CxWVogBX2/YI8gCA9wu2wKyRas6jltpXe2IrubgaquqYfhEl67l9p
zcfTp1xBpERpRS2f1DJWJOV7NafrhLWGLeR/AG9ECf5x7jD0ouqwhJY4eCD49QSIeMifNKw2ngcZ
oQwM9fofBOUZuLW4OL6UiZBtz3BA4bDx5yY4u+LmWGTJ7CfPY4taxFdmN0dv/0DqKXMbDHKzZNjr
66S/xEa89rLkVLop7P00VQloMN6+w5e/Z27RmuwgR3wM9nr4oh0voE4FNeSajyD7MLDNl/YPefhV
14WLgtrV2tMiEmiR3lfxb/9Z5c5rCZlf5yhyAAtoQ8XlD+aG0bbb5i1zQINHdVnbMxbUqx67Mise
jdIropeuLPNqHzRsfvLolNVLuQpWwxa/sEUeIROBriKqNbSXSLyjRXG9cb0UUodCqiCGi3F/NQnp
yFHdW/XBp0oc184UoS0ciW7/58sh8sHzO+DMEv7tCpXTN0Xv3HEixa3AORS40a4qqK2NsVj6UxFR
QwozMZwI1/7O4wpPd2X/N/zc4JH0rrSxmPhSf6DBYTYOZbfAqoErwcjKpsTdYu8UFxHX+ed7SHIp
cpiCgjMMEs/+mxJ2SavHac3G97tMixeVFZ1IckjpaP0K92v7e7FdWmEREue6TB+a/1Rcv0xoTvO6
G0UYNHWXXSchynNyiSGRAynbIC9JUK7a5oELXIeg/ILk+JOod/sKBfHxRTtM3wxrPj3xNpikQqa5
xYkYB4EQ6ZRAt82/dcw1I9wdbbchSMtB4ZlTOWEXPxKonkvcPgMoLBDPu/xlZkn9AcsJKnaES88Q
nUcDKbcQUeFjTutU+gcvWCZZHny5y+uyi66f7Gm0ADghraXn5i1SC/yNSsZ2GwrPnKms0qVjKG7B
vM5bo+9TF1GctWkqXczCwSvrFNnybjtzXVfdtSsqgs9IEBpNpKtQOkzJ7dOGsTVDcUvxmxcJom3Y
Ekfx3iVmTECsLJpHLWzofwBdC3LouDLV/xptNlHADjXjbOv4/efZ5VC0MsggCFyZUb7b3bEv4Obl
iYgSs80klGVBcvvZ2UIiDLDPgAfJO3NZsPA90ecicfSK+UYkNjafZsBAX3NR10kfQQ+86z6XXsJp
N62TdiLYBNCIBIobpC3OGHr/RRkebvJ3SEyCtrQPxVYgEstTBXk9NZe5qE7t4KpNx0s3B58yodEp
LhnDU9zfpMMKvqxHBlGOCKuS1ql7m0/qQ08RjWjv2xMW7w9OzF040vbb41LCIdDfa14mtCkDm1f2
E68Yxl4mJxZ+Pc0cqGq2xBLBkl5/oZJan5/0WuZamSRJLrzGLTClLaoWxyI0hSB8Qhg4SW/AV9v+
73LGh8cLSjBV17MOwzNlLuhEF2iPS4l8x5ZMP5K+wO/5OaKQDctkfOUwxh9OUuKdGkTxBaLM0W7j
ILjOxGdr74F1xqcPTbcgLGJumOsyMEHTFQfdpm1ccY/Hotm7+GxAZ0RgGg2Cvik4F5gG3KI8yzEi
Jc3hze03duo29S/RkHaa3b28uxx+EEDNXtkH67NMb7oW3hUfWnQZGj9jEOeqofX3c+Dqve/oW9aN
Lc+FWSuFlSo612xsOJiDS/Sgf6Bkmxa/okwa1lb5e8ZWvwyX3wy+sI+e/z+7J1MzcRwkxALXseKN
NJEpX4TNb9LBZ+RZMtwp+HlZy0EeESu46xMWoRt91RXB6S1xFZAu+9kuHB5Nf6p+T0u/Ngvx5pe6
Z4+/ISQ/aPzqXyJSRMBPnsVMQyUDFg8A6jdPGT04oi/nyKNexjWdJVo2X93wD50P4E9OD8TR3tA7
0Ftt495oS0AlaUGsBjx2qa1g4W+mS4mzpUMJXDZmZyzv8fij1TtcK1YctsZIlWQKmmN283XQr94H
qfNV8WrCoSuAiPbQ4YY3MRwelosFSHmR4kfyiamfCNxy6wh0yeJX3TsxpCWqLH4jsDX3wbyneRtq
l9LdcDD8ntBlvsNwl52yecOOtIw2pUbqAhP5I82KKD2VIebY3pxLvtdt/pSdSSmwr3cEcpUMU9PN
zrJP9cEyUKLPEuj/AC7wJda2Syg2Y3Ha+qVj6QhNXj+UqjOQYmn9AD5JSQ78R9YU+shT6CcYkkIJ
TJR4EEDAScgBhjs/eDnDRxvZ8UnAZrRshp+z0929I/xtsG9aZObx3ot0pD4kXwDbZQOUs4Fp5t/n
P/fz88JyuHZm2b1O0N37L7uOXrjDjQ4FCI3Linjjyht6oRZlRRSkGGjypcLwa1HUPdzyLqPb+9/8
sF9oJY/ic058hzDv943begFKpnanLWdk2fZyZMVWbGQdx13TnxhRrliMpa4mFJvQU68xDDqQAjXp
4c5Y56PZlhuIu1kNBcXRC0RmTBHOAIIrliQzQh8K+pf0esk1e3WNZLejOSnVL8B0D5KHfTt4Nc/1
ez6vGDwpjwWrfx4NVUHtEg44gOFs6WhO4CDkdOg06z02DKHkxk0Le84QHwHjYpA7AEl9cFPukL2b
O2sHSSvXD7l/qu7sgI6hTW5zUDDry/J8tj0n7yl4Fchpnj/fnurL6DsQ7JpMn4IblGBssVLAHyX7
RYodvjdZqU4Cr7FZ3Lxn0XvEpkN1KkQ2zuNfn5pBqpCkpp8x3LpS2T9nFTlGXRZxFTpz4Vk4kmXu
tVfL5/MWZDE0V8Vnq6X2+ml/B0TlComaAmXXByHlmIT7tEozCbs2FkYJpopGc1xC7opJo4JsaSez
9Ywlv6VVDWdHedqLc49UJz02ckmUV3tNMPDZ+37QSzVF/Ekdc1KKAnTUMjLKUUfrOxJHn0v+mMR7
ghC3IRBWZ/fes/j6ep0QB8CZ5rwdku54AmM/nsQOO4K3rfyPGHeZ/rBt2BQgCOhsrf+Xt61QtTZd
wLu6kJMsNY0y3vSzO/XtwCZzLFC2K7ndOWFU5qpLnUe0NHnveK2IyIXtk7OJ6eQ8GMbnl63ZIxFY
qL0F9jaVFXqpktbws3Eg3qen7cyaT1qF78t619KI2PupWhjhK57TqW65wHI48FfpRm9XAYYkvU6K
Iv2xUQKWKtgsDLXNDSpo2nPM7K7UtyC2sr+yJe4v3xCoKI3pQyW/Nfm14GWDwqZJNgo8Skqz8TE5
j9lyJGhZkI/PllGtOqAJl8mdQONnRGBqTcsrvrt5ECHAx5BTvdm+as1VL8gJTY4k8054sFASlNYD
wygb4CKzxb+SLMhHcEfLijguWmCn0uIQLPZdndluffgXjIiP82qryLN0Bl0HRyJvQ9vwkFNpUEUK
bCfKizAYYnEfSOU89S2YdKV38ihKDN9uynWAZGGzB3vf1tNyQqtjm6EyxxdR300v+dcIB5ME5OP1
V/P1BFn5EL43yh9YjTtoBZpLemhsIBBGyvxiQtyjX3JHiEqN5c8FYFzdfkQTbDkTkVnPHGvA2j9l
8Li9TdxqiS+GNXEgs3E7tKc15PCiMi8h1+y+oroKJNhPSMvRl/mGLzHXca8YHe82U5BbMFO/Tpoh
dxT3969pLGoTeYexcLDU2SaUsH6T5StOEpItghQx0ksEKlxsYJoBTWfFMzl8MrNaoYZ20A9btYo9
baJo+PedcmzWCMTVLHRFruHau+iXrex1tXiM6VajQBIt8SiQnNiBPCRvBJ+Ft3UmNI1wdbsm80df
0pErtbO9S4lyJLMnm/jqXfwWIuPZOCQCvJNdTCW9hcZ1yfsOZW3qDrO6kUY0u5rqDtGbu66hxmtU
ZmSULtQpVHZ77eKuH3FqRWC4i9c5+REJQzJ/DdWIDdjRBXn5C7HEL054yw565dDa+2yvb8/mpMv0
LAPQsDyMunUCMtbxy7MyLPSr6pUojI9++Y++/75edZyjSMdIVw3LNBCjc4lzhJzibX/euji6d62E
sywzGRlddij15AA4hyCAmD3LvKKyo6FQ33Wq9fwh2DDSIAtTeDEbpHMLf6wmMPOGfNEvTNkHXD1D
fW+AVNxv4v1X130yTV6HBz6AEqYVeDnkSOIHAJT+3AsWzYui8mm1+5Zsk/pekrkzFVmFgmWMjrL9
HwJ+la/N3lsketheJNh59dnQ2QjVsjnkms2gaByv4dvS35mziE8d3UTk70JHfCp5ml4+6qjVReqU
nge7WCabvPVHrFhGKSFly+ooiARabgmavFPPWkEpbCbRIycvlh9VoF9/N9jXrckpXzgZBsqlC+Ap
00j2zop0fVdFxdvjGeBypPYAsE6YuJYlEjm4b2SgjJAA0M6JllJwPpsbpNDpJI+4dMUsFL5N6MRh
j5zapgexNjKDwHDCTeJmt2Al7SZ6F/HzX5y9jHupqCXdQVaOLqbNvD+mf3GYAHz67D64paN86cWm
jLQzywubx1fyS2hVJ57cZVzVlubvHTKQKj+2y1u+AVRyEtXaQhYCNIMrHMo470nuxJIWFwT13/Gy
Lj/5SS3dfG9yPgmc7l4AFmYfp1/IzitBNXEwFQhj/IF5NNEEGmSxgRVRTmAZXzrU8fsFu5qSl1ip
jxxZ7JQITuXTFp3TIMhjKXJeb1TvF4AVkpSKDwQu2wmww3Q+tTzsnY2V4pRDPoTwm4MIVwp/zCt2
NrDmBby3nFQ3lt/Ohja1EsKmRI0b5KuWDjolkthtt09CROOz6KL+Hxo5J2od9VcrfnycOsa8VLXR
5rdGA/W+/e85hp7vYFGkED3R5oDHYPJrevNLuQy0xoqIZwIHyoDiwHQABDD0Gr6y5d4z9fLlH3j8
EuA+9Lda8KKSts5DVnXYAm2VrnL+XCarKMziVpgL9HCdW4w/NLHoTCtugJrZG3CbbSOkttla4smr
UCzDuHJvuBpJ3ktMVPCTBEQ1ERk4nnD/rJqO2aMTPRFfPjyw5H7gF7IGnzTJcCBhjAJPQDOHxC8g
7dXsmxf2W2661IKWTaDl+tcESuJQsfig/wILqyaKYVCV2D8MYBplGzCj5+O5+zDwNt5M3WiwqxiK
O8xEPAWy7U4runbKYX3PWcHcA1sjrHAbFfCEGu1/13R30CrBOe7e8O68kavH6+90jzP9trHoCMtB
W2AIbuY3DX0w5u6mtvZ4DZASUvNNTSRuO5aX7/zaodeJ8F32JIEccZqGpmzpbmUTPNhsgtUMIo0A
CaUKg940AtT2/a7A3XUJC6EPh8Ry0t8chMgpN0du/V1aqpu7lUJ6dZPjllQyfFfC6RkDOIC7RYx9
35TjQpilDxGCnVuDANIxa0RbGPz2n89g6VZwgbcSC+4ZLqM26sjHECC980TxvnU339Yd7HyD03CN
fgqkG9acppty0KUUG6Jtl/5Mzvo1OSegHkYKZvytzzj2lIyqXk+Iz/Qjjrc/q9umZjAs+XuKhWiC
0aGKyOxQFDTf7A+0mnIl7wowMnH16vmjaydZX+gFoqcfrAe9NviJb6iTT6cAGAA3OUSTkZG7HPJz
gitqfstfpDUzcpNUmEAGweEHhEeXIM2UzqUQlJ4Sr9X7ctObQOkLYJK1+CNgr7nXDLxdw2uroo+v
FWb0EQ6VxFbJRSofH4nOMIoABMMNImThvtpYdenUFZrGFDA4zHkzTAk7kUif6gHIB/c3YWRSVMbZ
KvZBIsKRzKYFOJYrtj8NntnOEVg1F+cacu/+aFl2JzP0HdibWr61u6RriX+J/C2iwn/PBAG+mW74
uiLhAYtfRisQAenQUHqG30M19xbhhUXrJ+5RY6Ae3B2DYAwlf7y6DF2lAS28jiL4URHYGydYSFvx
zZEBXXzCLZY2g8ttFd4JvFJTrYvL2cG3Ws8k3rBqe8YVJ4fst/s3kovHhjqI/O4s60L91xxh28hB
Banjj7qX8ljJBsXnI9i+eI8jqf3Skwv88S6ucBVA1yGuVXOM8+w/uhTTZF5A8mEMPh36LfDo/vN+
74XtpWVJO7iYHndVbXOwGHqjr5s4V3iZnipiV/hGzeCJllR5MelmLSBb1mUWyKWgnO5+RrxkvBAi
uDR1MvKz663UsjQTW5g2dY1fde6NVZdg828jn13Byf/b8gAcfJxFflO/8hLkImQGfnSGaNvt7+vV
dXufpocrwFx+BxNkuPSTkktQuYICEj+JE0jOy7zLiiEkTPX35OvxvXBtxvA9P2nfoLUBre0J3FgC
qrIA10gFnJeui545yg6edvQTgDMw73sy+aTGUyAWFuWIGPU4JSTAWRlPLMmFjG+Y3DCPcEdmpyaN
C7rzUvagRGmKd7PZKOEYa44CovU4qvelfGql/voUEGflofbLIjCXMHpfRnPRjQamRofefbDmYZKM
Bwr87umqyl0ibitRjoW/RQkHTLNrfwqMpC3uS3q0ZXbsMiI5k2ZwV2OFerYBRaPNnnWNQhfAIrVF
p01RmzvhZH2miaaXxZtj9DYAzPxzo/W/om2gNvAGeStsviA5NFCK4LQemvTObf8xiI1Bf3tzA8a4
Sro6Enj/kFVYV1W38WFGuKyFY6ZYWrAVdnVudujF/gde76JydeSPKZcQFXdlLJwqbIM+aCbv2hGF
rQSfhRMrRP/RjP9wPqp2Rwge+1A8VofnFcEqdCmYhNltYXbJfSItcecHnvDu2mvaOwC0urCo1DtF
jaVVMRuAuNqOm7BnTlzM8LtLQAaG6+1dLfUccmGMaa+nuRLJ/KbBczG5hVOUsgUDTD1WlTFMQQq/
FGJPWMy00G3fxXqFXQLqMo0dhucJfrZ7kxPMW5U0+CP/KOTSzYumpkgW+1f3X75STNBJYhC/HmLL
5z8HUeKJus82Kkc6TfMfwxvb9LXxphtaR4Y7v/Fw/0yUFo0ewnXLP5T4ZY7LkxeErVK+jV83ypXP
EY8DhijBrpcezhdXBz/pbmj4p7fYdP9jc7xMKa93Uk6dvMcMTkb9hQKnjKoVUD/CK6glUVj4VTKs
mNy/jaiHKrbrWu9uFs50HzN4UAmj2TkNlW5iv4ChL7OiYNWC5MkG7Q6VxMx1Njf6BAnnWkSRzFkD
WtloK3zVPb3fVuUUexhAM2kI2xvIikVULMtM35e5I8i9K+QQ6V2jQF342KWzK203kqNOvbzfmwf3
DBsX1Hbs2++PRN6lHHWnrw7Dcnxq/q75Y1exT3VEoarM7VRUTfPzIaSUK2C1LQGfrMh+2CiHT6R3
U3qUcVpOsNWj5FvcnU3xxezVHVpJuEsSi/3vlY5/+rNqoPRJdyuwQefsxaRtt+bDg/38jvUA2paM
gVLRo3KOdKUuCIaXYWps9js1Kce9mMSDDyENoMA5jL+f/8B+vHg0lgkLOxVkAb8Q/KgKTlv0cldH
BquozYSxciZrQaJl4/ckOQITilJBtKUQAS3xyZRTs0BgL8ddoOmUlXGtql6bcH/PDjZSEdshYWgC
U3B3JoV2kSRFqmyqaMIs+b5osCCXp7yKCgYICH/8LuARpU0F4VBGOGD7YxWQ2D1d3YCDQfuh3mgG
gxwoesOC+nW612bTS7iGWk49leXW9Mb9FOgN09jbj3UvP+O2dL/dqQUDu++NelRw53+zXcc6PzJu
apEqKLzPJ477/sYvu3T7eyUFIEiIvb3B4T1hoaA2mWfxdRbXI8S3ibFSE75AkoEKhfi2BCxJxaE+
AfXLfXnz8R13uoJQkDE0JQPPEaCwYRORyf6PRouPg2QCFINbjjZKWelLTELCEfqkHsY6QEyPudDK
t7T1VH6JxJVeLT976ysUmcnUXO2WGAqdUon78D09wtLS0cVuo7+yS/14vIvjIjgyHwMXwy+LROC8
pPpobccfwvWjrreoRVj0/xVl0+j6lKVPBk5YehYV6agxlJTy7CnVaRffJuyEyfOdIUc4PfeZRftV
kpzdx6//3lWZilRQcyNFYJ4EU8yjEJxqCoGV/dqaF6oJyXR33OxhM7LHQzJeTBgA99DHe3Bs/hKG
SARBHH5hmqBW+sdWG2nrdqBS7+RJ8/T4HRkx2Gnl//iLm/QTdCx1dSCZ5is6EWeFab/YOWbMH7SG
cil/Ka6RpKIMF9kfVbcsoqSPMsvVezdyxukqnUzx+AmRMqaZrVqBdZ8dKflBwg6zv9oftFbBctYK
rlHmvQ/OFlCVVjzD5DD4HA1l6mPmtnfNGf5f6WkmKjeD6DAGzTJYGejcdBgSLbZyt1HZ1I1JzgR/
sd63NBMBaDRknfAfylyqXHXf32UqgYGuBMD/xkObDvAb9NB432Px9+F0RyQasWTGhAZNdlM8ciN8
O2HSghkPRUjHp/bQSClzO25HLG97gi9pGTMawgdisxFA72hBGD6/idAKBrrwMnrocSgyNGbJ8z26
vTKgvbLjDarmhvkePI65oQvCCbEfB5SFrflRRrr9qAsFaYbSyNQw8LnbXKVfgFk0n2xfFnY5Kmw3
REf7yUig6NWQe+lwkXgNIDxB0inwSexxc0ewOI5SmlF4W61M6TC1GFjYhbqgxuZfD0I5SYbW+neA
7DiwQBdQWloICcLGHu8MCfM+JnFAeFN5nQVOkdp7DCgSe+eLDuDzcnaNylZsd4pQSaHdXBPdyUJJ
oG6n53VdkNl37L6T7fUYWHDaYnJUbdXwgsmT38zwzCBuGlwcPelGifcjzJJh30KGDuMvDwx4cooM
y0R9Tb66lmQgJTrJT2EQTiaHMBBxdNPpDEKSwVL8YVJvdl8QrQeyO7VwdpHFuMHIyqt+ui83rRgp
xfA4aXH1u/T4GwiK0yAXPgKasiy71gSsH3aVtqFG6boOyKaxo8IIbCxulVdajBUd78qzCUmfNtkh
J5bpUUN10RgsRb0cHeWDnn0XsMateVSTgpW7W52ni11nqNfkpj/VJo3zmzArv66WoypCkC7OWWPB
z9Jlp/cM4WJSBLhCThDDtLcnDZ+FCjQChZfxEr7Yp0YagQRPNrcSAQvv6lj4PBZI+WvZ4Sm23n55
lrXQshSMXgUpJIEBH/ScmKrvumd45i7aL8IICflZz33fKUQ1GpYsw6xGQmbKPVKvy3OJf2lKR3Rl
yRRcrnTi3/Q1440S2mlgUleTj9L1FdR9EFFUuUdl/1yI0FH242SlJ+Xlbhjdcjqa9GNmrLtnsdA1
mBjo3I8I1aMNY7zl3hoEZVHa7kMOrmWeAaV/6G2REN5C0p4lE6bf4IyzCa4SczL5JLqtlYyaYwkS
F0HSP3ZhK1K1S97ZCoXsT5C9LGChq03fijaAMKaBU5V4uDzEDVhMmQl9G0/VB794bTeN14OoUWJ0
Qbx+Saewzm20YcPdTn/L+fl5XBLiBwn/muG7XphenQAX8NcTCI7EoEJiG9ZtchxyNU4hT9NjFpK6
KVGW897ZwCIdONlHohxnMF0CZwWZ+ZtOHhHZsAOWTCbBCORtB3X0jDTd2UDud/D88dc8HbRPqPXD
Mrob/Hg/phGgPIsVC7C6ANC9xuBW7qov8tP9+lxYR6CQsXjrVIQ5IVZWQuEyShR1PwpaRQ7GGGhm
W7oJ+gPRJxdpSb/wq36Q3fMcJaxoLhXkxAOUtBsRBJx7JM4LiEhWhcT+ZoUOnDyr7OywHlSjORUG
tbaMGxc7DzC13F19T8XHzv4vVsuQvHKH2aWWugHj77ahXS8RHymp4VTKCP3z5KJH3U8WkC2SgQC+
siyRt9CoDAUQtXOhnE8fUQsQaw7Z5wuQJvJRnImb6YZB93OBtcb3vqVUSNAwmMnqExCq1n7DTUDY
dyb25kzbPgoJe3av1Do47qS4+i0lZdDLByZmKTgnFWEHvrZbS68jkYjWnD6m9pzaNwRVer7XOXOA
k8gBz4isCHVayhIZjNtbERuNxIsZhdda6YIJIuQwls2Dha5g4cf79Gkxxlsfp4GcDIjhbsxosdps
OvCUna6fZoMrpmg5gZVl3KKyXzBJQf5Vq9DNITmFlkepIHvYt6qp8SfjlufpeVhl5sQdAXQQO8kd
N3aBzWrAOlWbTPVulRlH55mxz9344XiuFwTwgVpiuqghvU9CYqE4TE+mDw0KNjZ/IVyTrFmpmAlm
bBVwLqBYACX3lns9KbZEiMUgcoR8WVyEQiSAB2rVjBL5ZVWqHZA63gh8NEG2WILSEL0QbhTSukaw
7YkgeyfLbJuFj2u3fYubj8ERMqjyYGSyY8QmH9edZOlfdVfPZY9PSjmvjKmGapJ7syyZ3riYNebG
DVnYeqWJ6gJkDd87K6tRNSA9EOyKvW/6IPE9uhRTSzvkuHtcSHiH78kqv07OFwX9f0mA8K9SGiVv
fa0migS7SYQ4dAMWied65+LvBtV+P0Zg0FFV7QUkUFcBuOXeYTE7DVqp51z6QMivpDSJZObmLfl8
UnCpoJRrHDXLmlKOa1eE6y0YBVGxuucKgo9VRQz7qEOC7Cc0HGINdqjr1IuIzM0TX6KvYDSfM6JH
Ll51QGsJxOxEOUfs2OrTKPrKdyY2VU5y2BwbUlypTuEfvIw+UjiZv/iXx/kCKGAPddwxa6QUiOSk
jPe/SiJNVYeJ4K+z1V+T61YqkyBU9HrcKTPSOprORo1fUm6wyEF5cjnSkPOFhtrC8rEhnZR7mFIi
7l8f1097nfmz5R/g5AFf7sK/1d5n0+CGH7igc1VUxHMk5sSf/vXvTVuisNF2Fa4IFbafIpyPTUds
DDrLqf/O8/2tZS+EYrKuxPPuNyVAIJv+lbjx0CRwKpen8Ce8AKVxIpZuDY/0BwaU3D4htuQP6piL
z+I6GI938/Oiq11NUMTVI1oLGzQLB7WoaCxydCT10L34Ci/5vuyVwogjpTjhP14BjHSO04ow0IC0
mxp4dEyJE7YsaHe1iF8kI6y2jxc/3P8StqrJLtArjMZNOFzMtCVdcG7Cg5pEEtbkuRByDIjd/WVh
/B6X36JLhAdkEVPapbzwbUEvqF89d63SN868SsmiMkzHf/wDiHfki9i1xy0/nYUdHV/rAMJ91dbK
sHeq/JZGNQBuzpg4I1jLcp9O4m0CrhWs2CUXQiAz3aCcTRW+CfSefXpzNYkbEiPuGYVuBpNwxImL
fHYAidVHyNOeQ1ICekrleJhozmYN1TbU5B+zVu63LITSrDis0GO7flAZABRyqxEue77vHXi0TQcu
rreGVBjtwxw3aKBsKaaH4EovqSHCgvjGqL2S9UMHdTP9sJk9EN1bcTDG3VBDO15LZVdeOOKBFP9F
OonozS6bB+AM6cp8NAPml4JnFq+iKiFwLST9F+f5ywpzhfuOAALiEfjnee7tlLGN9bL9i+WA4Iqx
6FmHr0JDPc/1K64ZFcR1aWGwmer5EZJbpVJ4ueixrPfRHm4uWia46adfH6JDX87u7JWTWJTFCP/r
x/4Sp1brQ35M2LSDiqj9+NUDT3uzohCZ1kZiFF106XHONH3RNbs4QG2RMF1+Au9lDN9pyq4ATS7O
Fq1IPCYAGYphRVDfU12s9KWOWxDCpiSt13CgRQcb9vnr/8cC1PO/LhDPuu59es7LZK+HJ116DZWe
Vn1BWn/+RLa+4ZeaBqYGzQZs2bjs1h7ky8qfa4sF1sbyac3Otv87fXJ0l+ZNyblJ5AvE/G96G2I6
fzNyUFeZGPv+OBbkdkLd44tDFt9fPvWJFSR5sVmgjyuwmx1Fqz+zHy7wgNlJyrrJ0qvG54Yy4zm1
J1PvhntFi5DIMgzgHnxmYzGCL20c4JMsqr/w6/U7iMIjga5t/uiNwdN6a5Yi2e36s9oK5seaiRlF
tGNye3lbSrsUFjppVJVOpJXHSVPGtlpDhXbdyR0Mvyq/QungmQqdY5E5Qruq4YjPRh5v/nbuQ3xW
bkK5lnU/Z/q0gkATNmJSEB+fZFiddWs4wRjbG/ymwOsFBpfOY11B8P4OMqaXMsqtG4AaQPpYv0jl
1Qi9pvrdQ3AQxOzNjzJwtACbTg7AKOHuJJbZdTdnjAbsSLqrPvMtMEO+LGvZuXv2+ZwpzjES2mLQ
mMssVTjOfHBPgMJNxIewt1sDZJY1VmxaH7jGZdgmSrXmqecb949Rvb5gsCrk0OrwVyzp1h9tzyC0
kViQkxaEPHtMLJXwwoAW408dwuhHKGT7xlo+ocas5ORANCYM5uz+cZwI6VwxwMfu9SkJcxg3iR8l
yb1Nkxm+LBik5td1n1pKa2/k4E14ZAKe5L1Sc415xCekTgYtV34pHxE0MJSD8y0BWrEKRgJx7jML
GqKbHOR2tYYSQO4MCpXmbJ5MfPCum4CGOUbgjj2lmDyhuY0JCUWFrhO7h4b6VFDvhZJ57PTUjiVQ
vTE9AH73/Cp9ItuZ871y1/UGC9QO5jQ6XJxgCswlnTjzQOADZ+5BB4UshFtoe7zwWNz6If7N+MrL
aTr+im65At///PP1BCNQssHP13GLE5C/yrpCrjBt/SdxFCDG9mC6QUDD6NG8PL82yLoBDl0kt3pA
jXq0mJNmdF3W6asDTTP3JnymGD7qBAoV5MNSUUzMkqegA8d9Dgok5w8OrjaIu0bxsn9P+//C6UF4
VobBs3hsTlLv3c17bzRq/JjbUw3pZFFzZ6GLT0Htv00nd6QfVYcEKjm96MlFBjifcmQaqTP/gz6S
8dYs9jKPw3LmiUljHb3ZYV+JwvoKTljb6XIoe4+KnyXTUYoBqRx7w7MoYp4n6uiuJ52w5TTrw2RK
QNUXBwp8hQAjthOFxU9O52ZuAn5PM8aqOKxbbjhC97LGidtnkDLuaUPtwonVgeaxJEb+zwPxkbJV
OGUMFAyC66JS64KTUHDWLDB/OV4EnP1ahSf/riw/xfu9k4P4Z4hJf1hYrQMbsAGmmfRxgWh63SAH
4t8HdeAWOAKcbB2z9KRcoyRB5V1djCmRt5VHgihBj8XXzBNS1FCzl8T5/kiJcoKmCmDwAt6Fa2Do
xeg1lGZ7UzHrXv4hlFm0B9fopp51EglL8mMHw89SFTgTyKIPrXn/E0Mua0GQTYnxE/qTQOky30V2
T9LoOV8ik++BgkAKA9M2ismxcQYBrhE0XmbpZ9zdw4Icof5OoK0XKLsbhLtqfnr4P9XGVSEVxeiu
+O+Jy9vpaUMjODxLDntQGCuWNJ7NM2+sT43hTHrIiPPh8SGl2Yo394TxtNPOdxh3Y7iXsKEc1AVM
s53a7/AwVPKwacNi4YQVZS8ABTqxtHNUbq6LiSECSGRYgxkQ+t7g3lsqoZ9d9BMDLORboTry5NFf
4G+CNhcpjyh1eMs8sKvaALoxzbFPaN6lTnjn6TLj0NE0Ve/zYmwTh70cWFm5Vpj8iveJcS47CBc8
V/JksY7ZbBEFT++dYcCcp+blaXNXX4Zpn8kKLEcSZ6r9vAXKXTntUClggBxuFNPjgsQzTWTp40/K
MuxJM1wYoJNfxEYVkdJ24rkNOviHOzzefxjId9zQJTd2BoY6o9DK8j9MOQ1N24C2WXgqzL4+z6He
dloQpkKO26I/FCrLy9XGHp2b9WCyexXhzTCHBL1whtIGYzcxP8uU/zlDBxi6MX1V8fAeA7Zl9UGp
ciNhKlVYxsxfHT5QK4k23xzWuOJ2GI9tBQWvTrNc4MdgWt2QDwi14Ht7QntUzOi7iq7m0kfFtFsZ
Dgct+HN8H24tTeOPOfWZRmNvL6tHByQRgpC4kBMmp/j4C8/rp0ca1y7PaE9Ylp81kRvqNcIXqMSK
u03QS2kVdMC0kLnykKuqcCINU9d5v05PEv+4TBhyy7cYHNzo/yso6c3pgd7XCMZL7MxqfMF5tfJh
udWBbLIrn6fn1MWPMUj97lIajM1h2v/ayLfSn1mvXwCZheCFfPZw1ypKYkoz0EAELebcKsqHPKUg
TzqFHFkU9ByvtajnUk4St7MpjtfnmRDVDtoFMost79m4r1vwwe1o2W6E4trmEVjb3VSuZ83CBm60
ETQvUdwH49qUEE6eORnP/w9MY7J+wbBJkI44URDbsOTP9Qm+s6qyHdeVPk1znMpVcHSa6yEsCae3
VOC0QNvL3FvoORI23gysDdI5f+wFtKBjqoIzgHW/bgWM/lRzZEzpOtatT4jnTR/rJRfJrQaI2055
KJp8uK5zkLTuinOg0a09tYCxXs2eMuNzDD65BY90NRSvg6cv0Pcuk6+7uvFEbiNFwkE/Nj5eaChz
IYhJBWPIRolRfNbNcvH+YFtcjfwwffgiozdFUBiT62HX4VDMDAG+WurhvGJOA9gWQw4yIhH4gIm1
dFLM11keKQEydDBlTIukZrIrmysnctJWQ2mAKh1PjD0StuWd30zz4S3R6sn4sl7KFUbbx9aaCk9o
hwwiqsdbTDQcjhQmXaoRZlgsANLzYbcUWZRnliL5dR3hKwsHj0f6RAf/vqFhSaFYUJDz0FZ3dF8w
aslJqtj1qy4MHXy/Px5MVXDxm6HwBIeissVeN9kbGaNXkspMURk19MZsc1B2XS6OfVAKLf6QPSI9
Tg+CEdjd035p4sngUwT7xj9q9VOx6hNhUN4j86uCIsClWfeen+k+c2Degfb3sXpVNa8ZHKedbq4h
cN17GwPQNa5sQxxn0FCUPrFlwPciEQhSZFqwbe1WT1goNYkRImOyxCqW0HmnTpQ/NYmAt4kSzj9h
SNeWAV6METlqHHWz17ZPMdqL813arC0XsOHCupz42AeldUjqm3eZOUMqNoFp7p78dYm0HN3/Gwkb
d5B5Q+/T3pVFiUg1j+kaYMEuImfnXiJkz5kRDaFt9zPoZFM67Rjh8UFfYvOdVhpBgh1t2V6mEef2
HdX0ZCinAO2aruqcun0RaWzA8yF4+nDb8r0ENHhNPJm4sFfEnv2aUBtQRLDb71QpJ/TH0lCa8tyx
cmBfKQzfMy691VkLDzlYxZPX9YqeuxfkH6ZJk1nJqCGRFqWuPtu4UfHpn2i+JLOrGOUUCuOGTier
G65OzXfnQRTXJizJ2wVbhvngcDzdpe9tnMgn402pi0CcWl27ots4k6xVciBKWD7PpKicGvvnpmnC
goMWsI6OQBzARNpQRBkNCPmkT2t6VhpVbV4o3toSK+/9MK2xnWMSnFj8pkCZt/LmQ8BezYWG8fM5
Nu7bJpVUCbae14Yu9xjRLo5JBIY0lkmVpKV9DP7jPAXIFCZ8A/MzChGd0XGEMM+Mk5LdJUoTWof4
7+uDYNLsrFJyabjY+T3WlCqRO2wWh6LJDRGzaiI+RAOPx8zDpsOR9HGaSjMD23AANzaADoRrNItb
UYJJmuIKn3gqP1nS0iEh7FPoC/ttI8pluBFyrGd1gWI9pOJBXExAAlithztS4HyHb9DbZnuwC2lj
mKritQwh8g+ziCtfqaCsbxsvfRchWR39BVre6DIpVgJbrpxr10vbHwQ9ZxYUjTeaFAkTJqvl9pSA
acjGLmO59glLfnakoKvLG/BPqX1Z/Yw+h9Abm8fqDzuReLXngBxE5gEO5ed+1I/vlz2EtbDVCuJh
Oxs4jmY22CdRb2on7hocAr4q6I5gKs9/lCO2Glo0Vk1PiQh0NEqJf1Qbvwztao9TvWfiR6iWUSxl
SsMSyVsXk+28dF+uKed1B3VZfml7OrPN9wi3AqkP2oLx4Eh/PFu4fd7hdLKptg8XQliXtc+LbSCj
SjNYRGE3uvx2gWwthal9F2q7z3Fi1PlT2LuxIUw22wMcjCQP9JjdQiSDKPCNPSbPko/dFFcSAWW/
GfsN4Yk+9bnBUlS25yijrUeQIzqp1L0/0inWPWtUP4JPMm/O+XqPzb0ioHhl063t8MJfeYfGSALh
ny6KfYY/6qSQ3kFz+rOl9yyXxF4PsmVcMXe4ok+3ERS/E36wz0PG8/7yFc8bnYoCGp/9Dz2eeJMD
qWukiulrks8WLCZ6TkEXqlDH9G0S2Pja4kYr5kviJhAM66yxZnBC4RS3zpIPbaMMuojz2sNciiQt
kmk1JJAFjTOUl3LC2o5qKIqBJwZXIK5fAg7fGl/l2wiUtUkvtZbS+S1kujtKPvEE75+w+GCVT7Zv
t9nukcCoFvH25OnIWNkfhVUmf3x03q5V0woyhN9ng+pDfH5X/IdwTYySYx8TVm8cWjv8rDkKG9lQ
tc78LSy1d5qfNcyCSUniTzdVgU6ZyaB87gF2hCU9ofYsFjS+v/bB8mc8Hxc7C5oB6VneCRft4Tb9
QInUwTV9blhp++uLpEKawWj1Ys9gEJj3d+w0ktoiEJwZzUz7Zvew7hThmhnQ1Uy205i6pqlW9ZG8
ETUrxStviNqUzIj2bSd4eIkum3WnlQnrAdB40uu0M6nro6UO9DTIr9JVxdCDTpPWJ4nM6lkgThP1
pr7/BBDllJgOBru4s4gsM33e+p9FcwCi2kUwgGLSId7M5/XFv78O732KICfHlksQltT0koCJuwK0
hl+k5TljFmHSG8HBSML7HCQR1DnAWoANbhrqGQedY8Y9A/ZjJ2TvUc3jU1H3kmzfrcLQm7vmZ0+b
/0+cbzgGMWGl1TfWeZfQvJda7osG137iJjGDHV7yEZ+yKCSrGaBXWDt/AMgkP8qUTQpnIJDoP6ty
Hjz7+u1F0UX5so2JMiOJl2/YWOg/v2utK5q97sg0DwBAzhnno107VInZEyvedDsTsnuRghU94vwI
5nwqgStBIphCYbxR/WPxADtZs4Klb9fpmvtaifbEZszUM2ltefNfi6ztB6eCBdP9Xf+uum9KHbSH
ZBoedcsjl6O35evg3aNKFH9Ro4VC+gGr7pfTU5nwd9DMfopVMv7WJ+uh9PxZOVL1L3zmBOHIiPwG
HIhf/ueolEVQnHq1hcwX4cSFH0/4ej+Yi+Vh0WNMzhWTJCH3zNKV5BB9AALiKZ5FcKaDeS8uWv1x
uPUPJiYYXwr9gYTyfCpM8XN0LMHMXfFUaelWwRraeCgFZ5PQSAphbv0WU8uy+VTiZciHVmilaCbm
NSCDHG6ZVdSJV15WEgdVCOv6YNyNv8xNkZT4aFyzizFDp/abh6fwbgZWw8OznRQU0AVMZn1cYVrZ
gx9lotrWc/9RHJgvX8fKLt73bjfiFLq9pDCBHILVY5ntBK0TZOVPvZhGvsroP+p4WI2v/a3H90d4
U86JkJHcO/X75rNEEzqyQ84VDxQhcZr0SLujgzkcBnNDzaNZG259rpslwRw/4ircTRDh2nD5fQAx
MuUGo4kypb+oZX3jNFfj4asIv55FOip4YHzuXEQmAAL3JUZVqdY66gNIoEV3tw5XDi/uVGB/527z
i/2qNHf3VA+IhTtajgmfnzjn6VZ4Gzl/JAHlus1S9gH+uNbn9rgAndw47OcL4mi/sgRJisaFBQYQ
P9e5RbQRug/8f3MmZAEveTBqAOk6WAKNTnPwy77C78jaigUDxUqpoIIAmgw4TejhSNRgA0v534Ge
h0m0Ys4E5sgIxLqPBNAksloaMdzFXsKmc4xfRjsJgTQUNW240uLLmqLZqPXMjPZezTYEBSf8NCkC
SNHE7PVaUbxgoAxM9q6NWTjcqjk5JVwgSRn5XLy9gDR4PFVx0d5mFwKaAYkrU7+QhkhqKTOsarnO
e0732rRWrsmNltDe/xmRNYOwtz+gAcSEdNoHXCNNT6Fgr9HCxkv1neRq/RDmct32RvYJiOKke+V3
fzgjGgoDIndFGLtzgKb9iMqz1ASANNQ/N2w5PVOvQEN8WNFST83gHOmuDiexmeMWtij5TLz1qj9z
e7KaHVIv2YcyUqw2SYkbRyi4UYtWYud8m+Jb4dz7S88DGunR06v+BeFtSOTEQAZeb11NgrALxl9s
2sw32Z+UCZzRDwC075BvQNof92qXxsDyRUtzWfjcDGXOJxclJaRnbkSqTGqqm+jR4IYzVYc63kyF
H95X+41By1OIGL3a+5Ve7YPjLovihWcTSYVG9DvnEbASl6t6AX5Ccv/WBnk14CgQAElqu03iaWx3
Zeu/N93Dsc1ZkSAjDyUq+Kt2nyJaAPCiELOcbqQJ1Al7N8uxyUA1mmnC5whL8q2JFQuCqrwe+z5I
D2rOHCYvWIGPlpgUh7JBijldEEgWVg8xGXUHLEtXhin7+4eqTS/QKEYjXcqIoKwwZWMwQKx4KbTG
GGeHWMJYEKuDxal870Phl/4r2Em+uS/UoNBY41fE95FqZilYZz8ciZ1SurZRNu+clwLuHt6mGtPU
JV+3/QX31RQGAiuQplO93MKqu91WSIFuEUL9xY2ATpxRUmkDue8WWPyjaEMMTrsuU7tKWymPR6FP
B6rB3z0S1HtjEVte/ai266j/+0PiAe8SjYQTMy4IdNG8hof7t86JnwrtOXjhNjyEHxuaY3G9hZPM
bry/uBctb2RJQMUPRXqIhLMpOIPrqoGgFC1Nt+mIBZ5G135447APD2Bo0000Er0NQ5zzWr463Eqm
nryvBy5EQyWRkdxQZAbv4nHTSC4U9s3cmcZrEojdGtgz5doijVy2rEHdxNovmbRuPnTJDg3CQgha
uAVgZjHY1UJlAu1PVwIbnp4hCu0QnI8ueAXkm9tRDmQ9YOzddr/ZOF/WWBmYL48dQ0ygpT5KQ/ib
qc1hsl9IzHedvIad/9JpN+uKemPhx/D8xylJzhfvkgRZC48FSkjryMeceunPa7yzOIduKvS0/VdV
l8y4bncOTizQAFr264+7/aHaA8WOuIHM+/G96uidDdL6btsrRz+DhGZRBx1/SoGrBP+4vN4oFA9u
BC3fphAEXBNoC4KDuK/BWqSJG3vAGDgljLK6YxbYdGooW/MXyCdSpryAbEzIMK7WOHDhsCKDRztA
//cByklQw7DsPI/jQAQr9KLA6k3u9BOweygHqfIw5pJCRAjOoJRI0KrymJDFmwH5rZil9NtJaVWo
ihc6LSC9YNfRZBx8FyrwQPhl70MNJfi9Evk6mF08as15aNhjtR7kM5zA5n4OqSC94ODhWYQ5cN2H
XtWtxDRa/+I/D9qDOwLkNX5NDa2pJacoNWoz1oONZilldAGS6QvCYgkevPCPDg2Jb1E0GaNb8KK1
I0VipBxqO8dvt+b/CK6KnD1+RCxbVPmB3JninFB+n9WmEFFkhWR0z/tJJuBQgVKnI8NnsftwlUlF
bwGg/C3oXfU8MReKC1uM2tWG8HAlgh3NcYrO0tPF1szTsqhNDZ6Ibcu09kwtiLD7BF5kzdvaUHk5
3jW/a1FF76Xn4MeUjYDCgX1zm/2ewMM4Pf+M8X1lBgQNQwuuc5oA1mqg+ymaG4ejD9kC88WP0QJl
VJonnVofgD62t87vVYh0ZH5BMB+tJJ1ppDcKXz1DfMDi+QqWZzbdCxzO6XvC3cE+wjOubrlpDJOG
sBrIbESJUQOQwwC2QwPgSePyLGdDsRv8X9n6Pl6F14sjuxF6aX6nl5Y1UuU4F0f09gdF0k+oSsd5
Zmm9W3W9f2AHcrDkFfb+vFWQCAUNrSWQMFPTLHTfm08YIVwO4IMRVeIXmFSsVmOe8urRyR3GHZ9w
mQw/kfU+D57KIssulPSwRNVehr20zoiSh1YvdBXGJ0aEa3QntPB3nbk1Yi7uChligVv0B8kQsNYJ
khUqm45BOXMYR4QgDXLeMihv0o1LzlWoWiZyfyxafk52XN6tYkakZ/ov+oItmpdhKD/oh9ORxWst
7H5fSNXgv1YlIPPWxEgnBrQOIepMXkSv06eX55pBOONqZYrxkLY4rojj0myqmbo8sFPTuxClGU6V
fGTQNHoYV7IPhG5FlheSVFuZ6Nu542ZONs/f8NzZP0Cmn1AI2Wnzp7eG2mPmt0tC6OyDBZQHYxuE
wTKyCSw/O0QtWS4nkfzzGijWLP8ZKLQ3uT2GORB7ebpzHzCkjKQdfoH7yZ29lMz8OR+LzA/QUkPW
ZTQ4J3l+Bet8HAzfmJSkEhHIMyt8nQw/1knNhrHqCVs7GBZjeQEK+ir+nZBTPUxWZ8VOYO1kmD0D
JJSYb4N/UAlGRw+InTQWdQVLZ1bfza+8D6+ISRx8eoC4QAAn8/ZYNp+MCYT81KRJyZ0zseI7sjzK
Vmz5PNPSY0cPQD8F079UnQjqsLelndTi/5LzpYsEqv9YdrAYF+A7+uy3grb97GPRI1WuaP9Ka/E6
v1lRT1lbRiJlP24ZpsrWBz63i4xpZ+Ei3LkGTrIJZaaZANwO3mDfiGBI0IHzRmkDwLFYk7t9/F1M
wX37Mtj2GkB33rJ8Sik5TzPJqw1B0cBZu2a0ENHQli5EUB/PlfwjsFiPwyv/N3Fm6eJ4iEFY8c5u
y5+M+cq6UBPXcpUMBar9UfrF3PiZKEFBqm9eouU7jfAyxnprZQtJWB8Du4CyifGeU6ri1gwE7qKf
ElE7LGtpO5qz/nFLOs9Hjbmn8hpFH6Fh/AWC74zmNdYvdwB8si+4YxvoDG69nudxR0xC0ajPHN60
hF+PAhqjliK02YkT6u2cjhMeqSBiSG+v0OXCMwWq4XGUBxmbb+Pg3mzgIvZB0z0GLNeXzsZs+WBA
u0vxFhCymzz7DLk7T2Y9UlkWNOxh2TFKCgRUtpCiulDqLmoaVVeWQU2aUgky5toeOt6DgMTyXZnb
h5sEVhY3jLrViazFV6b7lxVQNCfGgmf5+sp1q4j0dJ/ghr5go7lNb6lpJBQKgGuwDmFn3hns4L3M
Xd9OeQ96q33kxk0H4RlZiQeC91D6qTa/ITSPeoMkayIMNKwMkaMfSPij9bxUU3CydSm0TPEXTou6
50KYFAjSQbiORqCua/iHzmI/LC6i+GcgVXszUB6w+mpGfWD977J7qqDh6LwtpoNg7eb6fpgqYw/g
ZT64kddtBUUwY4imWAqccXcOegImXaTTZ47SEYIzL64VheV/8IVP7X934rimmKyar+0eBAuuAuw4
IaWR7HZ5fuH8AUHx/zkgrUSdSKSEY9i6LTgwv0kG69VPurVPVrGTYtLH+i55SSwY4Z1zXb96fCmm
J0jJ1KPoV8ngbViPdiXss5+jkUqmoFgciwaciiuCqF254RV4oAFOyhet+j0VQtpIAz74TJ0exSju
eAFZ7lGP0fCrj6OKyKfMmAYZOhzR7sWb087y0t6UAQiJO1RLYceTeo9GnHxmujNtZHWtAuJEAoiO
4uGvjqNDpNmIB0jvmMAnXHdZ+CZdHbBrmnMcBgIOh7YQFens6QH0D5qeizUuFjQtk9Q3hz9zF8Em
1LZHeIP9TRoC9Bl1RjIVT5chC6cDJj4Z3+aEucG/YS3Dof8A5/Mzx/onW8nNqMhOX4AkC+5lGVri
pYi0PQHz6aKMDTlySnMnFuu3uwUA+ksUxzCox9IzTA1LwiSRP1F1tnOtW/mAkovHmSf6EkmQcrDE
35YWeNXG+0az5yArmoAEkD7ILyGEYmxuVI20/6tudrAWJRZ0yx+0sARGhPLZ8bJLadq1Aobv8cDm
6gEUiy3HgfT4uvjhb04PfTc3O7SMmMiIhF4eKXr08IoMYmf1LBP+ux0n9Lpo6tkD7iyc/l1/XOpZ
TV1LwtMktXApA8bRFVPvt3VmefaVLHFyKTCHIiCb5ruZGD1XO4HKgN8tVSG6mz8Mp31fxCz1p0jq
NpEP3S276zVGhUWJp2u2GJQUWv4n/FaLQb6cpEcMDcA7umrjW5C4U/z7yKZOwpmRHuxB6R2POHmm
ekxD9i17j9WATIhWvQ/oU0tpWooa8f+1dLy3fWBYLOSftwRih2eMNaVmE0VxDTfSfC7DNPYQHRUA
+I7S5tSM7dclQ7mSkSugyhhwAe/IfZLyWt62y3VlPZOcArVAuSADQz3z1u6K5x2Ila0WrmlILQGk
mCC905n4wUwjx+UVUY2xffF5wm7f36WMpssQQAYiZXO3dUTVcPHGPkZRUFrPq1OzoVh4z/JRvOMF
V02tn1arC2oPXOgWh3Ih/KzyLGPYYzlD0uduxR6IiXbjzh7pyHBE/aEhip/bZFEYT/AxaTNnIcEl
3E3KeTuHsJ7Nb0036hWpiEcZdc2992JJ+3etAsVqtuKae1tpx4yb31aaJVxrXDpE94iPmbKVF5LP
TSoE1ussxqhv6OwdDRqF32hgvYgb6Ki+GSpp1ZjnQSYOo7PXnf+3Qx1XLy6d1t3JdtKkqLoU+VaX
MKyrYOyowQUkAmOEUP9aoidu+pxTC+wry2JBWgGQHPc/bMoXR7tID4hFiV+Q2H8ESldQYAhKMO1r
/4ja6fEbgyXCmlKITIPTew8gV0Y35LbnyrkhcaQhBhDqZ34VkqvJktrLaGJzODBwVmCVyld9wX4X
WOsbRwDuNJwkk9AnPrniqjnzFzNFAjDE22QmQTCksodEoIpyyxeCVBBDQNxCEmEkrqKTPuWynXFM
R6bJN7ifVh/Rl7UgP2T/Q39gOPmt/zUIRY3b38uxgWT56Mj70FDKd2QJiYrk5EFShvUZe3CmxC8l
fQ+4OOG/htteJ6tKeG3T0xnOAZfTFZGWc+tr+nt9a5hMx7JrK4qoX3Ndqwl+X3NnSMzfmM/PpcJO
tk4S0RLgxJuA5IEuGWTF1naHqARi28PLRJLABtM9//QM32BeXbn6ZT8eI7Y8gb7jUjtqqr2aoXAe
T55h+i4Ls3SYYJPwqarguatgISF6/jBscOAi2uIjfNSQhGxrf2LnzNnd/9gpCJQEKlHFYMmIwk0q
Djo+Eua3vdSn69Hlb//Mw1237VICYxKZLBvep43VO9ZyIZedMsn+Def1WxZYg/w8Bz9KjcsdLG9S
OiIuzRbLfcRa7qYO7xrkhKNP+gSd+h0TcZ0j7ukezr11uTZWMT5OnGAtn3G+K18TxT2fQhWnl4yy
PDTx498SzDq5/HZ72t1StbiROpyWKZ64Z1FoJqdvNq7PjH1SIiSMqOEkXPBZnBnyx63IzT62YFpH
ueaEkVkV73YupbgremBynWWHzp2jleyC/Rxp4j05S8DEQdrVY/qNSf6YlqisUNfrxtResphSn/ti
UeOCkmJ8ja0AOMBPvhOnR4fsosQ9oleZjGzev6nvN7KDob0wS0RjwtrGuPBPKtKaDzgr/rewDaWv
T9j01X5twWVj7MzjQ+kmLDrGWjJ/1UxQ2/rUuliqBVHoMg/OKkePOjC/twtMabPlxpqJsNJsLO15
A4a6C0hZWP2GkWqTESkY3mBVkqaO2b66MZiv+DZswIq41fqqY0pNU0RVp3kIvMGgFUq8AeRfaqHG
We7GO1aSFv7t+h1uboKFG9u5ufQUwfoZYF4nltONn3DNFHY7yIWc+fa3ChrDz7srBbHVp6d6eV4d
MF5Dzn/Oq26GfQjeCqiG59byIlTaavZrAc4AHr6he1z5gsva4q7hkDu+Z9arERSq9sgPok2un0Gi
UNEeQP9bkZRocRH2Zv0zr2hdBkuX20jNOSmWvLo7dduJJ65ZhbtzcKfbqwDwpITz6OlcnlhQbtOf
aYJCcIqMGmTivhMNOltgD9n1Noo7qAUmTVgGalzyzEoymQOqeemOEnPY4u7pPtWZ+sWltcuRDsD8
yYxn42G6zept4Kk0gJ5jrM8VYeYYJPfpY0oZJRNiiWwTZrHcE20qNoWioy/7Htkuog4V07TQsMsR
N9CnfG070XaRaPl7wNDdWe9v2kzQ3mUykDcNNqPUkBT6FGOGAjGGnVdKmeAJTPYYQ8D+eTxs/ibX
0eYfrhhxoWsWABR1AhRTv5189Zp+V41afL9j00efG0fVuYN0AxVVNKkXa9JGNf5FQzKwhoK/K0sP
/bBiOLTPkaTIl+ey0b6uhkleVPnsqIzqS4lkXhiyRhah91J8wjSnaMwQeeIj3gRM021x8jtggx9r
TIMuLckGEyaMft3O/BmYigynTJ+MVOxHCaGtrM/jadhQer4c0kv/Ph3KGJCuqpkt1iBs8PBCcAZA
hGPVydZYR/IL7MFsY3yzFGTjWZI+FtPuDqWQXHAi85RrQO42Vt/0QdxBivt6NR2SLqfnbWagUrus
JCgkd24rLglhPObffzCrDpnZFXHeOhyWCk7B07aY2fObK02GjHhxzLaLqC14drXvSh3gT9FKTvQw
gb7gGgSo/ABt6TEjCrpFBbsiZ9DXOOvXnrkFfzC3O9S9sjS+rjPqn9XSYv84eR61buxuMBqz/LGU
6AI7FMl2LE37P/oOonxCsHCz2uEsOrTQ/e1w7lyjZQEtIWXOHVLc0gmxDxrKv+eTIEILwW1GNMcG
oEOSqMxdC9EJ5s9H5QmmppbZuzkc9jilPF0I6kq2WbD0jhFmY5F3lYpMMzTnJL4UPMsbZ6UIM1B3
e9K1ukEnEmm09hT4mvYtmrMh7v/DGo/sFcc+aLnOg4g6ccKTpg7KbNzFbwVjOsrczyAIvLQBXJrI
JIoBoxb4G1SgjlBpJlDuauB5CuD0VT5mLevMl/6JWOQ+wWGeWuVZrQrqO+5g0odMY75J0LdbVMss
DcGwerlKK2DxCyFM+TYJMqQn/b8ZGEx2lPUfnwq3vmNKK19HXPRsoEBYZzVBh0Agxf3eIYOHgCHV
z4DE34gbcmCFYh6bNOh4/fu0d6PyiJHiLX1z7gKN9YhAfT7BAEP8uwpJYF3nvbWT1fyrsp9hRsIK
ALdgOT5zC7pqquuSV4Vove0mnJM/+mTBmxavS5CbiSyXKhETp+N6C2p1Y8pn6nfymkPLVLqVd3s4
O3n4cHSBwpFQ132Q7bASTbf61uo2eqXlrf2KufLnh5ndFsbu334xPD6pVLjKo58kjFq0SxJ02slD
j4YIV+vy5hoFNTk+8dZmzKQdo6MUvM30u5SrZcw9fEOeZIzHFrTtfM6MrWYt/ZYW4f07WT7uxDi0
OmEs3hnIpIV4Njv1HQ+N7HHKp9UCunvI8RMfszQNBs4IqB7ffSaSMxSI00lWEmII52ZZqDZZ7bIp
bDYTe5kFMKX7MMbnsNjEN7CTnvG+pbUhQF5ACsflyp5QPj6ttQVupXnRNEsJ30vrvoJVSflS9MOA
tVzIx9OgBZznEWAbREyPs1noYe1m1qqZZ9UIiDlWyJiPLF5MNRZ80oNmsuWBxW5OGWiQBVUAKQWk
IGLYMFRLbRnn517JmNUjiq6flBg9LrwFkP4gDgIkiuKHdHsYx9o8bTxO8aim73qATS5m7nYXJ3cU
9BjBNJvwTZWev39PtOni0Fjd63v/dixAApTox3AaBm46Y2O+C0qs6HJZeLXZGljcLo2Stc0EWo0Z
ViMbvFbFpq+htLdHZ0OsNceVMdKWb3a9vYvT1YNgLm7/L8alzmGNeaz7fydg2bEsoxY8k5MEh6+z
g6mwspoGYm6n5F7m2e7hI7RrPCGnZfJ2eFM/ZnHeYCfU/eA8q7UFRbs1IIoE9a5AZAjTpuYJSiw1
zvIXg72W9T0DLyutmuY9laosF8PQmTy+PF4nAwu8iscvZisqnhbWobXXPy/sHH70hFtSCL4yJgXJ
E8icKp7c0P8exqKhpoou/VWZjd4YFcawe8an1GuY0rGK76zuElBrVyBzPkfEdcTW8yrkyilVT13S
R/P5gbKnAlWON31I+TzKpP1h02urT7W28RJ/3/wQho9EswRYKpxaQxsz+qLrYnt2iSwcEp5Dn8TK
AQ7gRT9O5ItNoMP8w1T6tA+9BAvm7Rx6yeUW6ohWqGq97WFXbnHk/RvcaMX5AqWxC31GMzPKFUVW
Drx+H9gjsBOpctsJHp/bVm2zr2ZEnMozTkmxs2xM2luNzBcsxtFRA8deYcEZXZVcQCGQHo79EPGY
lDy+EKoRY5ZD4Uef/wA+XvsJcwPg9NtC/CZ68WRUa20XNz27GwuKFCdO7bNvquUW+EDyuaZ37rAs
jzlvTE4yk1hLHvfXiqRPMk9UAwfUipYYoXC0YXQApDBkB02y90jnp50WOcRtyYQH3lsORQEFqCRC
UJyJKfHS0sIMbcoykQy08dgbEC3n4zHv/398sAkChl/BFuBKafkzIDzxPoaBhqzr9ZN/A7UyfLWI
iOii8fBNopslT/jccfH19SNp3cj9AKZJ8PgwFGeTXyId6MebVvZhUjyPJ1dIt6g3+3KT81sEM/to
fc0cuRc8/EeSKth8WrU8DDYAb2BHIvK99/05KrnWjtVQqjxmXrRP+L7fbgzr3IDbPp7RefE9pchI
u3yjMql0eSuestWQAbQzeBsBDVT/AfGtfp6Mtthw6y3MnJEX5m5w6eTNGXIQDGtlbPoGdbH/t11f
ZaCvXambdcZWPPvMD0pcIHePJgnin2UX+ztENgbdUGdznAmp7/tF1r9Br5FnGT+HjKEH11Hu/VMN
sEhsPrVxUMt6rivslsEIWSc+PZWEqfKh9pcJtHzMDQq2OK13ww0Up/LVeMrf25LYAqZTnR84OOxA
MnJqEHscuDD5HgS19+n2TfS1J6ceHkhO/x2kVchf1rT49mBigz9vedEky6lCwoGJqAdtNYU0w0v4
sB19yoq3zPMgDGh1MYeCyrE3GNlI76C4ikad1CZezuKloKlKczsDvyjpErHrzo7x2lKzLlYTV/np
zYWNe0mBLXTTy/TX+n6m18VJYHcylsQn+C9KBU6ie/pUMTgApmjuSE2koyw4a79GH8FhuZvRcOll
Ha6VtBn7WyM4dD4u/FXde4JbDHQwymp2YfRsmVMsGO+AgDqVMfBmioJnymSq9z58/iQi+ZOPD/bV
yHkQujwVCf7NivvaOBuE2QgN1YF/vXNW4ugFRbYsEsIKxoKPhtVDOGQGv7QrPvWb93KV50cYxyyu
omsaTAb0GM1p31bf8oQPM6n7PaK9e+c4sWZKOQ9lZJ2b9+Jvsx8mXfh7CZFWzm1wNH3T1xbPHTiR
OkoB33QrxMKP/BI+v4N4LMFAFOs09GDRgvOePmOypzxQwIVmBX6+ZeaZSdzBfOHKGj2oiS593rB/
am7sWwqVW53YQvmGn3qUwZKZ+d7z7JGG5+pqnhc7kaJsxH7NNFgICi/HFWIoPrMxaO0Qgl8X45ud
a8da4Xd8CUwrmQ+wy3rcPZCvJRBtC1AiO5Dv7+KrkeJLdQCw2P1GYj7drg6Xisxl+EiM7/q5FYvy
W9VRnYyxlLhUx3K6wHTrCJdT/zjAfz280qpEtqM6nahDt1texwrXUmg2d2WGZpKcx38dt3IFxpyo
7RTZh1PTot6r0eSH9vN2yTBKiJ/4LzudyXjuCDr8Xao2tPUHB/7sjrawcjzbMf/7fgGfi6cJeThH
W/AZZ/iKnN+6fIfg6vfDVskEKICYjziAEk6JenOtndH7Cquz5U91BPn3SLg9OnXzNEiXJnSnp/5c
7PiUU9dzLYlu0ZPCXKBt9h8ETlWzHDwfRoO6KrJ1fyLCSowopz77L3t3uBPYf3rAcU19LDQXHOnK
JBHJdlrqjKVz2UIBeZjtvN9A+sWnvtO1h16dLTTfW8/zkTHAeb3tvJse9zgSVBGXpkwE/sfxGlw8
1y1KKIeyT8HoXubP8L3Mxfe8FgUDnUKuA7ALzs8gun4MCpoGkl0b+conpe/nksFpJ7scuYgd0cQg
1EDHJc7AoQkyOyLpfsz/8PCYRHCbRJWXN7fkCxM3usoGaDb81IOauinAnRekApJsxWG5WZyGyHzI
HCmzUdG5yUdFlQz0LbU/MUEdxte4XEG4hLWpxX/e/wD1wPkKicoRGR2C7/Nibj5Piks3dihI/1n1
hQ6uDKmdrSaR9BytRi15b4ymPPArDW6bRskwNO1lFZ9Owr4X4CGhemZSrcsNK/RXc+3My0cF/5tR
kaK/uHNMCF6q4ZHS0V8kZqAgg+layJNNbhUSbH/DW1XiyIlA2S4d1MoTdBXEbtN07zgtmjbex7Mv
WuIm91hXxiYDzHxKyutjIlGx1wBqg5AbEE4zKGO0VSZN/VPQwQXZn5B+wGwV0m4HkNxsckV3sTr9
vsRZ2LvGR57e90qGhbKE//aEnJwvo2stVbVghAD8pIniOJckB4ZuAS/Nh1gU42a4I8tST4EPOR19
0OqbIlzHJv/4wsNez51LFlxU8tSR/V6ugAghwUJ3bZkgbdfJUN84YApuZz2muY9u+iQ08aObg7WD
p5oA/m+k1AzMyEUSN+w60QlX19UNo6bBdzHQ7YyE7XkvR9NEpijJxqGkRgFEWjZz7lf0W+LumDnr
nNM9OahtIv5hubQYhnTEZ/iGrB/fF+X9FnRr0CjCmM7xLN30khmL6kFYMdC0T1/auJRFrXOyOD85
88AF6Re5MbIu3tyJFIV40w9EZexSwbW1zXEKcgLU02sykzspiHA9hwWGp+HpaMFcwtfUKk84zJZo
0kFLZvXi1dh3t+wam6b0Pyilp2qBlN9N/7e7QOy0e7zQajhs+w7YZI0rcIq0Eq8wjPDOltPg4xyX
b0+MGoW5vc5kxK/LF+WzmN2CCbOzX9zYHm1eCYXLeO5DtDXE+zBjb+ytxbkzpn8RI4GjtXwTT5tH
p3QIp1ReU1HFpQjZoFqn5eoAMRkF8NOUTbPuxef6KNoQLj46jKX96FCkjOFJ10ern8IDdQ3DdWaQ
9Ek0oFvzttPf5ArVuYimlVLvDSk8ghFTKitHqFJdzx8vYDd5wNhQS7vQczMQFePpGa/GmyhHO79/
BHwwTi9wfda7Bp+ZyFVwPmMmytmLhl4zeINCvG9M1vVmovyoH9vh6jXhF8MDVX1Tpjtd2wuHvD4d
Eytm8j8QGi1DGiij/mUzdnx3iZLYcRMVfarzcmGcphiJ1Zrj1OBMFhAyvVBGhyv0QvfTafOyBLN4
PYicMEA6xuHDDz+je2slTEvrjRmrzc0v+D7n2MRjTmS6FcoqKnt4XYwJ94Ai2CP46Jxh9WQZoeKg
bsaphz0v9+/jfK70npunGXKLPvCAnebbOBgJZxqFE8Buw0r65rOzM0J2rk/gFglnfBuWIG4ivCWn
0N+u2RLEnJopFIOUffFZUIvt1kKZmU8ymg943we+6mXcSMHmRT9/GyeU8JC9HA1CY4s99wk4n9iZ
9vUaki37Nah5v5fKZRSBLD0U8xRxRBTJIeom7hCZXkxCzwU+ETPuHC3WOMcqDPRn/MaMVDgj7WH3
C1xvnsr1l0sovxIiCIR695qdjD6T9kWgZU1p0gEAJNA5QZX2IV/ouUHM9MeyX1wXrG4ssjPzFCP1
Um95beXdxXk67WqdC6hyvyf16SRlPXOwmAtzNOk/c8EXPhze87MSGfZlNcEVAbGPnwkfsUaVA9PN
fszjscdk7DH+rSJ+X/gbYqXXXZ0svb0bpOYNUvWe9OuajqV6Io6cxH57jXRcQ3q9eJTsjZzxdb2N
eaTDrswJtLAnYpR1CQ+ks6ZQXD8qCirY2teg3IrupToRR4YwKg0lUNqVRG+p49CuHxK/cAPSwEQa
fVfmcGO/8iIuBYJ2n+NeqywatOCJWWQ9ohVxwF3a4fG9SVtbcHy4SorYrV8buj4HfKZTezNlevGI
oSLyQQ6A3JyQDi8pqgV5cKmAcwpKgiDRQdSe1vyan7fxo9q2/iPwI8po3nTeP8vzZ44xemMTOy3p
H8WA+UMcqAsK+VKMnMhg5o/Mg43jgM1xMdizQTi2nN4ZclOFcLH/mlUhKwM8wLPq3+vjA3L2SUwU
tJjef0PRTMhEHxwpNQOQVis3pkt8znDBNUV0tgpIi32ABsVpcj84d9lHDe1pavPpAZSBlgg646ts
QS3bm8G9WZL9cy6f9LMtH4/6eOsgL/CMFnOEkuE3Id9TxJmiGlxPoU8Kjn2ac0xNJDXQ/Z95lu7d
ceRQhzhQuB79FhL4+Tg1mtmoqIWwyBYJ2mNwWFdRQzgeXv4npADgXThQzBmQ8stXVCcgU5GDhx8L
FLi0IedH22vj4b/PWD/S9iIt6brNU2eiHSTWkhyuYemhYWwPQCcL/p/FWgtNNiWLHdwkyQBv9n2T
0Unv+Mcaw0mC1dgxwHsQ7bVLe9AX46chI30gTYFq0clEHxxHuC/2BLkh0CokEpK3JCZDCG3SfgfT
+5thRdaretzPbb26VrKfvhtR8AJRLKQwOJCWMtaV6r30AHFyuRGE193vZDg4QEypAZQlcwMrV6tB
9uHH0l6jT6ssHAIZWBgJ30OjZAcUBAZX1SMJTx6HcWx0X/uIxCGPxrhuzC700lzATtx1V0qT9kdn
McqIHNZ4ekhhxlJ40LwJ5hLO+jjNtVsNNDXmdO0Cdm0zYnq/aPcBqAnTBPMWiKsfBBQD9fYq8/f2
p+ttm0ejQzVhyw1AJQN7OFYjozqBx5W0OYChcSeu/0Tod2oZMfAQP2xysVcn9eFk6YmIoeQADOGH
Vd8uazcC76CpqnunhLN57M9lfhKOlC+Dlx+lqQSlukWwZuUTBW/17vfmTirKEJbCP2lPlGQgQ+vD
KwHqaNfKtfuWcbN4Dz+A/s79/bqnAFJyFAjJTZy35GK1EW91qUfkAewB9rPywBjpL2aN7iRPAcNL
rQcWIevYkiXdZagBnhq/aaTnYt+F6UpUNvVp14iZobcIRo9v0dI/FgWoTBYg36KjDUl8AW2mX+FF
bhDWmVzqmoAkQeImamiwi6+GRCy/vrJ1uI/x6iWVf2VjU9LPkwc2/eetQkLVaPIPzMrWBnR/AMVJ
cW1kClLK/myKlApBPtQ+2ioGRB/w/NL0fQtf/nVTpzYEn5xLkpWvtp7V68/HjBV5OUV4qvY9KHt0
Khqk/jrxaVReTb72lFHvaL8cDPaZ6HWpS8cV6JyMQ15ssOvwoBqwIXhswH4vZp2IV69D3bke40jY
xJ55CkLLZ9jS/jN9TDpBd34yTZrfq3vuUFBJXbLOlz/ayu/qWwC1aGYBUU3kYdoEOXLcAykc3oNT
KELa6MoFBekAI6lO4n2uY4XRg1Ab2jxyGyw50Vv7wli6Fy9dmiEZOOaWn1lyte4x4w/am7NQR/sh
LxLlS0uODBLzxeRZslAmHUZrWf1Vr02uNR/2qRUWiEoQb9YkX/ycsFe3nyOkuFj2iW20ZU2Mnkg9
1oVqL574AYU3VARMcHHOYbU85vCpMwyTfJFaKq1YCFOUXIkWcP29As/BtgFOpylGsgszkmdk0LFX
Qvqo6R8y1HC8rvN4dnyEA0iIzlFTjXjW/rRRA+c4BGjN9wFMYdCmutDKlTuJmKJlNkKLGCcnqwiU
FphblPc/isHv3RfJ0tc7MPkagwXHCXXU/s0jb2v/odDV8RwCHe7TYhal5TQF8VC/Tbvzc0sVxP1T
Ki8wT29gNcJ8nbOfUPLLKZu0LChZ0ZUCgJVhmLCpOA67p3/IpI07yoSJk1riCiDZHi+Rb2MY8vu1
Q9XbaC1KzyjvTDWInXkHaFqMyUJVZrZeEbM/rXDgFekaJT1gkZkgg1w8PK1DFs1pXl32OxWbOoMx
2ey/tbAiNE/Xt+V1nbqcVWZxC3nBvu6qTpBRGK+hlfZYRUbJpwFKqDe/9OM2japWBT3/kVvq+paj
H/Gtqce17wpjEvBEJQza71e4VVdzv/Xj1Q6yB8IBRgtspg1L0n3rp0syETXjHnD7EiIa/P+hwNIB
WxvKrQx8KJsUgzaB6lQbt0GVyhdvJotRvo+2t5KOQGkYlK+iPnXSoxZkydUo8eh8rrSm0PRVf1bB
REX0bvt6+IkdRcToiAMMtl4riS0o/N1oVzFS6E0abrQhXIrtGlyU2UxHlg7vZFVRAReKPhLcKBTa
zh6VnhD6bFou7U/fa/qBbbdeHI0ZXglCoBh3XJxqGCeATLCMz1ihbsihRZnCwaPkqggWRLV+TgpO
qhNDC/KP/WZjvWY22Cu/1O0pXu6iN/0q7i6gR4tOgApe7eFffA8Nu6BytQIxivcG/Ec5sjxXIj/v
0Udw1mSaIrT1cvh+ssINEunJx9CKVgqB02Yh5jt40tpGCt3S6t62JrS/JDqVXtnFWEP+S9m7Jurt
qx9q81fk7k1fDmpp3HZoD3OG2G0PGNqPRIaWORBCZieuVc7EIXnz+L9FGuOUBF0wdswQTXcDDHSt
Z3PeLHmvEU4PkCNOjA0SQthdnk28DPl6W8rGlf2bk/L4cviM92XBEJIakfClLKq7EEdHqaU9BW1n
1l1vwt9qFzAZUH/SVweEctfMbOuqlHXthTeonkBhQ9oUvhZzojRzqNtDh0r4FKPTSMTuRR9P6SCK
Y0qZS97kkpmIIPd9baHNVC0Cb7Ff6K91zavjsSHzMS5wCu/vUdShlPOvoR02kzMd3QRSyRgBzU77
XBQi+LU/7smtvL0h2kaB0fRNvGG4WlDeg/euXOeiZCb6PPpqtC3AFARbh+IBjJs/FEaCMpmHGVQg
JGAyqg6LCFYFvJuYE7JpKDXdQhSIZVxOPwfRc3UyseYS6IPDo8q4MvdDb5qWcjPR0T2WmXKTnfIf
RiQDsM0y4e6v+cJ7Rr6IPwbHx3n7TVnEe2LfZTmaS3MlEJohaKHFGl4l5ZLjSU8gdyePWbSnjRIB
/aEQwyVyVlRbVkJCVjSvlbBv/IBlhYqReZaznwF6f91iooDky8WiV08pQmAhi52WMswIDJKSWBl2
EYSDOewo49rNKremZYnDfb99+8d8jGtcJ3MhMXHqtoJ73pwBpT6+tgMwVPqSBZ+PDlaauICeSeOH
pvVuVrpPKOQ/3wbxTqjxVNTlteGNtYFzWQccx6GPAGINVo6qRiHc0aw0/xWmW//EdgliOu4ej/av
O7oRO31qZOZCcOezP6xDvfei0JDhlcIw3bu/cDhcqGBgU3YWN3Fz5zGxPV3bSxhA45NFW6DSNOpJ
s4seOFXImdlcyINnEGpi+Jtv4GSjH8s3ZSpEHcgHTLvVIKzbTnJpfkOX3b8SJeAIUgwJGo/0j74E
sCe+oodomUtrVFwMqiPuQC27FSRBvfkRMpbOp0qUrPBdJZrwz2TcLxGzqOoff2eFffOcK2j7xhPr
bS/1uo6EcX++skUgjDxA//fthkrkAPRh3GJZGdLAtGlWiZbT6mOnbOkhKF/HfQ3fy9wxJF75foXP
NLWzxSyQx04LOza8q8kH3zXbcJupqX3UoU96rYXaMVyouU8mIeh+m3rL7B59vqZaPr2jVNEOYFvl
Vt8bOmyxrLTOOI59EmfIybazMaTNQOPa8fkRUaiPRMwB/lovzeNokwarJ/xELn1JfI+ZEE9kgcjM
0ALn2wFg9u7IKSYV9Cod5qBRNMWDuVfNn2B49cyhNWZDw7G+2gKAFsypAKrxTGSu2l5hjd0zd/La
fRbDDzr2iD8e56yjHuhb+a2XdA5hmVffg/Il1YgDUay+txyj5qCpnwlDFR0fqMdKavh3DJnskMf6
o0DcDwWJHhO3jvw/zAp8kdXJur1WCw+SRZky4Rwz3ex0VstaT4wtNAxkoSrX+TYTD8s/xMbFM96K
CwoOTnBTq6x5LGF0exJ5+3AtSd9/uBULI/mC9mWzTHEOMOOin24Q3C3ShuENXTvM5pNSZBlLigJF
DHZDWIDVk7ky30CQyWi1UnbiVay1J+OxdlE991l9d8Xg7QOwmBy+1NCULacC/quNcT1MnCkJU/cq
u6PCT3V/jR/hEIGL8r/2et7Xd34w0agBh4DGUm5TSZ5VqGcoxLiv0I1qMIXlqbc9YxhTuVbE91YM
qHsjA6ULxDF6Vui3m31nf0KMRlz4I/rGhm6T31USyDYNKTuRlXWq9m+vYEoAmSC5OQg+xL5XeI3k
CcpiS/87kj3e6snJ4csMdq2VotEto/SkxAmCCK2Umf7BKzpg3v6/kJ6yk8i8HBRuSsJw3Jl58laG
3PL266sra2eJCDGCcoHAwD8SmoIM9jQ9qZqK5pPa7/XIWkUaG3bT2JODtFW6rSFvNKbAIrLTjUSH
cCuBkB0qcti1yJDFKH396fBeiyIfoqS8O8v+gb/4CNLQLvR6/x4zLVsNfCBOXB5jLLQC5ZOEosut
2GSyWrnfeBje2cQYGUZUCYcHmFnqynvYY/s/A9b20djufP+LypYNQw8gOAdX2THWCH+/a6CThNRP
4VCPd+nOPSi69atPFIGzM1MFIzNQz8xEKaEL+6rYyL1QP64K/7oluWjJ3U05AS2fz6xLXVhjToVj
I8roOfVW93ysf7OhDbxyo0vUliZo+0sNa9ldu3CpYzVNYH8k3CI6mDCFUbCTIEThA9F3A1UqQdEs
r2fk8IrzULZ1t24mXfGW8zCWyE5fXGo+20mwyxqXrWJJXQ4zZkX8sVGSnq4XLC/zlVXLUofDANN9
ubZ3DQr95+wBo6wbcmMHYUa/9hvzQbzyfNegKWedWv20uEF+CTJnX4kXNribAQjx+WnWJ1LGafJO
oWJOIBtrNeRAuEaKJnC4Fm1tORzL1FMXjZjb9bSe8VOLpT9h4ToEgRI2Rt+q7vxJyoXMeMNdxrPC
5E7BxFGBUkuAxUluLiIE0DaGpHTBRN4NuZ9fuo3k9egM9uFeert7VCoDrmEGiXi4C6jvYYEdu4yp
p/Mp/mxWnBtQbyR52DBjuMkhP2JicReeaHxzQ7/i1KNH2bTHvTGvfDYfFPumyrHi6emcG2IA3C5b
mmb6wedxYuCW4JGN5+hcNIRmALxRX5MGTBDUs3GL4FC1KPKbLR1h+GaAo0vWheV8q3zJLpC4ggbC
9LgvMGNZd4zoPP4u3rbCweheZc9fIvUlLdPQyqOSgNk4ciqKXdXnKLEmw8qLQcjoMXzwHZv8Pfn/
Iupdw64m8i6PnM6aluyIWGG5XrzWCtL6DmYrSgo3XyuC5HLCM8jAmIbI4K0Uoh++5HXjTHOmnjFJ
VBZKm7fwsHYOI8QBqh1/DZRCvS0oGFkPrA+Vn+KOuj0M5aWSJ0HzzEdYC8WwK8zvTxBpX6FaSeT2
KOXIyfgEHbehlva938mwbY1QvWDXvcWjNcAHIIOo2gebMdHLT129UOhv2qH0me8rROJJ3DZWmE7S
KaWqotxnhpfw0t8t4CaI9uwojzgdbJP4OmQLdgFSXKFV1uuI+lEU1BufZrJC1c0i19Qs6HXZ7n9g
TFpN5oGbHBHhZaZhSO0zKaEMq00EGgLG0nxClnJMAZSQPEBDXHwQdAVA9474EcUtCi3CU14pi6zt
3ai7gwoENmE9kVvfy+QIJ6fm/y3o+VL66ls+0F6tbIwoI34GHSL0s5Ot0SoXUFqWdYtHzXGCcBPK
yC96PISLjIF+JXEv+yVBgPMsO5uXSA+ZClfdwLUeD8/nt+Cb8tkF5UKdcEv94OBKMstjYoj/rniI
fZOiz9Cpfiy22Zf5wH/fQvc2VboY6iosjOpUZSdaXlZBI5cI9cbWbw+46QmNQs6vIDooSi+cKWZ6
9cicaxfQdsUzd300dGXMPIajNXe3aMPXiqkCuxcf6KM/r62+f0zAtaW0l9/tB+ln42vxi/d9Ttk9
CwyffHCgnqTSed6hC+9Lv1T5lAzht8c1zopkIHrsI6veoUgYDLXq5UJFrBUbURqoM1ipTJ//exm0
xun72We8kA0AgyXAZLxh1NfqM/EyfqJyFGxtU8KMerSHuoguzKS3Naoj2my1HbXHmV142JiD5LSH
1k1ayJQUwA4BGGLfSuaLfoIQ5PvGJ72ZB/GxRxVdNt946EV6L2NQWfcYnCJl2eBldaqmGgKtcPRd
4TQrmF/fcFD1Jwc/9M/8bCn4s07dBRBhg38mS1ZnBOGtD3HH/uY/AHnOQDOQRgVrss3nHpBtn4sK
thXq6e7gQkhsX+z5qDa9kBwXOypbd18fCc/0WZ/AWkBDiiL2NoDARpJPxYjrMAXM+Z8iwMjG1pQG
lxNGEVNY33UKHa9wA1KUKJMAiLnToq+3m4oIWI5i1XTKJCWausnJdqRTaAxnUYbpHp9ui0N3yBiM
AyxV4oTMkMpeCdvFtgs+4Bvfd+xRpupgfxS6iRoyaP3EenLu0yGu+HDjJJZqJpnOgIEUVmr2E1ju
vLuhZ03t1Tv8qK6ETwHJ0jjdFophWaj48rXB8NL8NF1e0WuflfEbMst6uXo6iQphgiwxOC9/b+v+
lU27nDUwHvAyP20kV1+IwEpvhdPrZjs8AWMCxd19eBU+jwTnonOvZRwAnilnFhowt3/2pX93WcUZ
dx110afF+BR4DvpVnbp2MV0I8M+M/xVC4+EywBCzdm8mqyrGZ5799VvzjV6Cm1sklSM95DFXga7O
ph4B24RAKgltz+XyA1wF/Ln1Pq/SwZADD2qG7QWad88V+8lX6EkgehIGjmOicAF83y1lA+/boTek
v/7sV+dvWPwnYprFQsrNB4KlfQKSdBEDioGAtYavzso8+9i/cwuN/LZpES29yDh3xMXSQbLteoTA
Et/H6dM8+ZPesSmEdR9jzr9/eYpJUVSnhYnR+Qbwd64SqZIvW5sKtUxFbj9TbmAU/U2BHsyKyiot
DQ1wZWQSK1CSiaQOlGrE8Texc6oBz+EGos7mnjrUjilQwhiLdlKZjDR/QzWns0OI554+CvNjLLUY
a6CoVx688AbktKrthptV9uzu61MiXFTmWn3ocd5F9bwA1B4ovtJmey2pFFuJ/qnq1QoWUEF30KEt
Wvv2qHn+m4Dk8wXZPqH8gS6/p4SlixXCwFglAAcB1djLnk4pHbc7KPxZswysIGcfGRZb3LkuEZuA
loyFNZsofjikiItTsRfW3yfoEjS4QyFZlMDMncn6KKBUGvkg80FmEwUK3u3kS30HG5sLQUQKEzg2
anXhp0+ny+TwmkW2DtaAxQZvA9+h0QPVyeOE4Os7ri0S8M0F+xlTRRvuGuYfvTpgXI9p4nb5uqHZ
TRJe0Rr+mFG0rrPJ1oz3AvlFhz5k4Wwnp8KNdQRtX0IXvZB8AXnbPMlJ+WWysDsLJqZ4XXoQx9ME
u5CRoA8ZUi7pNJKPEOFHRz6sLTAliK+yAj2TzQH6LqYT6ABsh8mQzfEoilb4tFLgJOcWIfe5DFpK
4ifUhr1gG2DoTZJqVB7/rBg4XjAzOGL69ZQyQdO3wnZEAoTgLQpXpEhrsm38ImmWmcQ5FdiCVUxf
RLmY64bSJMcjwuqR8OMNRmvqrFPbTGJKA7A3LU6sFv9zEnfpKj0GWBM7OBm5rDBjg+nK3axPMFjv
l+T5Qx2peFfrl9g6+6ky6v9VbZKZXBhuNZK13Yx/cjnaZC65z0nlbtlpi8cRtGjln1qx0A/QxW7R
+Q4LdfQbubE3ysiGXFXiXU5TICn/dcWu+DsCkMvZq0k28TAkFuEabE97QQsw4fIB7Sf/QQRTUBaM
qxSJHMT9HIDmtsRJoo6gggwpSaPJXzWjjKY3imyvIcQ8jvZaMzVjbvz6ld5VkdypWwGySrIcLiYs
eYNYPNHrZKWYATqGZgBsDl29dN+/7/KyfaDZGcu3uindcXadsFDHbYWiCb8gdiTlg6GBQUauEDaw
USxjm7uuIF9s8aosHfGMs/uL3zWiYvK8L4meUj+1XnU2AKrqvo/7cWSEhRAT+uCfjr1NglXqhuXr
IFK8OLaKzSrv1ZvS9hogSTij4TSzattkVnEH/C5GKvCFaJKpMVUxzsqEm+vTzEA9kBz4SqXLU/v8
GqCeoQVzftHLLDU+QslToiRFzZ3zUCmC/FmG659QV7WMxQRerG9IYLUxbrgUE5wNsLNatSbhHRmX
zF08zqjsOgL69q//vdhAXz0GMJQPERisO59K+pgBFN+Yn3Ma6WxutEm92hwuOFuWA544wAkKbs0z
DaoZMrJNCT2/rKJjhFqrDN98o/l4F0aNiQ9l0xWBStT5bNnap2+G+PLXUn8kw6bJKzVOs5R4VQ5F
GOQ5DpTHqQv9V3szVxFivFcWoCVktVA9PonF9OosyVIxemuH0zzgi1kK+2sfrTwBu0/EtS6pQsAc
94TMHTXAPMjwBThbTCUSYgcOhqsF+YbVjzKi+aV+aQ1NRbRGhDDFsfx3p8IfuJFbOKHRi+nxtuWA
dDVG+p448NDVwvmmGIXXmGuqXkyVfzEDJLQaGnhKql5YqlSziwJlHQx/ZqyElQezCcUV0YQ2NqN8
Qd3BArn4HeTpEiDkGS23mdtl4nLY0ql0m+5iISb1hAycHRRTFoTXruC5YF5oIxXLUFHo3LhOIXUQ
ruAXF14zVaS6FDtv0MjGycSiY+BbPugkADgV9AE8g+tNiMICN+DPX0z5nEvuefLTkgGtN/lyhf0y
vJftHUZoN13J+tOup/kKdVmKTxLbaT8apnv5dSwwon07/AGA4dd2dgnTkENs55IRyl6GixE/+Pyj
bTQRL6bQJb9rnPAdI+0FXLxK9pLWeozzwp1KbdW9xeYgKA7PHxsSEeKF7Ng5/Ob4DIp+lyJgUY9i
F9h/M0xPbGPuXwpC2lfOSNEs8YEH3GcGkns9v8OPojp3iv2sTP26LVbcwAZi3Yh4uatJHCc+L6Yi
h8+3UWC3AX9AjOtXFn6tBE1jzGCScNcS1LafD827kJVKCEvRNYJtgFdy3wQf3SgGzGaTzC0ctQb0
vRuoeQ5HAPvp1U4+mdU/o9qBF7PM1VovmO6Sjq12zAwWldRWTSeAqUdT2LUWLif+w5aq0K3re3xR
FZs9HCSzgEpt7HKbz1b5gJPSrsfmag8GYqCXX5/YeGx/vNq6GKNfx5AV7AtfKnkGfDhK9b+6Mpo5
SsPent4zMxZXAY8qn6WazOp6LKTGIfK+F0ivTxrfNvfVqpGh4SC4oQS+acxndWbbgZ586mUo1Yrk
0h1qFG6BLSdpD9XzTrnJZ95rjv6/ORir1zsxW3DDSdqykHNKp9tHX/EZRohfnGeX63e5YaHqZGcb
51UMMUmN5WVjE5b0qUe/NgYx1/mCKkEqIfkJ5QPrukoKDaClbceoAM3aHAzfBLzrl2fTN4KOaSkz
25lBwCvT3AB+ux0oe+eyAV9UMGnMAChEwnaPWvSswfJXy7nd4iDDWTlNs73Lbt1jrz6/X2zRtmuv
BvIWG0vARA1Z8Zvvirz9VFuytL/NC7TEFa7NhwvznGVB9sM5o6595YddH+SLZxApKpqh6l70BnJN
BHxEYY9gQ4oOh8q0TYp3Si48KdcZ2yLiHix/oJR/YxasHKOxS5y+aRwqTFTieeqCQvXI5ZX8oIFF
6sIDcJh8a/CRPEgTQT4jXTHIYRF1Z4H7ncWxuLTOiMPEiSgaIPj5m33zpAqX98yFZ5xhtGpoh9NF
95O+qocTfa4LWvJVBgrboJh6akeBGcbNujeCB5gyYDoYOeN2yuDtXr63yM0EQFWFIy+eBFLo6p1I
QQM2h/9ZY1PHfg/JpS5yqxzkq9qcyo+YVasO+PDPBU2f+3wA8D6iKp6gFSzqxPLx4TjLUB4l78nW
fzjDAhRSEETUPsmt/CR648/V364n9Yctplm3ZkcTle2n3TyF/k3R84oFhXBRP/AK7kOy7IM1zJJI
APPpzBLJU7a89o5e0lJlxsvMUz/aRDVxCNy2zjGx8B1t4BRh10tVbqPgh8sq3GWeY5pCOnKts9G2
yX+xyuxrcSNwF31Hs7fC5Zr77V28Ss/pPnnGqQV1hbhPZx1u8m46w78Vt6O2SUlTl45NCEPfAgEh
DSxAhbsfjlgPXQdgWJRBGejACyDIYobBNWXtvL7zA6g2k5UG5EeuC2cRozHpjABASY0NNyZv3JOZ
mCGK8RykdWIQ0pvt82bGmYDlnYn9TtmO73FcsXse209ClWXNTph9WFhq0ztMaJWlaBbViTwxjrD6
cVLx9l5zH3JG6KSf3rnYRwbwLDwtZpcCD6YfDEbbU31FxVrklJ4RM9R00ztCRzVrQjxqK8To3CYt
NV/Yybma6gUjrZ1iQLJjp7Z10r9zJvHNJ5niFDwld3YrKNBWYM0o3Ly1rY4qMcSLgpvhiEG0RHWs
/MtFGa1irZvJM4D16kBbsSH+0qzTp+XP7unhc/Iht/R3vXQSj00yG7H2z0w+KyyRmkypxsv0QmLy
fgjTEgFfCWLaTS16izL32fOO7ag8jw4r472pKDgh/0Dq30+jEcnKeAruy5Q4IePs4+ISi0eVa96t
cq+yfM729pzQRC6cYuTqh9fCDLyK2tVkprdf2BJZ2NIv81cx8mvdLR3SDwCUJL45tJ0Pl3aGpuZk
lQPEUf3fGE3G0zZ6wsGkLb2YezkX3Kl5L0jbwXeQZwStVyrUmWMZjRGtUpqVE+TlD23DNHjUlR33
JnKDHs+jSlDTwaQFMmJqt4w5l6QmCCE3G2qGAcVaicV7BbnsinvftSsvNsqRBc9U7q/kpq3FFEPa
KrCXCzE1amDSFbloJ+aNItBlbUL7rbHz8XTYDONJnZCGhz1iIULqg6dYYT/keaTj/6QZYpmBLW/i
GRu7lbPKHzXB6WC7sJRpTi2H5QlZI9cVdkM9Yp2g/ByPzrlYaHNZktwKqRgKrVKF3Y126rKiXZrP
XfEKw96ov0AtSsiisFeWvdu8uSym3ssXucIRE9lcD8LchadYJoVV/5ApvGPffr9wqpzTu44m8Rat
MV9TT75IMsZntaTng/mTuw/9/nC8GGW0qx07Pni60pNrs0MI6sMR5bKQ7vLqw9bD7GyPVHs4ZQGR
yT7U0lUzu7gj0ILuRD8eaciTTubQcBFg7lHYH52xej5x3aAc9eVcrj+3dtih/zWeBShm37meInPd
xF1y+XkUgQSOuHeVzwDuqgQAr3OtCr2nx3wT/m7eaAYVwlVArHbdUPSv3qmMwb/LEuqpZdD0+C4f
6ytu18IjBrxqA3AUEe1VH6cfjeytUTK1bgOPTsoOJbK2ccKxDvo+/lFqEOdZEjXdmdTOa54VnoX1
vWdtX9tjyQa+Ykl6iutlQWh8V+rD6I/sgL+HSD2juVBscQaRS6B5uFQ6fN9r1U9e2lkm+8sga0+h
nvQcq0nk+dqPo6rsDL6ar0ptOEUY8tLDdsaQRTk1PGktMNTNGd8NSDLDvlG66N7CYULqbJ7c6o/z
AihGijxPBiNFcwRZ5hl7ouktnKTlD/5EqtL4uhvwq6RAwVsUC281CYvN9gDWVystIknQmLGL2mHJ
zPvzfkJDpIhrR3zKU7ZcK3XViHNQvWmShT04aFrQrV8Z3kauLPlR3U8pDPpnFO4F8Px0GZXUJbYx
bXdI7MoVqKep1l5uQfeYWr4tz7qYysxHiXmshnD2eMGdEbgBDZmt2TfbjiLFNM1XDVgu23vb5/7T
L0Q2KAiamlHoSCVhZLrFrAuGIMLAldsVpv0RHaoC062m7xdP+EcBmZOxLOw5K4Zl0mMGncAXWMLI
NfL7/saRTlEOaG/XD2SNdwtj+t0zm9vf7vUiau6fRlfOtCh6gd9+H8DAKPD7RotzNY1ANUFvhmiP
VPbT16Il+sWiXk2meoKrvA/H9PBTIxV0vYL1ttYDu+WeL9gb7tSnVlanc463ryOmxcjtwfhgi7nC
ToUS37DehougkcUbtRa69DYuWHrKgPtSe0rF3l7gSfgrPHe0DDW7UrQWDcmwpsdYB9TJXKnPNip6
Q3gxBJmUOJ0yNE1dwW8IQm4jCNhNvcYV69k7kSXzrMu5hutdcX4mQob+tdpDTnhIylAPQmOzouMS
YpS/nQ5lLtFyuD/hqR1HTmzDyeNAC+ySkHcv875tiTHD9dc+XnfX3+Ivpq33mM6ln1Nw/n0ZOgcD
RBk8bjlLh30a/WTd/eDGN5w+OHw9IvluShieQfUo5c+p1l72maRRt+r0BII1g0VqhX/MYW0KeqY8
AGwAEdaoAEACiTv9S5SflcyngjoiS0cV3FpeudKWM+VlCO4KGwTxMNDd7+VZaD+0WSIhd06Z8LCw
r1uDmofyR1rLC8bJmPNuLuaZBDak/9Juyz/1mg94aablKhRdA5hbooi8UazNTRQAbhErUerUMH5L
8D9/KJc9FtO2ZNSCDCUYQQf9yRbUy81g98ZSkjY2CwiL8XSROe9O0IqjBV8woMqXIckrmapg4evz
cw+HcGxjW8WdHTZwMlIl+Y1BCjf5nmLtLZogI9UgBLuw79RiTfUBovSrTfgURn8XGZiAMqZIywzT
qgcyilUQ6YwD10C3Of8yrPIUxm9MjDc6+Dr5PSYE5j6O6TTIuVz9oq3JZfro5MAKb+SVpx/iqWW5
swjw32DKQLv/SKtvLuhgN7+eQxO0dF8QaYiFmIDh0kUp+1LDBufWmXW6RoUMsS3YOoCOVl2DpZzy
1Qr+tr0V65WJAR7V9bHdFpb7jxkmz5OIiCC90Zr6rSXkYaPmFT+VwK6iSxe++b06I9/ThsFQO6Mp
HTd5/FjSbttCt7+MvKA0F5IYExrimuDnjx/lZ4V520GpbtgRrZDEsgLpKWsrxjozvn0bymbz4VmY
kigZVQ5oFhdF57zDU55xacxgR3IM1JI8CTG343AngX6OOC3qVY4rduX9f84cEeZgKIFK7FqcWXhP
N0wZyTfdCeoLX5Ci28U/jNhoLzXtiVen57EZvDLpG6AzxcDV0OgyU8gD02eYOqWW+AGt1b8awpyA
XmVj6+m/p/7ISjicCf6gG3ZJ1KoNFFQcFrsoxfAz1JEhqS19zPgAxBOTHyF/NVo5GjWrJagKzAkz
UUkqQHA8x6BPjKRjPkcv9hFCwxNonzyHMu1p8giVy1Mj1pskkw9nPYT+wGTcYVSogaw004qxOCaf
tlPHn2mETGxr7Ah+pbNZE7hb02cR+ZceIU7GTybj09o4H1OreLbgUlXnMPwfCf9G093i/4D1uY++
3n18+VE9h6Eie8xE2wYwxg4VvHsHagkuq3DT+vUc2wtBjXiTv8TElWt1mft5tSvwP1WqKzY/PBAX
OwK0K/Z5I08iyIyb/eaODPITLGKwqfIikXyVZKp7y4p6AKsQq+gE302jGH4pMHWH3wcQqtKpasUo
JlKEMfUjU/m1XXF0owSVhg4NwODURIfSaBpNdKoZEdn8zYp9H0+LqisItnxXQNsBiTBTiS3RUkg/
0EfMZzpU1pTE+VFO5wFpsBZNG9eKbSKST5MnLC0wJpF03uWUU/ekzGWgfILFs8+cMqFDzRYq/hoH
FS6hHzygWWmrVYEauA3WfFjSbJ2QNsD4mDsNDcj7xLkWcXimQvuhJcTUNPkTO9rR50LwP/98Asm1
vVAuUUkCAEFaOxoY3MeS0dgtIrfOUBF2ykqAGLrtORBxI3/p15ljSnkGRcyw1r7qZbIykMWextd+
RrDNWeBh2r3/8lYJruJvbP4fk5zD+8qCgMinclVe3TnOiFdapGc544TvAvV9dULYTzLY61Zd94l1
JUhpLorcGs9K0KWXKWAnHa6KdRrjekGX0ACHwlklAuIbyjHH55ZnnGcL4q8gArkR2wieZp3irsfW
xcUfsOiZiYZr9UFdud34V0Fzyd3l0u+0fi1qex1cggbgd4lMPwCpaTvIBuXMAPaGswK42NTNIczd
/q7MO/M8AD0/yVZp7OKrZ1yotWvBcJCloTuvIQ1X7vYyheSvj0EapSlHUOxnLogtfa3B1EGSJtcB
QiU9YFA5eG96BEXkNbXRVfz9wMjx9sK1+nLB+juIju1PfjLanfj+Mrkh+iPKuteD+O5Vdfgjvq49
QjdFQv/KpuriU192seOI8G9x5uOKsbRE4r9V+k9GpaZdJtnrTb1fj42oqnKDQ3VpUIv7EihlO1vG
BBJbMfEX2LXE6B9durQgXg99NDiZi8B4bbO+Nav1U1enFR2dBbFHMoTX94VT7T8HG6oraEDtsfQ7
Oj25dnuBAM8AqipuwX3lSf2xAIC+Fsyaj8pBlmI3reziqTxguNqXVJBZpqLvz28NIn7vigsrQMEG
4cbLutTurv6mvpQNKN49dRZQWawBEAquCLBZpmWcwj6Bu+XKisM0kx8Iws1B+90p5VV9oLsPsT6M
RtUr8kW9OzSIvER/VzpG5y6TAPJHZUW90/Maxozur09varYMwu6a+w+UvCcPbrinkum8gEx2fLGE
toX7wdvmnlwY/xH/NXSJbr+tYBskMzx4jl+IVALi2gCfauhdp4kIwYgj0Fs9rjBx7uFTwrnYncdS
DSnb4J6UDJUjp+roSZD7xMIfXmDAhiTnYIcWxqow+17pqkg8c4LsQ0fwkmz2/jZc5qS1pCVqUDks
wfGhKQBiM8qQpECnToppm9BVg3BkzahzxZrXmfVnW50765bVhc6OAzBtAMTPfucd67ISu5GY8uWu
dup5u9D51BpJ7VMiVDJE0BUcpm+q2akMrWbXuIpn4i/MyQPIrHymHfG/Ak9Nd7MvA3p/A61c7cN/
p3tTkliF4N1BN2PtCBf3yJX243b0luU0P8eJOy8cZQ10VarsgzlypJ63Mwzl18nP+AmVMkV56N7y
PUJShsx+QTSsWe5vWDWkE5aVMCeY3NyeJAKKF+7ZGiWuVsdXRKUYBL5S/NX/Hf96xlYH3r1wX7qw
+XObXYde2eOzhC+DCfRfAJNFFZAL7YNN1EKxfRRY7ThKR1VIAu8v36mua3FAFJ3jZRYxJtgRsRV1
DnPLzMsZTjEA7Ae4iexHpeuxKK73to8u95PqfAcEXaDM/9+HV2sGj/YB7MDFhGyR0ax0dG8ObkkH
3OAm/TRiS2eDY/+U5HE6krkd6sEGZMQBw899SkgypgGUtMmJb/KOFK/+jDO/feAKBqFisjjpcsop
IqFUkeFgd47nLgWtNOuFnkr3EVFldBMEu8XvLnirhlFhp8aJKyfx3xZdZX7d8h1kOyst/dLSZrgM
O+/qKPuo9R5QX1FG+6fFe8S1AX/BFXPzKxS/N//XC+U0iYVcKfoKms33A0zUm1p+1wLTCmnn4NKv
Pxiwxc5KbtSCu2pIlOB4RY1JprLLGMAGi2X/ko/+cKkx2oBRq3g+u3B3OZetBnB4MpE4toZ0tymZ
57HEWoCb5A0L6zAkY1UbDLin9dxr9VA60q+YZAv+qE1W33LKEAgvCKwXoyO0b7Cyw1Rhf6Mn482g
17e/aB4rUKIKwhXanqraG5/VsT0Ul40P3fX5uxgBZ5muuiMizWB1fXpjJWEtQNpz14ObcAjl9B40
ypODF3+85c0W087bdOm21J1B0FBaVkeC0x0KOttSQ5ceVQdHgHKN2bNY1KCQGorwYZjgXy0ia/6z
vj2p2HJpO3OcaeHoPXnWY9h8jqGPiNX/f0RRpeVg1ri+H2plYxhMgaVk1H1E4jtHozzEBSd+FPmG
o9mkC7BefcJj5XSV+5v09qe7+CMFJEnGXcRz6Xr2QbzrtpSSRcEnWjzsHz8pjU8QPMhpu4iRSyAu
CmPSm2SAxZ2B5+ILT6sm+jlLlp0mQzwz3sY+NDdcx2d1SJ3ZdWQq6B9SHJfL3+xl+8m/11QlA4Ia
fSmgAwp9FUsIajRDiDK+mH2XoOD2glX3LQRaMfN3lo3+luFVFOrM/n/+6AKMu+jEaZtO+LCd7Cfl
D81wk+vKzaxrwobRh5D6W1Jd5UnBkzGYiYOdTGOXFZlWwMoY7RmEjY/S0xnT194iAXz+QDO7QnyW
dMl9CECEwEs1RLkKDHYewNc4d9rxUX73czoWLtj0IeZ38A8/cd8dLuh4A1LlFvg/EgWWXVKJgJGe
fcNxaFfSHJ/1CN+YPORv6HQHS+pWPWjDtNKmaMTyJK4xIYgITFg7xfa9yQ1vc+E/adAlt57lx6FJ
zdiDBK1UIRwKtbZ9cXAD4DmExxoC6L37G6RlaSW8i6h0QeyBXXfY2HaMxPr2b2wKBRt9rhbXkHJ3
D+YAA2f0Dt+9Mr6J9q8tkWTDP0zH/GhImue+rh5bLxBANF9aDtjcadU7lFazeXJZsLy2IUCuWOsH
1/kHm7dllRPrTXd6fOii1nvQN33y0XpEBzYd/Q6RdSv5ZWH04Lp2uwkIEIcPhtbw8IUSccbWjgqF
qHtgSfkntxyQxaz1w171dfOCyxwyCh4agezeyS/ktgH7T59JIPaoLGgwEvraDxQc/rv8pu4VG9FG
vn8pHbNecN5HHexEtJZ7LmPzFQHzl90uANE333tEL5pGppB5D56UPiX2yflIDQVMLClroz8irfXy
Q1sDeMa/LGO0CRASgedxSLGXveUoXCoYVWE+e59NW9NVbQMLpZ0q/3ljEsrAK28dYgKxbPkGfjvv
0p1xdwY/5s05Di6bf+znDjaZ/pR5nnh+gCkEUagpEq9STlQN413neiXEDM1W0zBiWbYvekLN06RY
ByPdqsoJLKr+ehacPpAh/lCIpGjGoPjsomls2cL/DLqr44sux/By6sxcrUsMtJDcql+OAquUIkQL
bnqX/xw61ywYwC4cJZH2GNysq0bEu4hJGFnXz1wKyTXV94lXyqyoSJgip9TFIG19d9wocS8v59Mu
darCsdWOLww4I6wYmy5Sil0wC4YO7aeqn5QAhb35uVhcYj2DSpNMZctAZB1qcgDK+SEAiV/dKxe6
HsXIiwTn1Zh+QSA3doC5/coD1BBn6eCHyM35mgQZN/iOT6YX/HIpyYx6+eN4QAMUDchn7vHyjQyZ
ZnbXIR2WdBJyYipbtm70vZ0WH82BGtUf0EPxN0z2inS0cuQVqZQ4cf4CgEkJSveVYgj/FOOX5QQf
IzWOYJG0S9OHZt5ou8f9MHslCrUGX+wHTx6QqT51UB3inZ0bZp/iAUPovmfyoi1MF4fytmJSQtjF
GAsiQrQJ1PI+EiGZrYgxBl5rUdwkGcE6bTySZkJkb1oRyj6UbsGSGWvqVEFF7+YpN++I7QAoYw2d
zLYPjst70Lol0NYEcmu+u1w2/5CY+eBww8qCn5QJUpx2Xkqk2YUZ22Cro543lQeDLJivgnwFmcfo
Z2RfAFKcbGGsBFZ3iydYNr0qPoFbVf491SVEAS+qizN5BEoDcbKSaAicS3tjvj+ru8w75ymiNPHP
a1Hzd1KQtcGSnVZ9d8Mr5MJsiSR/zZy6IUCMfYIH5lJ2x5Vnw/0HrHfFuKlr3LSINtKt99rIApb9
/NDWyp6Ju94yG7gcPrJBCm2oMj5FK64DEg8KhiLgjO8gYC1aM9ce2ybH5sO3Uhdy2QejFyb26OB0
ZY2tX5+iicE/hhrTqU1Cigr69MKDsPxhxeq1yHNautU1MfGHvaL+ocB7fgqdzEoLclS4A7P93orl
ff4BLopDAuQGDmSX844GU0iACPVmsWdbsEz1x2YKd1J9Vb5IUEn0hs3xGFyD5Y0C1KgFuWupef6r
6/ufvM5miVn83w5fQiIroSbvVNfDuuDsgfPRYwi1siYB/niNYXwcwBzbHlAha10ddvcT1xnZQ/EW
uUtHVcO2UrUKYqWVC6xi5KlkO1kB6ekoob8iQni0TW5cILmdMoR5fYhcqQIdR1nXpp7XBY5O/IR4
0JoWkcO+wEsK44Oet5bYrIC3umucR02OvHDRNR84nr7kObmpCQnOqliIUATM2U27e6bH2uoVvhue
h4grNGgqrdSd32y3PwRxnsJFjY55aVF5k7lizkRupgSceAyC15yThaUopg0o3S+AHiY8qiuKTDsE
U0tmLSUmHrKODGqjruIiLUm4FJdDfGAFIV2Io/UnUfqgvqbZbh6kqpiztvGtqDZ/xBErGp5e6Rjw
WX549W0nU7E+8Txjs8DWJERflquzzANGP4OJ7wgqZBQnKl3KkWupda1fAJD0WSlcY+/NiytfLdRt
YD5tnlVdxObXBYuweYtC6WlL3RDMpy4dx1zmoBJXj+TkrNFPzxxZD2n1NszV+ghOOhBEBni0xLSm
SuIVQige6nCZopJN7/bNoQXAst1uki5+OJ3MbROo2aJnPElEugQS7RuybXofONAst4PJwrOps7BB
FLVxQ5hHdwWXZuFnnGpwFmmpzUzZsHrCWUL214uJnHU3dTRconppDo0UuOacV8RLUJGE7lUPGLgx
PvxCLjFMINwZ1xtX/UjpFvNyTExli92/n7ZrzuxrTCzq/WXZx8ae1qRiZQ62Cwo08OPkqugM7aqY
cVmtpOEQganbT3eIYh5y7KCRvxnftUdAuoql2k3a3Lp6EIkLGjLJpk4l3hSeiNA2vbVDYG/Xkmlf
kjzkkqwyLQdQt5m+Jc0xPJWAI8rQoh94RyoUnavpGIn96YrJAcbQ9vbDpKnMK6pS1+OkcTAKek6u
zT/H/DK9s3MPMV/nM0FkACeMIKDrasqAzBjdUthS94Q+l7bXp/orW5iVBLqjITBcnLQE3mFgT7nM
q2wBgW5yj0UqlJri2ugRTgeh17Dkn7/xcIh5AE61jPegDisrnSNnOEv1zVwlcxRY5P9hoVAmf6Kg
Ixsd3enBortGow+7OyS/DBbDPEYJMx/TpwL8/1g1gIOxlBD8uxbC7fNLILLGM0YFdSYQk9B+iBq7
mcaIyWx+Df9gsEDBIVLLfa2aSE7X0cXoGTTuWyyhs+7hSKQNKydmAS8sYGzphiB0V9bOCYBFernM
sXiHUZ3pxohYFgjPfwiiPuK2jzlNmvo0vOIGxfE6aPULmrWZ//CzYsNrZASJpAL+P/ZzSu5MeSVS
uvLPF/VpUUqAChMneyxXQfX/mRo6+0kiT/EgityLKqL+kuOZrj7dHCSKQSfJ8jL/8YJNwX6tYWLf
XwfX3d7Plwhmyq7JBHozPPnbZbYKan6ql/dBtrEXCiDxxw7Z4HgH59z+L2lPJJAA4GBnCoZUIBSL
35X47106GJC0nwq/DqDXUMYhRd5V7sHvgi3yl3zf0ZmkdWh5IY9i31JOKyh7+VQ2E/8vct/rH77O
5+BmgThpuimmP7JK0uHPiYpFHrIIcQx3gNArJHstm4pdTt/OCaBQIYWPey5/GllyhsV1faykusVw
d3nJE39gf3/OqpwxbjbX3mqYSddnK49nA/wtQ/CPQjAV23tFjAX8t3vTCmhAYBdQVFubm46n5MV9
bci1OhPDaCwZyuq9gIzYsAnzkH7o44LWLfPxxWAsNekFDOAJiK9/Gs+E6iznmmgY/0+OnircukzF
nXlbmPN4dw8y494TaRZyx2bZo/m1i76qjc67scKaPgkxC4zJ3A4vF5cku7iFEIzHp3g6B1PYawmi
B3IVjV+dejMF7YEseuQJX4JZTS0NlCyyax3AWU3cfmjOy/UYVOcapuJPpxLLFrRrbBrhJSsTinLQ
j+zpz84CGeQE5BxeMQnlfg0v0yD6qAoKcdJqPEonTUrDSaGUTjSvWdMH++GnhNDgGSFIhRe2Kec9
x3WUJh/FiunJU3eDRQxcw+9AOy+gZYWvPdBMR4nFu5o7CkjLXTyNIO9t0x1S7Ecm8ntK/k8GswjG
7xDOaplCYrDIKXnMCj9b61obMIRgwxlMf22qT4x7/nYdYG4nKBY9CrDusxzNii6jCCq+jRJcthVO
BWhnzEr4kxbeREaqN24mFGbJ6Cli4F8SeLMikRVQ0G3bQ4MVSLr7hhp4oiUq+y5qjGPOcqHl03XW
iSZsMsndDgbsKBp17Vx6+c65sKRNOo3uwxJL9RIi38q/QpRxLAJHyzhfV3BazPwydVxZNl9Q0jKp
VS6kPieOhiPPk+LfD6++UoCm4geHvXite2sRxXSheD3BgoIBHj+4YzMNc9wHUjpnp9sJ6W5wtL2c
A33vnaJKma/RmGr5n01iA3f3sDeqQEc9xMeuWB2YUw18uCzdsSjPxTnTujafVzFEAOPcu/tTyVW5
mU6VvToZRS+6Oq+K/k+25XoaQIEsFYQ2fz3PoOkc6WUtgGBnJtBuV9iBz0REd4ltDiQQv7EeC0rx
F3CYNtr3MN9a0EDb0KKkBsXLvU2t515fTbK6KPmJy5jcoS9sk98P1nIHy/uo9ZTHPahJJwdpiaA0
os018TQvK5DPPCtKyky2H1qplbW7bciUChGKOaQO9jMFwf9JncMe5Up/6mQWLgS2plVGdoYPLTSt
7WWvF7UcOAqPqdrFg+9Yo/eQ0rKfLI4rJ0jYM+hJJpo/bX6tZcpMcYJwSJR3XHWcerMKsHPW9DIk
pG0EM5PYMt9bqGMlbr0Z6/HzVcaxzO4NCzjeuH2/9pUHZEz5+zNjF7qDqLfbSZ/pKVrx93RabMYE
+c+dF4DLiVuVsnPUpo5h36UMejjpbda9h/lLFl0kuAQHrTFeHcVwQFsPLR+zcHLynBa0ZiiiHRAJ
c/Vcns1LBM2xytA0weTPw4VjDj94pOV0zgpYEO6hGhFhizRzO3ms/NkMpF1S64T6w7uWF31zR9+/
hvqkGxy1g8DQ/6ahjShtsc99y15dLPhQQ5kOypJIIW1grHPADJyr9UIbIphyjJIq9GqtYP0zOF1e
IyhoBBoLIcWXYC/ToQCLSijXBYK76TiRuYvcEjLWDFYT+hjzTDWMJUV/zISaZ+P5hFm8OX7nrAqS
oKghVeLo2l22oXMnHfw59aaEC87y4jydhOrfWEerYw5DUwi+PTZGl6jJWGQwcD/ipa+L6d1vOfu+
NsjymlzgeoQextvcKdRCEx0MH6YpEvx2R35O1dHDu1s5uHlL+5wBAZQHK7uQvU7oi+C20Pzl/leA
FOUPiDRFcIz9ogbLXerR72IsofsVChwKzuM75bh+F0I979iGnZa0gjUEmySj0NtAhn/Tlmcw+aoq
xRkbfbW0oOsTNz+xMH5yLo5m/HLUJmBNEl5RFLXlHC0M2RiCuWNJW7LgJNhrn1sjSTAhFMo9eDz0
yVnue4AtbgEr20LWdc//PKHmfXNGKMcFjA2Q6c+6bSOPzZn8BW3clOMJKzzgMe/KQiYHo2z/MQx2
fQDn9S7rOP2qEJn1FC0ZKJW9UZbQuoA9bznlzL+PAS7kE5GQbOxkjtD6KkI+UJ9QoliR0T0RTCpE
tBXHeSx4LFcZaK3cJQcDcDhD4Eh/FqAEa5VbAsC3KH6H0OMMcNuGN8dgOUArxnu2y/OzXwdllqzl
v7TjWTuOKwznIqCLrWRw2UUDbe8xTvzWoE1Qk8Y86U7gtPlY86Ud518+M9H0xkyaaaAxC4UbGKxV
wtlMLCQ8tpUfMpMOb4/Lk/p139vWweEE/l1swFzi3AF6SAZrzF6cI5pus3TkWKw8CshT/El6hj8y
yEn/s2nFOHz/aI02qjfsolxJ8j1cH60Phr7I2JFX+nlwmIH5RN6pGDqaJUrWvwr0QLATbrrvDyCq
jUXCRsUb6hEDgRrb+BnSub0eFiRwUWfIbBM/GRRUGZTTpnxmB3jpFnTpefWTRL1A74Ax+6nSEEPL
MUqEWI35EZIro9LBpRDyanSObnbDxrugUbuj9L2QX4K+Mz3FCjut/SZqlFrLFaw71djCK31UogzG
9QfM3+BO8wacVJox1TvtiB+4uAs1Qf4FceEQkSv2lqbzbL9XMHOFImtRPtGStFse/NiBZuKsRRXJ
ccUyoZrcc8t3V/68xZo6rLldiiTTfJsx/NE4PzhEOkUeWrQD/O9rDxMnS7oVaVm42vWpGhIywg4r
sZZYJiBtwRkH6w7envxHPnnE/bqTliIB2RyFa0xdUdBJ4a0dG2/gOzpzkeir8tsVXR/oMkK8EU71
bZvFC9p8Gy6jg4duljDDcdMQ2nwEWfumk0OMblPw0auNNfTjqoqMn+twtO+CZzMKk3ukhm5NTvCk
/ClIJIag2H3B+5EvnrlRIXKzhKal1IBUZEtuyGNi82iXRrquHyyXBNB/q1vVbR56hOFQ6Uvvoc2Q
gZuz1fpZKDiV3UUToye0iHBcW0mJSfnxBm5lAuDNC0TK0p3I8YoBZ2AvoRUG/s/2qtkDtnBa4DiJ
ISnWOLEsabiFrZcPlmguYedL1yHHUWu96dSUlVsQvQ0AEb6b8ZosKKzVYGw6Oco4KdPX/gn6wJBX
SVTBvGXhTk9dyATITTHfKvAANoWcCetdXMjU3wpbb5AoXjJNtP9VQylwUN2+2pCet0G52r+XFR4Y
n6zqH9/NOejJmmh60yNq8chqPMZ9H51M8U1ol3vF4dfPopWpMosRKcZl0pbJl2vzUTKJHmP2XHKU
eRpxffGeM8rANxxVW2YHPCUYCHC8sJHDyRj0Cv6b5O3f03ekt9rMw2hZYJWmaXVubn3evjrx7+Lo
/8ZcyRSfokEdzCLA/JDRNtf46W31PPrdUdr2L4xA4zfUTxk2n6FhRKKk8yBuPR1S10IOZ4mjpa3s
gxzTYke2Z8uTvw6vumCc3rmUNnhRvLjpXqce8evpcUAuRK2X9utEs6LNgNpsItCrH4mvIyL05/Mq
eZemoiXVZ4meFF0SeOZ47e+AQ1JSbgiOcH4EHB3I3y6Uot/VlGFoICcPcpQ9jUjD2vzGrSMSXXgO
R5eupelFkWlyS7QVQcMO6melKt1iQ3beXa75tgWqlfA8ZiOCKqpJyOpaENIQ3yjhra/5Ze6yu7+D
eR6nxVjVW6ldgYkvdjmibEQyTI+I1ftdBKoCiaS15dokw4kQgYpwZDer74BxzUkQyzgnGOnIZJLX
37HiPpwK8aIdJa40wsg7UWRqrHSL6n1d6M2xqnUAYwRKlv3qn3XcodWiJU5E+e1cF76UKEC/rSWc
LLYtZFko+rP+0ECQeXsEDLhWjxX3t7pOuuUdSx0R6LQkaVnoSKhoMVhrZ4QmUfvIdH5/Pj7clpC2
Y0i/x6ajYXy6EoluS/eNnC9GRuIHY+WCCAym2eaq9nR//PKvYTVvSGFzzcZ/3LZqcqVigiQ+qRft
9gGM+F7vqnej03n7fG2a2EKat25Uy5QUOKXOvFMWzHVLZJa5cdc5LEginyCImfnDr79ENGiERvIF
PZHq+vbK9YMu2W52ahaufVGYiOx3O3oxE4BcqVn9rHwcDokTLJEYRRZqH66L3HbogoZce7mOzqKe
AEVO0qBJwmwe3rD5UlJLfwcUNmMnQoyTAvohBBYJ8RqM3aqHHbAO3lP49Y7Gx9jwobcxAyPUxxGY
/4c/XU9a6lxzTdlItmMIyhzwV7fr5ASAeMVq8NiEVrAzbuskhQU4zJaarxUuDxMjg9BvRCbYgaDJ
0wG4hWdX4JvsYB/jZ1gzys/PFtBWHBRUtbjZVzBUFmatoKLBqgUAKfHv8HpRBlSUhDVvMsV2UE/S
4B2Ea6sSBAn5I/NvqvMxPeA0RubTFh5OsTRLzdCj/yFGCtlGtwWrrsrwMwxtzPzDEH5Aw+l75sli
pIATu8yAzqUEst/pXnHFeGtY6Z7nks1B0xnJSohJZurTuni1ylRMLUwln9ZneZINU+mTejG+0UkX
8zJv0UwnyZQASEQBp1UfLOk+SaV2FtPE0Dar9hoFKYwg/Zl/7KqvmfADIUN+5VjfY6OtqeAmKsfl
SacCOUs56lfuH2nk8FEaQpz9G1ZqUbq2dwrC7txT1S9O2HAMf/wXxszmmVv+SUMs1x1BnpFyx3wB
8o8nOCuZXlXlZRLsAozdD+vuCKXhSXCVxkXSyd5xmmiwfwc/noJVO1N6IM0QunzJomdfrkGd8MMj
ZXWB1fBEj7rlmbGQJ1pvkQChIN9EEZHMjHl2odj+H4G9Y0lsvqZ/XyhcwRbUQD5sfbrdjW6SZ+L6
1yUoLb9T2yRT6br1EsWHZY8uFu1gvFAnEqsZQxpMgNFRTpc9s5rmk5LTghWFUTXtvxh+KGtgUm6b
c0HBTJIkQ5S+jyZZm7Ltc3V+bBGnLHyeyyCbih8Q0HVDkmOqEaGVAFH2EPwHMtyVG6pI0w15HkTa
RdLefsaVhtNfAk5pdamUoVWC4pfR6weH5XPq06gUiqXT1vzQ1F+0AZDBnjlOPyhhlGQ2HpWr5/Rr
k4x3m6WhvGuW8+NXh8tFKiXJU+9jHLQvS/XOeqHRt1MYbxVJ+pm6Wx5zp+rMqiE1dwU1u5cFGqsn
iRriwMEhBxUrnG+eooSrWoR4/wnyl9k5wMWtFq3jW6KRNdF3sjMbsqXL3l7XLbkIKRAgfoyblB+t
1pKuZp5ySCUy3wPpE74usqxl5bu4z+CJglb3gXmeADneRKkxWR5JgizcoDY1wKWrOELeQNr6qOfk
4jF1pDlPBbRJSPwqigCAPQQkxEqIRT19mOczSGYolVpvo0Nj1SysWv5eDpXnKfE/rLVrthbdm4qA
HaSIOL1sa1cNVEzuCA5KYgxP6FcKn9gQbcQo65qFtYrcGnHuRCMzHruCShMt3Bki8s5O2cbikBn/
GWTIiNLdh8GCFdBjPC3BEI1OMtfX91N/FXdgR4FOnNn/k44luqZyWSctvfQc/Bev7t6r0SSIudGe
RTxj/fezV2czYZWi9fAlZwZNmau9BPWTpXVk9qsqAkj+TIt5SHa0JEnYapcz39c066pEhGx5kjaI
O6LUeh/PhUIAGnShk50Mpc0aXYrDH0WpSrFbOUVEFZ8jr3fPtulrLE/SQ1spQgh9Z6Jyolw/JskB
oXm0LITj8bsIZf3qzOa5mIYiXsfAnp1Op0AcbcAJiwTJD78j3TFTyOLRKFuUaAIwu3zRpPFCOZ8v
1qf5jwuTcqlTQdoA1SdA1W6M1h0rM9BR81eTGWsRdl+PzmgOHJ/xjuOM8c5VZ5e94ZSBKFyOOdSZ
oE4RfD1Z7niDuEEFdHIsZ4NwJvcW6rJ1lcLowsjkctLiOCvS/5fh5Er0y2ND/S87fXhxDNAo/nTi
yaa942d7WcCvI8En071mJr2Nv0dLPTo391ID/GPflIBxCekSFh0iKMUKB3twK58GTfG3UAH2G/SG
HVEdR8Le4onvu93x7Z7pa2Q+GnScJylJ5s40oT91GjrpyxVOSqEFIgvUC1jm4I7Mq2ACQMne9eck
SYy7Axlvyfili+lqbvH7RoB1Kf4dxuw5bn87XDoxYla/oX0znPVo0dK+e9mKbDrvy6yz4gBCOL7y
i0V+5NzZT7eHdkoVkMV8Gngtq6D8rwGDvFdv/GIbrHPZhUA+bHdUAhJAb+KgJxTEf6BT/WWddbeL
DjK6FfD91Fw65hUdsG5768hbaCu4VpgnxcUInX/ZPV+uIobYYamMnwxqAL2mLm1wcvA/8X1TM6Aj
9OeX9xOy8CoQNhdmfP3Oa+k6C29go2f1jS+1iaonJGVRN2x6yirfk3I0XelpVDHCidPLRsPaLF4M
/BIWpB1xz1CkULzfhwP+zuLYxK9BeFjBmA9hbB8q4G8VpwjXR/dR0FRGXCZ00ysNiPqTY28yOOTX
9t2cH8QPWdp8m5aI7wpO+XMoCfW72ME2+TzQbQNF5/jvUUaYpVBaEt6m1fy20ANrDF0EzDoOxqfb
VHhTKIRe6HJQphtne+QY7ZKLxxncZYuLqcM8xWwfaHDdIvA/tzr6CRclehWODa62G06wNg2yrdWr
231YW4NMdapwLC8ohhqbqQvEy6ioElQ+2lQekBz2G4MmBMyedMrrN/GACrvFuuzk+/Bm/+TKbJG7
MN4SreKAEsi3y50XNBordTvYgZLjFy/m7MvPJ8/aCFdsCRj3qUgqMsrc45KOl38rJK4Mkpy8Hs95
hjik9LRjXYlBN4juKC4o1hZrnqOCPV26FlVnCmZD5PyS5UINbzv2ohi+uPt1rgNavUDoBQw/ux3F
8Z8LJ8eqijEU8m0d18Rxld6bqUBcvNRBSGZwg/Wui7dSBi4RxmzXMKROeNmlUpfZm0wkdsPvJZjs
wAvbeUYzUSWrKQn91WOH7MFVvTjbjGku3d7pgKKW6ewRrdK74/QDqXPDlYloYFs0jWJN0bAPGMkG
Ba8TQJt56kXzuc1CvIrEHC3I2EEThT09NzJ6Fus/yNZtejoTEQKWnlt3xYdkLCY3FVIlJnuyp4i5
blbSFIZhd/twDo2BeHeRQuajRINnyr9TIQrgs9uNcXX3zKmbeY9fAy27dKREMEXwc8u32JrvISb1
Wu4S7Wyq0q7nrrkndsTwcNYM2aidyJfsgiQwU29hjMQ3ZcjCj4NshBzPQlAULEFm4G9eyVMdaWcZ
dftDpKm34F76IzheB3Dk/KPRimIrjl2c0nMEstzRI83vhGKahsnoeBt1nuc0vTAF3BSWBUNEnbTB
yiYqMdd1d5DH/PBCyERt/W/VoCH6Am90Ymgxa/ydRX6xh2VRbMhr15Mhb3fKpO5WUuTlc1m7cJ0D
HuhvTHV7n2LDQM4QAuuH9JO+GoQ0yweSBYZ6wjAfgxi1OZ20Uz/zeEzX5V0C2ERqA5G1+DYCDi7C
4Ks6EOkZCZMT69oC0wMAJ1e1vvV3sX/cfXtrxw37Rgd/q74vZEkgZQB+tWhYX7/uPq7Hkg+fau6P
ErzVPvlllO9woaNZ0aX3Ufl4dABlWbO5R0NLU1dLkg6Qp3egRVRu26cX5fAqU/BnSBF5+p8gORph
UlQN2ow4w3PDaoBhlnl1FyOg7gbq3ckX+EHj8WOp7AuJsCPrWJEO4EY2cZ+2LvqEfA5KDxvGOD1H
6Mz6ZZmn2seDEEPXyD40+mxcqBZMQii2i+wFRHaR9eqeFNXmnz3vjBOTFDK0zjAPb6qTOWmzW45C
1SqB7fIZ55IkJg7DK1nGHhVqexowGlWRL7sP20VtjCAFnW8ERKm37G+T4fJMs4Rkx8Hu+4Qthk1z
8+PTYOIastLvyNCwkECAjY584NsObX9InZfydAcohrPhkeU6/jpYCQXz3fvrJUHy3BSnDH3xtcwV
1/yZmgknVB5MHapiDVu7nD0R5XUFrRi5tyfHeavGp+RYM2YhQCkuMb06Huye1kMPdR6RqYwd7QUn
TsiMPBImQOlM1bFo1A/+CpcS7cEvP6oomaE5XClNkGdrXd1hCIk6PqPJBnHhmonQpKgq+3VOGoyH
i4C1C7nPJuKXKUxnK2ql4ZWcJNTfCTGFlOOdBJBLVbIYQBekPOmLiEo2LQbfYqvIx+lhwz0IxBCW
IGkq8XFyGI7eOxh1eWp4BMmfu4vy346Ja3fYqlKyKuKMCEahCYhgYAjkR0BhKMfDoglM7WXWQSy6
W8gkogKiW8NJfpqid0djx5eLfS5by6Q+SCW+7c5qEgwE8lLVH5LYa/3drwVG6nF/aQZwigOmBuZv
cjjuux7Bulv2YL0DqFNR6a2BGzNfLWPb7S8h3gdjO6c8/OeaC3rhfKYrWYxthC/VnFzBodS0dBWL
CWuOGEomdkEgTfAopo4yCoQ00RkhvddvlWlIqBBOozfAkYg8ymHNCcogevXjErwY7A++vnm5JueV
TSt5ko9z406hCmq9qUcbBL2skyYxQD1KXB+i/qeGYJt0ltlbScSehpH+eBHYk7zdmxd4r04+30Sz
FfG2aaHvOcqEpinTHGTKcDdHW1LS9JekODk2K78iZ8GQYG3v0dPV8GTt5nNdtxXgVkahNCHQ4FBF
aeKvs0siVNqnC0aLPTrqxAoil3n3Q+ceeClfJN9UFFUObl5BRYEGZe1fC50rKdbR1qo4igt99iNt
deoj1UK4TUU4LvEFRWfxG9yMx1yx3aWlSECpHilsxgM+AGnRlQM3A0mFTVY6pR9HCb5RcvG2JenI
fsZl55yU4rXhTzInwhu7nSPaqG+l96dTR/Tp9GQow6vFNENCvb0/yWIL4LLWNJWvLu0O4wE/591Z
5K9AcXCi71qWpcuk85TVccPcxbZykckTO0+B8Y95Hh8Ojba57QEEgbSFWZZZ9bxlA0vxA0Pr95R9
kgrA07NaPveVbDKJggLeI1LAShDJPEtUn0liEx3u2QSV+APCyh9f1aahUSGti/16yIa9xlyBtyyb
4Dvzx5R36I6mAjXY5xFrBYYyHo1l3va24mT1qLQtMjNqbsEPBP1IKwlBoFCSf4hxxHpTR8HaxEJh
5L1ouqwATK+jXoxN1hu4WtABRbjgU7Xf3yijWACWANnAD9LvWGYaSiizMU5LaTPMNeHwnFrbuEsL
rrzSyWTSqWrSPj3Wy1V6PyMJBhT5If1ZxZLGKNat+2xDICGbE/H3O89+nvBC+XgnGUAPgARhVDPR
TTHAmeyew55mc6Ws2wqcbj/RUjaIL7PZPLL7746kcW/LWwGQagKocCcM6Tg2lTeUN6xUuwEhzfwS
U9VFB7gulnZAQQL8H8emkREuiqLlN+RAR3kM7FouBlYla6GZjW1VfZzpWCOMLXb+jlQfSffz9a12
EbBbuFVq0pDFeRgn6VkyYa5MCwGrbzW+/Rs+wcXDlQCxKXn8+MhJT2G4IMlHkfRP9jritjbbmxB/
l7PhmkE8dWMPSG1iP21cY/Ts4NjZnRf4n9KbYkMq/2MMVduBU9Qmf5Uj4a8Zf6Gr078qBraSNfhO
/NhQOfTpuk6F1E5Pnl6rWi7Q0lK+USU79Uoq9Q6EaI4u6Lae/uNVGHpbp94in8bP30f/YdN2brRq
SaJ1VdZkwdzqgK0kn/4IbGw8SyfWOjJmA0noxJtQmQDHl2Btw0+tD5Jv1JuoWNPL42loK6lp/xb+
I0855HLlNQB+CSNRf2ACDEuLeNw6dEUZBenzafo61W/t6ZSneos5dnUrXJRbdw5wIQFFEMFpJIio
FqnWGQOVa8oRMbNoQ8ni7h4ISh+l+ZdNhSoLvMLJGtMKuAg7cZJ+yCf+A+v7xJAOHxY0pYP7flKW
H2QSsBrdG5oPs7k9EJVJKqKl4cJ/afAekET+Qbmr6Ec60glXycnXLaybDG7Apwb9L0HcPEZlx/uP
TE7GPciqFrQsQpkcCq3oz257EdqS5v/Wk223SxiRl6AsevFVBMQtTVNx0bKFB7oVYDsS7tdV6dAL
LvB/D/GTTjBvvUmEreB+lI4yDvtnG4owIUqNR1nWE10nRHsqhpcIfaT4rHy0rWtJSCLeHJab620l
dkGPT+0iALL6Tx+3yqWOAt5rmp3dnxfGZ36th7Fu4Jj968AHscIb9+i92hCIs8Myoes32EBE2dZK
HP1LgFJdUTXA0360vg54zM3OjvpRPLd7XutMtbMhBMxsQMvaFzXBU1OzGOH7ulaOx9v2Owe8TMsq
h495Ia5STYV42GCgVPMrgQ6DcUeVuuH00dGOEi7odCvrzUg6OWKbta6STU6wzCRJ8Tcfbr2QMEHf
d6FeZXFWojsfMrFnT2tdJ30Bwt+T5ixChQDpxyupr/7L3ubKTKJYp1yRNfWlmSOGUIO/UAvNjfMb
m1Ok0WhANa2P71hYMHgAfw6H0eGBZnTr4zz1uDGzksW08X6WkXpd4uuRGTZkT9nS3fLz/InPj2RE
NV5X38tMmT59Pz/awUcCxoLwNax7gsHYGZQvvvD0XvcfCno+ArEZYHfCCdZ4Sr8NH6rtJvlC/1RW
U6HjS66j6F7VQ153D4ucLql299qsGMV+K5x9i7/PVfZy+ZHbRbqPXsYQGIKfNDK4Q5D63gHeKBXM
JYElpUygGrEl+gqr5xFPfW/V7n68owRkswamLtTNwLBi2SBkRYdUENa3Vripbo2fQ2ZFkzKUJgkG
A+8OlEXmrHxBm2fPICxfiuybmKZYW4BFruPDA5qEjNCn0u0IzK0G4/bEKLN2dEbHBYc95LrfVw2a
OtcL/PuKxyhmGFLdHpun+FbK6Ar6ZgzEggIpv/NinoAYHo8knw8uOPltqVQ5PRlI7SfOJK7TKCRE
Kwy5fXwSwmDVb5jBqpUBlBDfcU6Jt32y/59JPL26qdSoo8qsLXKuoW7JtO5Pvve8ITX/lhKY8L9Q
YaB8ZnPQtkv9fT4i3TPSD8m1akbIeyDMi2v4+OUt5KxClMRPlqoyGAvIH8AVkE8AjI0YuzTdaiJD
BfzkS90CMQvRtuw5RmDAojXpUR21ellYMr6h7hXfm1Sm6v/SZQ3uS7ADxnqHhcuGJB7+2Tsc+pZU
K3cnzGE9K0y3dhTGvYZCW/T8esyiV7Ze/7PwGxJlJeBCPa/NZMau3DdtboXLRn63fBAOoXfsZ6x9
Ur6o67QXAjMMQTb5IAUofakSbHIb4Kz1hjwzpf7Wl/nSooZD7adEWIqFBpdAMGRKLXaairb9iTz2
p+SL2Rlxaaq3j5vukd5og97XRlw/BdvLZoYoI5TBKFPGaquDIaF6mJOPQHD9Z3NbqT3DtUcQuQc5
IIcNULWF4J3nLdl7UIe7NAHckqF+JDyi3kgrwoTpi+s2CDlGElyXwY9SDExGuqKiG3ger6XP+HgC
cErZBhJ2tuR4nbPe+lmC3TyKMJLJwLkHkzPNpYGA66l+IvuiJJqQvgYOe54DPxR2DAXZLdxfORkR
uWRkJatSQMQj7rGOu4N3YGHGBjOanRA95wArTP37mvFAF58xxyd4uMUV2r+StP5RRfapg2bTHiDc
4Pk4zLcSPaV4lhroljqrsto0AuaEreEqp5UbgRgS0lzOmxy/YfjNZv7T0gGquDt/Yt2JBs14oeox
KKkoNS6m6L8QwYDvjToGsSk26ZKe4ZC6YJalvPVHQgqUfRBs4+TYRQbYl/b5fJGaAZtemQ/wBmuY
qWBirdoBNPMLku3x8JAwIlNBAMf/LvQ0aWriPL6vtoXwVgG/ZOi4NY83jkdlRga9AK2nJ3YtuQgF
vWwmHXm9qt+7WB8Xlt/v4549MxG8/M7XPeU8TAOgZUo0D61MiOeTf4LnGq7fvXlL2w29pMHBkUJn
ZZckh/a/t+DL5XeTrX/ilHL3aAizQ91yUd1PDXnSXIe8zdo2Vejur7oXCpSl0TKnYvBHbFFprtjD
IsId1X5vk0uDurzY+MMcErZA6cLv2A0GNGf7Ls5zVzBf9bQwZJRgeeb3sPL9h/bHYXzawKLvyYZz
UE/uZrkCGI1jOVy+LAx5prXnj0wHMX9J6PslPPSs2dI73nOYDavUbf7qrNH5bN5OIWclg5dA4mHA
TAtzAo74tbShyfypuc9/QXD8zjPdPhe3hBY7LuP30emnTrS1ffNSwwXLRFomZwmzIDiKFs4eAGZ7
GmGmcNWJZl/Pyjcp6s61g4z+LVuYgH5c/nDlBcGEdgkdG/PzzruZTDb0MerolG8CRD6GXwGGd6fl
5uL2BYAAyuS+h203znAX/IHg+49arbXqcUxftDD3UBIBeJnazRx/BiN7pPlDQceMaW2pb9CsA0Pk
qPrwoQkSBNhsRVxUQWp7BCtBZyGJzIgt4OARfxAc8HaSj5E3dBzCGSJQi4ofOClWEL9waSNxwtbh
JA0N269JpdpIyzzWJqkHcfhVy+cEhx0iB5sBc+QOKxy/sWFpXKfQejSquwWHJIqxK4UB4Uz04TxN
RBF3ELcbrpp3ANXwn2IKdGMfLy25IGJsZy5iikD5Xqwu/xboez4U5EFB37Pd6TXtlHg7VBb/XjC9
otSdDWi4mUmsaKlHx3y8La7ZRRY3EOwKsrGS+AkErmPZ/rmwRO2/J0WXtkToKdRtlKxyRta2DIV+
jRi+ncJ01ZqIuv93Re2h7hg9uRIfB6+akoA2u/cybPwlVQ1C4nU1bdk4lVcyc3gn098kgSLEowT7
xU1HdMMsF5utGdpDK4dCXCuWCLI1+g7ZEUbTgzLTDVDq155QyjIZVhEfNNrkpudnSpyZ9m6K6xIQ
hu7IzRjVA4kl3JOFtreI/L6OxazlyoPodm5OR5e1+3Mf9bM37IlUJeCkqR+s5We2/ZpO2nOnE4YO
h/RakWvR+P8KBYduaG6tfyELwykgJdvj51JBZEzBVOaFtOG0ZeV3va3oXkTX6D91ZM/YNKnx17PJ
nMbB/IOjyEyW7Vt+qV7dxgT2nLxVNDUAwL/aqXOprA0yWahlvyQW+5HoEWB2IP3/ft9u4e87jUGH
2lDHIArT3EL7jrKw86U3ZT/2hUhHcj98vgA8sfYjkj2DjZzzdFefD5/Wz7N5Y9YPGTiybTzcgmv8
KfK0ZsEEsP4T08ypJVDTCFZ4vbltwBtot0ckn6cNRrGQ/hIGCbxj2Fq5+o17xa8u/2SYiLckb8/7
0YmyeKl3JEEUhUsesLvoailROtXFSsF5xqxrO6/cFC0LHxMqaPOc4U/ROYvhQ6q5N0VIKXT7prSd
BfofFRB8Z5kqyHGArZPjhyuBw4stdhB1TqJsocjSljxDXu1If/dYA2C41teYQxcTUKV7aaMWs3yt
wPifEJuGXnNtlSfD2ioVjt41Zdvfb/a23OjGFnRDnZZbsa1RKvMnM2rtbIhyiS0zOSJ8Mn/UELyC
h2YO9kx4f2DbkdJkWxEXNmDbQKqT3qZbWMvLNeTr4Wjsx+j+8QimeZN/5YnEY6DIkLAFqyEiT2OV
IUNpCdv9IWhOgfnmGJyqVEhcACY6P7ulMJLtWXjhwGmzDK93+Mj6pC1aB1Z0PQgeuOTZU5p7sc9O
o/eHnG3lSH+zqCq8gfG+1ZHgbC/dd9X+d5diZko6V3/s6e3ncZKudivaIOF5wLEGo0LEqlLzBnnl
0wBY1uEADAU1svCzFnFdkTEEO6yAJMLddPzbwy+K/YIESTi2MQcHuKW3tuu8RKxocIiePiy4jsE/
+FKBYCBBlZK36zIujHgiRJbf1jYLnlUXpwCVTj8DFC9U5JftrBPyF/WWCzy238dtd3JPBP51gIDf
fuxPJq+vPv63no/3e/72TeqF2RO62//7a6qA/S5ctMjE7Gd7T6paV6abmlBF9HCYdESbIHyO/RJH
d2KbdH97gjoOpVKGaoE1hYckB8P1B0QPsZ+CCJwzl6vK48YvqL5wrEdrv3FolAuQmUGCf/2xo6Nu
L0CUbpk+GHUj/EoTMVRZ/62CzP1igSsMVSDMVYyrQYD74AAlaIVWJb8kwF2w6R2bZ8PGiaRrdbPr
g2z3GF0zuRQSz9J6mbuA/aa9bOGep5v8WGYGEwzX7+Ag32hkWSZzUrXLGywNspUBueztgY+LLxJO
BhIdoPYvfzuGRD8kJNkzm4fD/mbjZynzvWloIKMumHTPIuKH79jSvvW7jPwo1uqxRnlp36vHOWzu
HJJlGP4V6X+rRflMuC6VmP8SrFCwqJMX1Bb2wg2dIBfdc2ZPLk21aXfqSoRubKjjGw4fGeGiuYgP
XU0dRUQ3C+i5UXdazyXEpbNIEJcUkp6LfH7gig+MPRwdq8WY8mD4IavvIdKCmhnQy8UUoFYDrcTI
iqDKDfrM8dmqcDUGC8U3pT2N7uI1orKkwwc2X+0uMVYtXnADNYpt+0cS+zvZFQdhQ0CUE6cOTMnC
jSq6QwNQcRcqZmLmRFXQFZ67zEPrxSwx348vVz9ACmLGfzKrLakzoIhnzfti2Ir/Lh5OAwUiNlQI
PULbP3t+AsojZqk7U0VbH7V5y/Jdc8Z/2QS3v4GhhR6j7wlAlZs5UoMT8k538Lus9b9TFh8JKNnJ
UxIUYPVEGpHtag7NY8PSjQe0cr7VLpZizXTyys6qHNt3d6a0bp110mzgqEDMl6jTfO2KEEFxH8cD
SFTQrvJDHtMx+nMFCURjjHTDjfE4MI1UaIGnovtboYexQP0jHFaKX3mmMNoIKLF9XHWFA3ydl4KG
cJAdV58uTyGKNtypDHfSyOMcPMOm03JeGS5j0l43cOlWuL6buiTJVS3h5zB3ltc8yWGrN1nV0fZr
koYXVxO8eW/GmLu2q3EL2Pa5mNAB/VPC9DQKkk0oICBnnvX2fdZT0eIa3X4zv4Llaeb+nGnfJQk3
oV3i4xhpa4gm9SdfifO9tK3gokIXZQSnNBfA7gbW0jNMebk1+CJWe1Yx8Z/nIYROvaK9TBaD0DPq
4xgy0lXaRXhZCv0Ig7wEEt7aAfHRkJhZbmywqD0CRBW/rRc16zWsJZh1vI5J8YCxe4wCz787zHZ8
J08kvnB/rFL4WloV9HF3L6olfmHFZbbAypav8j7FqcNnIxWDJRGypugVtc4wN69fVmp4nvbtJna1
li6ENfnukzjDFOCxkdhw2Xg/P/ve2TIlP6OUsb9vV244DfR/qIKswzgGmZ7vn8IcEZfclKOOKi+x
jbs+phqEoNjlaeCKIVGv4GGtR8C8SuJtuaOrWbivNEFib1f2ovpAaU8OX3X21+3+6oaOPEwj4wTk
lJXcWIE46yjbRr3otdqizgYKbGsE5lzyfrIUGnG4lQoB15rpyu1tM4kNc49ySZSZm6QvUNIEyXi3
yOJWyc2OgsVD2nbP1ocTlLybYWEDX6NWA9cLzdI7ByZFXEAM/ea38wzNhR1dsg7osL+twC8QYDzz
4Sb9rBV9jLBW+2BMXhvoKlWGJX+JCa3UgjrU4B+ekqBdI9AEaZxf8SJw14ZL+FJ7AYtLhW6rpXub
t6DO4GHJR1qm6QH7bIq6rI8Ry7N9A1x/6/O6X5LE34qrrYCkvH7TcY7b+QyaNrO+dcjrxzr+aNUR
HEJqatV1Xifu3MU5DBXZZ3/IlwFYgN5LxO6+bSiZ0tmw+lntvnWylf0EKoLAiQvyMFe4iuYCPppc
672HQxy9L/y62i9YOyoSg7+XAYOt7/DNDfINYWHfq8gvzBEuMOo53rTWgSAu8zYLzfCggxvQkOf4
zssTx0QHoGW6Zdm1nz8TYTvNMLx97ebDLg2Dalz2iIcWzYhVbfxpU61x/O4Do8gShVkeHko43VaH
0e+aiPBBaHb09i+/f5RcCaKVC/C3hinXkf2RNFY0vVLARJURQOqJMRKpJIZr97Sf8uFj0Z9c1lnO
3k5qUQEEsyT4ef+sLtvm9mK3BIC/GDTWAPlAxmE5bwJ74Luy+KopHY0NXfeJweexyoZqrGphMh8G
MDasF8O57/w24fiXjiT9z44JpEIntto3RtMWBOkcacW5saGWN/sYi1H3NV+MGdcmYSLaJhx2Gv73
MScmwQ+fAqMINNo0bGq22KFR4NtdvSUzgz8KHRbyKtouz9mKEjrNieTeAC0wtwx3lvJHCixgem+2
4+ZqBYtoPztVOOpZaHkymeB18OXfl3NlGgm1ZUuqS/IbYK6Jp+bQr2WYcpzZ/y85q8x2D1rPKXnQ
6Mv60WaYLMeY+d29PDamEiSqDwIV/6Q0mBac550Dik+8c3gkp90vkY0yDb7PDqe4eA6m6+HZ7vXw
rLswii7iSg6V5Y+lrwGcrxAngKdQxuZohr+cU6JFcFAChpRN5jFarFN2EhGdDBcWEtXOeZEmONCX
PSKIKIO+6ChuOjzsZ3pVVJi7qgT/vVEU5ZfHJsSAVg+SPaLa7Ff/rMuuEoj4p4F5hOFFbH0oCtQ3
d7hof3aSuAvrtiXxWgun15hxpgOlmILrSuPAeyn4MDYn4v7CrDHEO3EFjGwZ/6V9b3Q0GZtHKDYB
H4Peo3sehVYSjFN13/gFV4ScLRY1Am2PLyVC3P+rd63ttdw6mIDlLbUupVZVffTwMmJMUYegH6cW
p1cp0SbbpmrN7/Zj2ausnjZomDBFYW0t9+7kXKJB813u8XMZyClj5CJ8mhpKGIraaMABZMH973n+
8jap60NP+IbVpvhzcz5frO+ImV1skMTxU/XEoXIwpqfQqTtfjh+/4odZftUuvr1IWtYtWf1ZLmTu
DLQZjGLMiLiUG8jSCqjD7x5CcYMdzWPl/+nFlBDoDrrlNvp6ZTw7P/j6JYuWcnQicg4pwkQ9ENHQ
yLFu4L8ZO/kFlDUY2zApG0pJZ1tPP1rUIlu5KIr/EUSmUY3M78pB258WiOXGzcyL5j4xpifvFaD8
e8TggE0/eB9NmWp8hrUcllUBcNrW8iVMA1/i8VSiUPYXiUkshqRMNjzGG/syDrmEvKMnLz5YP0bI
bwqq0dqWtGEzd1+NohKQCyfyI8DOWi0NZNYPRsmlu5AfiYi07o65qQcS7b0NnIsPSArSUNNs+I6t
soJ0Obr3uFMmYm0hCCYn9EaBzJ95qxWfccLsLZeBdulppRd5X01wK1JwTk5qqL1C27SIVZT6MYpu
XJpSRF3BMiMFlDH66PCqiLowyYVoJ87KxJPVk4MqwON3njWjYcUboEhETamPfs5FwRAgX+c89ixy
St5WujCpcFJx60aaB+sWiAlJmbZJ/Efnj/oQw2YI91Meo9emW894dbLI7FEKSMSxgbk/JdhN11S6
qh1TjQZukfEiqF2ljHiQkXmKNxdBFYJbUdSGaqQVCO3/slTyJnSOzl2HZ1jmFi4H6fBHIYIhQOoD
YHPXIs/CkLZUuKX6zqT1ry9fkf/yZcGHUPbHFOZvvsUPRvpdWRNUCMzmpns3s31/nct7VOewMQWK
e2oxVQMVGxrhxMgmlcwzbPyJqw99I3T1L5laz/zgMdR4TGrgQagFUBTkywLOCCiLYhGE1c30pKr5
c38FHMcJiCjhy3a1LfAiPvH/5t1AMAvpCK5XdTVRHKc6SkebDUXxX7Lk0NlkxYY2JxPMykzFjCLK
D/oFdqjgMjahX6vJCK/sHMooDKhy4XXwnk5NzDLD69vtYkN5/DaZYKlZrtryLXGN94FwS+wBlXgA
qN0cXTlWPCxgKJ52eTLBfQ0bw2+bWYFQSNQ6rPsR8TdKOWr/52QtZmQ8KnVH7CAzVs8t13DC87ZL
Itp8MH4K4Vx3PoACtGzyVD/Kjv4UpTP7E8w79yFxwrM7/rcHk3pVnjuMnDLjRYMVLGfDo7MeCxtl
i/nQ5GAiQdt6KIso7GOGmRR+9zhlfxQIgC+YqcegHkfxHz7qait8WWDCF7xILi6QowAmWWA1Q0oZ
MSbWgoItlhSUkyeIP+ZFMF8PQ9gzVl4+6fb5iJFFZT4mDbAx0oiBJy5SL7kf8/uPBRCxC5tD8+Jo
I9NhVGJWP1OYfrymoUSOo2lAvlbMdyatUS1/JFWrO+hv7p9tXuKpVArfC0pB3x/VJiv3Nh6SVnh7
9mqG9mddrvGgF9EXlTnpEIJQMkjH2rXooOhJB8LrfBCLUwiNU3Sns5KXB50Qoy3hrayvuG2Tu/fY
w+5xKpdHT6I+AQ64E9xIdnn+hUfnWpvc8DYMZMHMLJXRf/0KpRVelL3+yuUFRumxamymNDcZjDov
qQdEgGzC8v11FTjt1jKi/2Cn2og24uiXT2Wdz5RSsuom5sils6ufZH+2xzH7lg9sBQ3VrV9ACxny
pJZAHp4l3ofu/XrUiZjd/wi3ZfINFMFT2bfbD4KulceSwv6GGN4Hi0A5iQhJl4Wa0sr6O56/iLxL
8HeHaNgxn+WNrKR+xQvHqtCnfZJ/XiIHQ/fwbELb4mitug9G7vy+wdwnIp0FOXpJ2xxRGJYWcgyK
7DbiWbt4UuqSMbLqrgSdg7lh9vGvlz3/G3Wwa0M+rlfRLfuHytc5XSueeaiwb8idFr6jXRaQuOue
uOy4VJql77lF4gr4kf3bvw9cEhvGqplX2P21t2vODmlRpiZblM11b3lHrwwOwVtV+jY+fZ8Rb96z
YD/xqsrEbmMLpv3ghYZjUlRnqdCpbEPhs0qpLSTGfmszr3zvZNbOgNuEnvQT0t/ELeLPGGLDHEIv
+Kd56u0iw5kcNCX3sRjMp7hQ195Y+dIfgtRlO8sBYM+F37Bn8xO287V6Y5Nw2DDRc0nB9GTYi/uL
v3/UGnAV6Wa32lGpDf3hNjZss5Arr1KqyhzThibJTlJs++f3nPxf9Qt7Ut0Nq2z5U0+mb9Tp6I7A
MMQppExq0hVQKEG5ztDeXQ/l94D5+82EohuTZQDTi/9dG+/qXAwPeRm4QsU/7iBxfFsH5hx4ar8U
SPop+AZZZ8h7AjPtGOUjVs7fg4C3XVvr+NX/rcm7tTRhDUnfNsIP8Fm9uNyWtz2VT7tFBmigaCxV
UF/tV7HDyKfGRmqFQSRpqSX2kOBuOyb4Icww9MqEuR7qKMuY6JhyQmvgL5+My3NlzNPC/Uc7v4C9
C1Kcv89i9wzWZfng1UhrVRjPFMXuVSquMxXDqqlD+OHDKUzOxDni8cmoco4kK2fPoZdzxpVW7WVH
B3fTMLBjh9GXlJUqxIJgOFjiuYG5HqNvf85kgCbia4GDoeGMfmKsgFmTVX7bgmmKx48QVZPyRDzI
qnJ9YDTOpYpnNSHqNYmRONhynfzIro9pVIbXLWdVVIc2CoAAqqzyk8VnU/UTuJSj6BnXg1iuFX/O
F37NExA2njAYpsH6XEzbEz+gmPm2fj984AGqhmFahuRuaHysv8lhEVYSp1YISBTtc4L1AQP8n6hq
EtT9as/4dGoM++uKofFazShyts27Y2pqE7xeMSqWFKhT1sJFYZ6qpLmyun71pkqAa4Xw+mCt25LK
RgT2ZSJubwRtUSqsK77SL6lCcfbJHk1PgY155eSVnhAR2oHM9D+3Uol9sRAxYoWxGQmooELVkXVf
9ygq0b8qBR+A/xuIAev7tO5AiRh3dmMdn3IVOV+yLVFOkMYX7cN6RwUhyzOBrCFJH/g48mrbYRQB
Qe9sPvd0HnGhgnvLGQnygU68hzCJ+cZbNj9vzeJLns0MJfAKhNzW1d8u3ICbDIXtWUuV/52gMCBF
EOKDbwolPaahdcv4WyZfzxDyyY3R42F7INyHxZNyKjn/BXGwHxtk2P9QggJXVu7BIyeAyN2cmUG/
uOgY5WgJOOVkiOKU11tcZrK6u5VSc60j5WPPKO0dneDuC7JxheUhNMc7i3/ezwFmQbxFZaPy/3Rk
dPngt7xHhQ0HFnk8GYt0c2afCmXT4TI1VqkEE1TVtl35nfpHy7eswtKAxK39NPHnvNUlC0u4CN1h
xNAZAiTFgp3b65ulHSGbgD4hbgXZ2KLl43tcld6oiVYu79UPiWTkcNytLz1A/VoYD3SsZbCJ7UL5
HED+xdvHWa7JnEyu5IbIW2VcfyPzn2aO2s801avmymisIySAm87co4Pf6Tj1YYTMh5VDoH1ogO0u
yRmmu9zZ2Wv1ycp/dfIeM3YCUh2MyQeTszcKByYizcVrhgemm2YJ4zDn28T4tbrTDUPqkro0yf4H
wHlVOUPRKMTSfIJg85iaLWWjHCI6qSGyzOw+tMq+KlVyl0edfAv1Ukt4KcHcfVqB4Zc+K1TWZ3qU
yxYG9hhRkWXBct9QoVgN0esfJJT0imWABGLmaUyuFCseRIMeA29tPS4E5i4RKhiWugknJKvJizk2
YWrhVtICM7fl6haIE15ydJomaqHoiKnXa+JvXATdaqQMs03yulLxu8YxWFkoJTyz58bd9WMHJw2g
IL48IuGRopccfcahUeggNyRE2OiL95ssJ1jm81o+yQhRwJAv97N+qOFZQgqXV8wRtkzc68rl5ihn
GwoGG8Dg7LcKuqLMITf1CuGL+tEtjFd60xtTVrfwSIWnEWBnUBfDeaztLoxcJ34sGW+AaXNLi3AN
x3VUiWkz3hqNu9N5MJ83mb497Fl8RwOoCam9+KX+FqwfG3j0spzl4osassrqcNHBQHaTqni0K/M3
dmeNIwMSrEz1qVnHc9pTr/pw6J2H2wxMzH5cNlIoLIgXT+QxyvNdzJpyGwXYVdi/4XcYKXMnsZv4
Du4AeRLPZvHsydfv8WxOyxvkdcDVtF1T+u18L/rOkWZQmGGw71C9g8kdIYPQBHjbZeV98OU/BwN6
iBqNbM2bPpFX5yqZGm3KkPACTvIDKf7gyIEri4GW1YNXlmY6CXqUI8ms5MngccKdDlMgE3mCyoHe
PICKdLNil8N3rWUkeQAc/nzVl2nz1eQSQtQQ3v9oRz7yL12m4vSg2Q8mwgqPAFMZLv5Yz6DNVvxz
HEtdNmTjpI6sjipsy/SJmxVcRvfAxeHUXKckOYoUGntz1QbZfkPsHwxKsUZGzsrQNmbPt4iMkU5G
Vf8ZsbCWlU5srnWhZxFgmydpZnE2U2LbsPxGMORcznNdLZl0knhgC+2q+YPq8iUc7xzwlZYV8V+L
gOc0UVPcuNkcqR2IlHbinplbwHAXfLXt3NDQxLUnHReCNfnlT80GNLcXXYKp3Hyc12QKm18z84TK
nHpYZV/bHPek8ozSQf3fwDEW5JxhJrmyT718hPe0v6swe10V0505IPeT5vEW6sWadmrPYr1ysNvW
vukTi/cQeJzQETJGAO9LSxiCLjJpnVajt1RLGmyex4A3SlqXKzFGPoIfa45UcHCNSp8cnM606P63
wxFSWvqqevlBUV0x6o00TcvucPq9rbhuGmlKtovXt9CnWYXnKSBmYQMecdkRwiUwaykixVKmu8Xs
DVMlxQ1CZXCjkd9CM9jQXESkXDpkzA0+0AuN/PnzQOB+d/bOMwMiBQIwTGzHdAaBix36Gla362yy
iap1Ceb198+T5/49f21nmzzPvnFB8o4R/d2+wTvihVMMK2MnV0VCXa8myaPEZoPcRECCEHb54Ro+
mF8nDqwGF3oFDnNmoTFnbGVn2dKmPdkm7cNfqmFI7rwDyIL4VPg2loxDjiPBdK/mqHdZlQ/l4NUu
P/4mH77h4MBUEgfpqrFg6S8tJdaMoy3biyO/djtTdyeKJ/pffKb7NpZVSFDaW1aAoyhYuQOCjho4
apWru2iMfM3Qp20GB1atCu5DClYICDa2mFFtwb6fBFYq2wan0WPPMUk1XZU163+X/nYZq/0tw8Er
ENgtoMEGHO4QWFa9KBx7DnCEHqwax2ySGPxVfQaHtMkve1naq8WVmW1zp7NvSnt6KnvtsbMov1tS
UAgtkQTU+dSJH9o/XzrLNtyZj/+AeqJt2TGek5fRFtgArDVjEBO1Z9oPYAFt/EHbWhhO48ATddII
9+02RUiBso2n6VUotoITFaraAG1y5/J3+/a+32JYa1geFumudNaFBjbtTt5Xl5pNpcbSEP8Shm/x
29EwDteyzz4LKq3JVzGrCyCpViQxHMF/xH4alm2odxptQd+7PGvsBIdn5KQBW+PFCO2JvVmevncg
NGCsCCtALC7y7KHkVvF3WRxs0W5Zhs+8K1qSozcEGG2w2fZDFpN46DBwsDzDrb1reIqpqgM0qw5j
6hej0c0zGU9Ie3Z8YSEgQSaX8PY+gazas2K2Ge5PIXoMQ4JlNiu61+paLmyxJuea36far/P2QlOn
QxGZWtJWdDGkrc4uwqgkw8XH76YXYmKdrWrg6Hk2nq5KEe9ZZxlu6j/HiEuH6Qy+/A2wzOW60d7i
AxgWibRG6N/hPpSiyCV+zfy66nAwmj9oFZ7+B3zYCYtyanwHKFt9oGfO6xktvJwBcLZ90LeiPneW
MYKCYcNPGAXMsHuE0iyNSX02rYbwnpQ01xQJtVoXN2UG8g0xdH7w2rv5NnpW6z2ObRhaB5WF/fo6
FqqTF1ZdhOfkUh35l0CX5Tacj2crhSG5LJ6EyXZF8pM1xYtRhESS8h1a760YhL0mId+1HGucBsLf
pblQcM6k3pks5Rg3ZuOu1c7wXb3RI3MvrKtfJq6VvxuqkUSIKb+aPWZnAfKvp3r/OTrNJLS583Uv
LzG6fdxAi3m4DzSW2YCQPeJvaxMpE/C1HuMwV4mpA9M66WXeRNR4lqi37uxTymdX/T1Zze0674ET
2cAP5TEMLFwB+ncvsLWwUJ5wN8RQOjjEnGY2bN8bGN19GbxONe2AkY4FzpN+K/GLHs6gtHEKLaQC
a0oLkGAVHKAHQRnJ7aY5B88bTEGDLs1Owf1fWqSi/jiMdf7reA8LoyZSUbvEcZZsjECEJ4JAzbAD
RA4QPsNyaE7DcsYjbbsscKAcojetC1Wysbjxhx5BfEhY+VYImugrmAj7Z9gSJiwIVDEJLKGbHLHW
dY0G/sdkRtmG+m2IuIkhePl7DPKL0dlHFUZM/oiL/+8Xj8aptx0h8t/TA4MUme398RncTr4Men9X
aAMckm2+GNFE8gPLsUogXjod0mW93G3+MMVyK2rrxVMJnY58ozDD5VsG78ptKMsDjpJfkiu1WLVZ
9RKEJTF+mWmctiOAGYSd5y7wN0K/dp1+VVKiJsy+V0Rfkz40I+vjCvk5dsyahWnelkK+gc+31pK+
tsB4ivQ5UVo2bHKssC+cH3AP6ZxuW+w6FRwnKErlmC42wmBNFzeR/1YugJplSrZweSCeVN9MM8N4
7B35K7RBFqgjTdVUuXt1+UfLMQEqFj0+b/51KqfEBncDocizVHWydAdGQiBZSAS8k81lV33CKQ8b
Wq89EHzr5w0mwZHpvrBg/EQSPQZOT+ksFTVhdWQlO7yn6q/3Nf6Jg4uZSmTSpvTalpLY+Cwz//Kg
TyNX1hOXmHipPy7xrFbTVzr7iWpsxToumBZqMyIwZVX10Dq8H5+timEEt/abisYbvm1Nl1THpsVw
Mh55ZnW46IMw5Dt/Tf6gC+11DskWodg8wAEdmyhe9xK1qvxgUX+OJrS9dtnpef7m5POrP/69tYCF
q6J3r3/dhh5oxrsVD6umG6nMC+OJq5VNkpXkPqtR229WZVP0IGBAJfCV3tBa2rsEnBxe2L5ncPkp
tCYkhNI1t1hw8Y+CKyocRrJv2aT6SBA88XAk0eZMBNgd0hRelHwn5LHq4elBTJRRyv6wX/S+h/ez
XC3i+/lJ9YO9gPDwZRIbrN7sWtRSUGzzzMhRZm1oXsb/qcvKgkNxtoS8Ma9ndAJUcSlD/ie1qHyN
wDOqw8HuuRIInly32+mjwBBBrnjGR60saZna/ueru4p/2lsw5pvrNunUzsESe78shw9wc+V73PHL
sihny87NlURXBtmavvR8O0IYceBe7BjQu42Zmwx5Cyot79plO8rFPDbyOZ4ycc0lKP28zDOWVhIR
E/jYdYy3TtH3gly7mesGVYgYio5O3r6gt3hbk+vNxdtZkMrufpHyEyX8/+4pcq5eJ2TVdPnz4PnO
I4mXBIUjqFeiWT+Q8HvEqhBGH5tMQiBAytRWPWlPeEppJmiyABgZW1Xm+MNnHhF5sBUHFe6B8c4s
2xjCrH8/V0crkfoYD6jmihx+xglYppibmAuErViPX5ULyaTnWYuZJFORWHmywa5VEO1OmSpWdjEI
mRPLNmJcSyUuDCXLQwtTcLXOFsG899M053uLYgdUN2YMKNGpzZCE342FJ1hwky+lE0RissDNK6ES
3qBwiMJMc1WUoYqabTIBX6bvRLc2BHMGgd7st9TsZoOic7R2Jf/SDxKyQBMmYnoXbGCA6fqV4uLA
2Qx25gPL6YrptxNqTgPQFjcSMvi++oq3iURmF8u9F/lh3RvpMbBZo79alfZGvXDELnHERZ95N1f5
AAwXVD3HkJ/I/PdD/JIk4wdbPD2sU1RBbGLSxu9O+JjBKNymA9JIXJ+PsrCCwdNZZLXlehgu8qsV
he1eD+PzaC1cbrdbM5ikF9wocjTWrDWwYlQLK4UlUHG1MCneJPsGIos0b/OReJ8PdJrOn2PV9k6u
Udkdxuo8OPd17evWF9H5RIdWccI8SSN9W4dSBnLloTRcxdNcdp+b6jpe787NDhbl4k96Q+wlUg+G
XaJ9S6VwACMQq28h0x61zHpwwxukg9zjTm/qVh5UiHQfI9btUiw9MbHUwZZw5Ro0j/5cPS+nQVjy
uhqgy/dHgpG+FXpa65qXVrXoj7PoKDj2kIdO54DW/iYKkAbrOZhnvic2ILI92XA5U27UNmIzhU8V
V++uag30ak7Hpz2b5GuYLrrYvd3kSL27SvfSsAvOYJR1PUV+HUuSAMxZ8iE6VTILrrbqxbtH/pAt
CFP3S/iOufTpxN14wXQaodMRc+mZ6MDor2Xk7LzgB4A7/bqs3Rqf2p57GMdtd+NJLhQQGIHIfIwM
9TWa9ISeXXB8BuHgMcb1iqKXCI3Pzh7lac7a1Bgyb2VyHC2TycDcai9lZC9DcgJjzUAyzoIfIeZf
ciMNbdhMmxIZxx8nG5IclABouqi/7DLeD/7UoPo1iycQ8rJgwek7Zg2xOyL1voCQBzOi+qknur81
MTcWm8LElS1T6j9/XphYR1Vy0mOPz+RE515dii0GPMTGEpedaAo6FVkk0JGsB5+mYSvJfi/X4UaH
pabhzNLLDOAjaUeTi6iFOrTNt6lEdDEJs72zo1lCk/K6svnZI2dr6fk1qS6+BzkxdsbbBbh6d4sz
QQU8I4mmPmQzpRZa6u/l8MOKEgmj+ZMhp4DE+yV813R0fDNg9Z8NOCCqLDD086rmNyqp7tFZJGoF
3RI4b4sIn1P0sCpPo9c3ZhcJtL3S1AWjSKeVW5ZfolaDS1fLekYT/zPYNozzb18Ble7OndA+7QcU
rA8uqMaVWZYPwXM98a0Tjk6b9m0EdiS1quLq5sNPn5oe1rvV+QxDk5UXjxAv+3aYxHLH8fYFWxT6
8hkUwb9ujN0giBjVDg3zEhAPI7snHIKO22KPogjHgdmtHjvKT2QliezBkxujwMTDnXwCWOvla4Zh
armiC/F16gIlX82H6O1MUvtE3GEqND02jcw/u4M2+cmy13EB6tXNonUJt1w9uOFH2YXq26lMCxkk
pta+4+nkLKEFkK7PRkBnWliTKlT5Dnow2VIU0g7XDNxeBLtH63PWOORV+TeohGPd7kdN7rw5Gx0F
d7gvNFOQVSvTo2rrWh6Xybau03gsUg44hez3TfaXsObUR3G9quToP/lEgfpdq8Q3b3U3x1AgAKAn
YE0JMSd6tPVmNRjvEEAFNMq0jeUSy8lM7b6dSoCnhLrbDqtbnSZtyFVSlA+5Bgq3qsY/UX2BQNMe
f/BAOQZ+PFQ9A+iNEFk69kL/bCKFPpCp8sacfN/SyScqXPJP5MhC+i3vT8hxhcUwkJUJIK4UVqaP
h+TaWsz93/M+4LjYJcVYPgLJm4U4At4OTJdwgNXko3NOAnnJ/qh9+Mxc2jtb+QMqMse68k4Jp60t
KhVkjHrBv0lUqWyLk0de8FdVA2J3O4Ev5j3zddFcWY+LhPnyr3Lwpsa5txk/WIPhRY0J1Ys934gV
Tn8hvM3BionR/zUBnTKWAguKiPH4AyTkuN/WFUcolv7pfrei5PbcqotOBlnocPSt2tpKYRyB+kBh
35fw1BC1wYsZh60cE7dDz5/UK4t01qtb0V3LGA7r7ZDny/Vu0jczRCOiOGbUvSYiotwTl1KO3pMu
WnfX8cti7XH5O/JgAWos9beuf1Tg3TDNG4dVktLhcJUNUl2ZSEQg/edIhu+6oojVM+1JigGQ4Y4O
VwbP2MPLZU+p/9ikJyLnWOUrz0A3pW9lZGWw733Cqzd94k8zt/YHWA/4/r9Lko6wsmEw9mpUj75O
eO9izLTIWpuu3/MdRpayEurx8s3ocCHxjKzGpAHOUaAhvmKPGPIl75Vz2o8e+3Gsi4PQvtoFmn4q
Id3xYa/lez2CRbbjRXR4PrXy2lIRKkXXQWre3eSjyo+sz99WqcQO0Q6+0sULa2fidnhGNPdPpUyr
Y+aMokw0/vB+zNISHzaJT/eKZKizoj2XXvQI7lGz65nL63layGr1ar0CTCBhdDbFQ+uEBqEpUWyl
LWr1IjlRRLl7C2KzrUFqx7CMyymmlJfHXOi+n3HRsvAHU+bYd1YPC8f/7Gt3HHHavcRj/rOYLWas
3M+NU3uAt3Sxk8LlWBkU+VStoKI/CJVhsQejCggvwr5aGJ+K3UPOWgjwLz9/lhwI2w6ACG1/4phU
StZbaKA1+HSrkFNnV7e6F0hJnONHrfVLy45QQLFdyVMC1nlTLaX1jtE2eiCpLFsfyb5M0a8tcN5u
U2GSiixzGiUl2fiyUp0IJT5PZQ49OpmA83r0ROLUzbIuKy6VEgYCUbpmC5NLbHGGcfKKmTaLULwW
u5Ujs28rcO+a1HEAmoCk4zgWYM/n6+BAq5aOHtFPRzX30fj6M+T54ZJBjRua37bSlWTUyru1NetV
wCKQ9dRyhLkzQf3XDcThIXdoFtwYUoDhr/p6uFvq0kx624L08H6XCXSLxoWoRfceATRSLCXwfNJ4
9UHcP+TSA9jB3MbSsVhvUT6pZ6v5eDHu2T1EnhWKX+A6phOjITLNCcO8JXJVW8DSr4MczuLqB1js
pvfA0ozCMnoWaVkrQ2pNMDzEOmtLHbBOsoUAwYzPBvY322rOqjPwGM5E1sqMjJq0sYNFfytDcuVV
J8Jz/l6r5tNnfrOpilAuT6EpAZIpu2pUaOLMHNB8VaAzv4oXBm9c/lUItqSVQlD130Z10kDPDtD1
NvcSxuV4dCzVu8asPvrtqEQ+/lhc208ybwgRlQFBVfQz80tysUQlpk70afsej+V2Z2q1LQJs9Dge
EgjoUvvWmLk22Ey0OpAdP21FZ9pyg2GxXzEukJby+UR9MKqsAXv3IeRKLHW0RJi96e4g+//6d5Fm
FEM7g8fdB5CIR54aVb407Fbmmd0y/qnbSR7ntJiUuxBtca8ZIOCcf0+uvWkWOG9TfJmNyYVfXDuy
U5y9kScb1q/9lccP6rp625MQa71ov+8wRZOe23YxjLv3FgaQhLjnPGh3DfZ7W0Tn6z7aJxr6kKwd
sRSQBNF/Xl8y+uu5kVyNmtu/wZFjTiXX3HGkPz4tJJp9ZewcYlK+OCB1AHsYIQxRBXQSmKlj/Sih
tvdi09sfNWT/icUDPVnm7RLfzyEhI5AUNF9/W8lHeXrMxRLIg+TOrbYG+BlbMilxEpHsrQpe1bQD
aZT1YvCLfL3wWGkwySzo1z61aUXjo+jvuuzgDWs9F2VX5zRTmgaTHl61mWlaf9aPd6QohaNVoKSi
48GRtsOez55E4jZbxoem//LdgJxqKPqPbHNJuXJIvFYL3D0jVJAxxEbjvAePfHcfeY9lGM0V5QlE
qadJloUeEFoV9QTMAeDTix7/goDuM8uHuT5k2taMVqBG1lJimCadHW8jkh/F5p+F5W4sp96KamWx
3ontcF6CG/pgXHSvnrgPQxu9ClZxlkCMpCW7RwgRvKMXD1odybuflx1mvoel/8PmB38zyg0A0pvr
VeKTU1Yusocy5fA2lREgK22dBCd3WViCez70FcgYRTXdOLHFx/e0cVx14gRiCbpqZWNiBkBf7BZD
t+pEMCjblsfNoeOTRi+iZz8UpW0eoijlhcILpR0Pm6pT96N7UwF24moHEKBJ60oa2TAMJV2ilg3m
kbDpqonKlp1Y3pLYeUiSdbbrk+jLMRQXc5F6bPBC4YrA4uzY44n0aQbNxidsay9TlfjEUleGxd+Z
xSnshHBFQoetEO1vx0O42f4b/v89k3qjotHSbhexAUTlGJ09bNwQHOIJ5Bp0+aJj7AosLOw3OU9e
oh4iNnoUSjBdIlA8dAGiq8J80dFGc3NABl5e+XLgnTelxraONPUjdys0NzU7Z/eyrsI38yuyM9tk
LtUzE8M5a8o2FPH1n8mNpDOR9BLikrCk5UlwQ0WkYf/rmjkHJbARYk0yY4/9UmxtKGwML+zfGf6w
nSe9OgLxMoVFH8lo1K/T9xmf6Jp1lQjDRblfIF1eu758tMAvTAbqsqZq4QFykDao/kubHJNpDuh/
slgcjYdnVzLsy1OfauEYf0k8dk0uNKAc+F3mPLuqVGH/R6eW/RH9V+/fsBzAZT6mb3VWUIiIPZ/3
oXjKmVo4T1J+egZbD4Aq/Uiml7/fj8tpNIvHJ2rAXzDpLdWH7UdEuFlwLgDsPghiHlfLLDlpvPo9
jgOxOG+JmI8VQ2ZLarGz172OaYhdO2jv6MWFTAWDPffTZ4m+td4LlzIUM+cIwvIOAuBQu8FIL4nH
llinV7jfedNva4X7kc+ZSv01r4lHZF/6qVxxYUdaIBiPKkfTdMXA4hfsyzczyQ5+NZv/SU7h/sww
3oQLmAmTjypk+TduUq0dWAGkb9DoZQjiGIbDrnX48Fdwbs3gdj+QXnJgdyMJgrdtlxuCkha7KJot
HGUWcJMzW46N9PzokyEDjMOdmiH1ICkDLqWaBWTqBdiNtN4mHCcFqM8CBV/z/OhjWlo33eIo1Sdv
n5sc6sfYYjKVLq2H8OAW/RK8GF/H7XTMK9D6XkLt/xXX8LVkvuVMn9kykvXZJqLECSLl1ddlVF9I
QrLPCmTaHIzk1rpCJExs4e65OnR+xXHbmI0HRxhuu2zksBYkJb+jyRwfCoUJH/N0l2n8pxQRXuPI
qgnmdoCRs21TrHEqVaFJ53c6cauJBfuoCysRDFHtW3hPkCb5kwGjw/OGKJgmFii/d90K086ZLSrP
8WORYnwUXhAEf8iYAqO73QbjjHyptUP7dvVtdRQ8bFLR6FKoBwQC3cOR3+ESXKTsGEaU/VuSmqEL
YYfUqxgBepmQatooZQ7Ffn2+EAhtSzlo6Hh80oZOPOrm8s4orx25rp05yP6nHoU2/9ZjHGDcEELp
PJwo2J19KB67MRondmjgOhQ1D7gUu6ojge4wZ/2xmxqIEfvKuoUg8Z2wUnqDPWoEpLk+xLX17b7/
7+gekfLQcW1WxTR0V7n8nC/Cu8AyAbf7VErgk+ndupAg8DZ+NMeICtty1ZLI51vImY4gFUX4R0oN
ZBrA/0/zRJztDSRm9P20DgBvKsz49yYpR+uFVm/QmQ7kzR//MlzOzH3tqboTbDL383vClKl1nobT
vXe+gJkkf6du+a+ZPDhRzBl/wLHOu1tCjdk/oYARkWUg8Wv+HkK2Qs51+1bQPxKwOU3iMhyidDHI
6R0HyVyTSEtBPDc04s2+3O6rwBXQFdYy+6CmKJXpAoy5jNG7fnkobR1O6aCNbitqX182wggjTZSE
HAqTb+nf920K1Cdf3+kqp3G1qrSpGnV7Ao2mwnW2yzu9rYUBYSrST8g9tKCYPeBUMD6n7WZx6y5H
tUJRnnrUEDtv66xoLIvxrNqHrMsq9dCLbD5vTKuVUkg8W6j5FPlsWHcvm+h33lLhx5Tnpfowh6Fn
c+LnJ0PHzFHftEHDBZy5/tMe1BVj9wbEftS3JEx5GkSKS+F9mEZnxn+SMlXscO89oiZS5Xj2yETp
TsrPcIikubN4XHyo1FjuPHk1cPcQSEGLX1d6jvqGYMZM5sJDMYbq2+3aBJQRh1GDGlRaicVjgfZY
8jVEdzJfZuGKnjikeBD1L+cs/Zyrkc266BwlLNZjX3P+17gOnG9KEq7NvNMtsHA3XHzJm48kFEFj
01jl8PLZSXpZ3e2vCnpjB5+V1WYAiTNsMkGvBs9QT5OMb+SHrmfH72JFwbOMwQ3dijhbjsWykhe8
1mmDTd0xMgwsk124Fhu+/QjP9Z50v5VJZf0Vh/MNjUUSQZ8Ft98OsMm9eRaSwXYU6Rvw926rjdLI
1vdAyphaAI2q4Utj6xro5+ebg3codl/T5wH5eY/AcJPh9yQ5TtK0OxvBd0kWtQk5VS9/UMWqBC82
GfcC8J3Cd0TXcPCL/NVifo2a9zIU5WVAENaGtcF5PbbTGqraO+P92+6raZIIyd8QS3aPb5TwM2HU
WRTE/oXwLEOJsWBel50zolV3UJZW2DJV1wnew/XJv5AMp7ulAQGhbyP6XMKfv029zV1GD8xRVHOg
mDqEAax/0/h0jrlRVhFohDi3oeVqzTSm889lvoMDvpF94OG27U6aepUIkU56sqV8s99x9w1yUP5c
ttN1DX/JiPPjNisHf8SC1Jip8Y0lbWeMODC3Vw6wdb8i94uCoVBejgX6lfbPf+h3HMzqymENTFgQ
ROCL3rlB/gCrb11LR4BxW3A8ID+GVDy5RcRcHKyunPJ8tZkI4hu3SVnbia7k6m37UgMiXxNHnfaw
oRzjGLe/JPrayUqyVAMx1UERmmsSHf+i/7auPoQAZx67MbKXHQizmNG2dD+B1K/5WpQ5AIXq8nPd
J/f0G1+FSSH9JSf3M1wL/gkomFzWRYied58SNsFRseL4uWhf7O2t/Rr31nLiRF1SIcrxb/nOsDpl
HdHQCJmBEBEYhJJbYqXX+q1ZzmNwjpETzOhlmWEDnMY7zC4fe8XZinMTZa14KDT5zoamgY4GOQMj
zevGh0XLE3zDWUWovvzfgpm/Z/ccpzWZd74qf8pYrUsTTPrhhyy1wmFtvbMCV7imoK7tRZtnAkF7
wtfn6eWV/mobnfcAeEA0CqGvbVhhy5NmR1Pml6XsJ57RH8F3f7luKnyQpW8OwZsreNmD/8FJcfRM
aRIXbJVfHIqfdTL0Tv3lrY30TYapuHIGWOG6Zt/oFHlrGMDjNolZn9jzXurevYFirKqVH88Bc4I0
KKU+ElHQv/KbyGb7ctrWHyEfhWjTNaUkC54myiKoDd3enF0lva0aYcfIFBlKZ6Xw5qEDgaYMz7l4
j7zLbrmgbvA9WXSVyIHZVVJWaEWJ11p8n6CSmYwQ5K5eDXHJMnQJ5nLULO3z+SQL2ySgTTuFOPE9
pfFLzHUgQyPqfCUWe2SV0uPEFx+xArxyMHqUy0AgaKxCDt75CpEL2kGth8hF3tai+jQ4YpAAziQw
DKmlq39AAd6yVL7alLhqRo0j2u9x+mfYyxvgUqJ52s3SsqQJUxPq23KPxRN44CF1YvyPLqAKR86t
Cu/tWsBfoQVvFK9WQAp8p72fp+FLIVv7mP1Eu+1n/luMM8i4oruQhxjaHJ4gMwOlx3Jo+xVla19S
j7CPXTzPygJqFLeiYftiNcwAejrn9ck6py+PmOBk/kvRJ73TDvq4ihN3v9PNZ42q+65hMeoB3opP
gzDj9KkMjmiw156u7fghoLMtmWsHe/ip2gg5w9o+b1ZVU4EC3VTsUj7E/leXj8jVd3I3kd9sd+iy
HkvD0VffaEh7jfK8zAdSE/Ayuzi56o4SPidJLfYBwDlPavxWLrzeBT4Uai9NekPybh0wmw/cFGuI
zHcO2hr1XsvpSJWIGgrSZEZQ9DthtlXwKcRO6ija7Oh8jIsE6fo6eWWbQdrlxrIvsxC5i0J6MS3t
/H6tPkZdXUIGUHNL33Igasjk8rMxm5PTXdsEixlNAB+xM8ervNRvDpyJcVkfMP+eoVX9BBE4bSx4
sNnnI4riETH/LXeH7rzwE2p6CXetjOcPMcKQVwbO7KeZtvlsw3+IvbLojD25A2hvOUZ1nJgv3rqW
yjSs+/EGY1r9prAKTTOxcX0ytFiyZB4Ozr+I9FmhlFpzUGExmOsUXVI5EXuu4L7dxETXSUzgp3BH
ahBOmKNRMieSgQjHuHP13PDguqFDWRfWF/Po64OAuxDujCvpzLl2c68zX3M8Nv7tLKsi2QrXV9qV
HQGG1D/Ovf1HqdsJ7cjqK1JKCs/nDYtCZ2kPiZBv0lijyNQ4F13Dq7b7+PzvA+oD+nETCpFsdLK3
02OXDlj//Uke2wcWRgyaj/JKI2M7S4+VOwWjnBV1kU97wjHbPiWES5d7yRse/cTXmL5ZkiJBV0IR
gP3O5ekveqtKX3qESIm8JEErM8yERRbS0LJiI+g+Xuwj0h7EHGxCTA/iO/AzGjthQR17YtCRaDx8
7RIMWFzRXtNHWEeBcm5XgfhKHp81a0IXri8TSYmczZpDjL3ykkOiDvRSwkB4V18g6UKpoib3/JJb
fYfZXL+228yxOmC/rXRrIRLlnJDuwYzwcQD7z8ZPYiCkwpXFMKcwM/MH3X2lXhcOrdeFLDI1HL/R
1KGNDPxWQf2JM9dUUT9fEOEpQiovAbrp7cCHmNzlQ97k9ZjCz9ovvitVW2cZcl4me8wBdEXz9WCL
nRy/3Qb76GW69LZPf8diEyjW9zwCcKdp7lOWURfrRTxk6JA+k5TChxZXahm/XqrxuFGgyTrwSjw8
Q0dvkW6w0D4Oa/z91zWVbK2hWy6zTkoKmCA1naXY9R1euKqiuiFhpdwdg//BY9SUpTBaNLlUeRpL
W9hDjOlSMe8TVBEK8W49D1M63Dv5k3R5Pfr4dpBGNJ6rr5ZytPYC5Md/juBiW4jctLXo7PoHsIFi
eqxHLMOhO64HgOUFu4Bk6/ZMAVSIssZnmyCcfrYJOQga+xQxSdLD+ft4T4vZO3S3jyVNnJKr4o9a
PZg4BuDurNljXUsBEtPuvMcjD+wxm0BuS6W8jY1YXMsmVv/EyE6MxyQ9TBUoooy2D7LGZeLI13eU
HcBa552eI8dVWXqQpBsqGTPc6dcnkmutVn29Od3Gl80jWapOVeK3YQ/igvXsyUfoAiMe2Bx+Y3qU
o0OYqX5EYVGTdHhtq70cA7EcXA1BxLcvSMF1lcfNMXE/whKM2dB45R61i6qOWDJ9AoKmJOjdi+RT
gVrtxLXnQMo57QT5/rLeoU04gs8zquCkRz6tiqYCAp27d0CpLpZzJnQGfh2cPAlzqgq0sebLW75o
rxQ6t8wX6xtWQI6fZmFHYxg4eTI8KSVnRgb0sqAV23YYamlBXdTTdJt/mj/bwt9EE9qaz4rTy3xh
hnkeeqogEdyxpQ1Kwogm0Q4GbstpPybePfEEPuat8TWWX8ZieuOGAf3HGUFcKh4H9zejmd8KuDq3
5UJFnwegiiT73G7Mv4Gj+w45oBU5ZBV3Er+XvxcOaGq7DGs7cIhdSITPUmElzDblyLxkE1KD8FkT
pSEoB0VDqYsqcxcbPzLcNAx43yqveKEIOuyOkfTAA0D8J7iMdVtZAU2A0/tRXBfQ7XKSR0OsyRau
ZQ5AE/0IPHVa0OqHID23CdgHlDa9uBlQT+A5E3R/qzjjlvvIpcHE6i4YaUCwskjq8ve8W4STIYOo
uIWmugaw//AQArEH4KP0ffozZCx02m7n0tL2+cNMUm2LNnWYTlLamm978DGDq3zDQqHhe5HG1B/9
VG7tqzQQXpS+dTPbU2EgpswLIKTRrPGmh4W1+Y2nnK4rgPvTxKS534BO+xrlLHUWiCw4Gvgd1N9u
gHrVt1Zc2F75JqZNdQ2XZvdRX9VB6qzbb34rNimKXHb1v0NvuIR3vX5/TnL5FfDmtB8Dz9NNH3x7
p2bzxYhRwqyfj32nquQUESXVpiWi3JXVJUJ1rLHWrqc8aD9ZCft/h7MZ/5arl6itKu98rJ8V3yu/
uCefSgHAUpNg80RYfB7Tqg8U7q1Ze6TbFkX+JMDuY64ZzSeEpkivj3TVS0jReZcwkIKSfRdo1Uqk
glMR77QB+R/JDZqhDWRi+WHU/wBpjnYQ0OphGzPTjMfcn/1UAnpfgjmA6g7ypPaI01gETZycEm5Y
Q0Hh30Z7fwvKJp08eSxfeERxEl3f3NyWug+A6HJWfCUq6XNbgrtdl7CiCJugMSvzh6ZB7pPgEjO8
YvOPxP2Mz2k1v/jmItAC/EZrNXtr/STR9uOEa1pxMUy8X35iqHhT1uC7KYy9vt6b1XwDHB44yb8I
s1yD/uKqi8ECWD1SWFgkCuUovKui6uPVyh3AkiyFQ+nvaLVHn+UlHPMwLBIi6i0xrt6XtLkG36A3
tHnSBSLzFh2fiTA+dKpPb2DrFekLl6WiLXJe+uGkytgJ4sfZaJhdFeJxqmO3mP/DIJR7icnMeWBp
BwuK4aWCrv9K2viOVlgfsOdkDWuGuen4QfE+Nxvbg8koHYDQHjmfWrCTJ50N816QaCFV9w8Gjx/r
kpy4s/jaBJKd/2z7hwZyENqPjxn4hlS1IGEKc5t3ot57WHygmt0b1Emh9kZtEg/8VIN9gKDSvXAB
/Xr44gr/CK6x7A7txMvVDXXGbmwFm+oVkmjTYz3d5qay8Fn720qBt14A2Vp2QYeHtEK86wffcNNk
6cp8bKN8PBCNC1H5C+f4DWAnJamIkJDGP5AXJKusY1TJ5JzfqZBp4h4U9Mt2Fzo+D+VS/fp29wXe
Mvjaz/wBW6cQ8obPDYjcjOMkDdKHNYrh16xSNSJ15mgdJT5QlF103HltSsgLr2XNISIhfG8O2WU+
W0qjBiYFwUVt1ScWCbnD5tzKOgR6C/+ebqS62Ok828uHbGJf4IarxGF30wVhTa3HBl7llTfhxgPB
PHfHOu0GbSWkS5M8PAd2Drpvhm2iiFxi+8T/CMxn2+7KuZ+PiZU3XiL/GdpmpCr+/ecbvFBxv0gr
eI7k7/C3qjEJHCSC/7fcv1jJQ2UIRy7m5F5UcWxdyZosUnw9w9mnM2EfsJ9lD4AccdiRBRIfawKl
jtY1wxCRv+ZfJ/awXBwnEldRylvBj96W0Evos+KwtTbBTpEMvbis3E/2adqvUSu+u3zU+7wKJRaj
9UpHeHOSk/gXq+HxvQ41lUZ1yo1NG0dL48v03btHBdYRS6jl308zTjCHGMBXqJ7LqEyCX5+dtOHB
K/gc9MJ0g4bbwh66Wie8LRPFrytixuxbXYk7PSbUG/LF5XFAWn2Rk6yaTTkIgWekBj8CjtI737Ge
1lLap5XHzeGMghMCgslnm5yiKHodBWTH9qA1iy4nm4Xm9au1pGW7+eYwt76CcBdWa5Y+d8LH98c4
rVNOoXSFYCgH8StpUZMh3ZX3bw/Y7dZj1JRwj2N9K7eh1eo58db/7lmyzrcotOmMYdFgfWQf6I+j
2ZUO0Dju3UMdFs0dRWWjImW5rvuL/MS9r5bl0q7vhod+Y+x0qNfBYYGFdAKMlghphOQHxNYQv/do
qZJim2Nn6dW/MQu5jv3pOvuvWgL8+aMiunBpShqGQwnB6PuCr9g+hw6lMRhtd4OfnpnHPcQF6SSJ
BXiiZXkj/wPsgTdbwexNY4VmOAbcBA22RH7Z/zTdxTAJzWYDZkOhQholW7T9tZbjW/dFvmlmTxzU
XYLM1Vx9vNr/xtLMf4Cnwrxw7syoK4NYZJmHqh5+TVdU9MvP+LPkt9KqagdaXwWy1BPZsmXwMtX5
lou/rGgzubd9OMfuzeTq+JJgWLKBKnI2LOfMxDfHC8GQvqCXaWAcZPZWJghdG4jBeGsPbeQJu3Pp
2O/ZooKy4Iy71vTld237mng9M5aTWyhSNFoWhMcP5MkrqG+Sph/XINVi7wlTZ/J/8D89YvNWcz1V
Q5zIyyUx02yVZeE3biSEP0piZfL+n2qzZOfccTrGJl+pLNRgM6YQedUTi9kpDX+SPajrSQOtc/iE
BF49mgeUOr9OGellhS8Wz7uvDiKGl9pS6a10ALUzW4v0SlOi5fIyj0fG3ytj93PHofv684kRDjXO
lw20oxVVslc0UjvKLSp2GLC84Y2TLPjx9SpzU92mEZd4xDJuqeqwphCEa1Mmwpx+WGkh9KsFTbsk
eRenr071bx/7wNR/iwKEijPUrssAZKny1aSkjN3uuF89bskFXL0Lm4C78UNJzVzP0Fg1Edvoo3V7
WshPsvn6fVdciiTjhsfnDeFrWBL9O3e0yvDVcQvoJEcC2O9rCschq0XTBy1ITJVuKBij46Haa5Cq
1q6nLczZl0ZJk2k1hd1GYQc8QtZruwZTr4o7DkmWORY1ixjuSk+Jg7rz58gdc4JM7IlhmGuGsEF6
bu/J/CQqcAmd6xAwF2J6MaDU0Q6atlbQalt99Q6X3hVO0LsgobPEpkB1xq53cTlDxHImFrsw3uSB
QwlZpdHPlugFrtR5puPDzZKYfSgO+K/pmZKWSp6GtnDnwLXtTKdkcBjQPC5aaZEygs3sZ6rqqg7e
F9wOu0/+T6lHg5hryM47ur7UPWeTC8sSUnDK8Fpsc+bAdQZqY3+Is/sC1kw831SVUJFyvIT7r1+e
f51d1b2DtaMWbA1LJWNXO3XxrDayucq4OAGL0t1YO9+/CAp53lvtKMFTBa361ni/ChpGcYYyAJIP
WQlQBGRu4UsImP3YJi8WqzZaGEC0Kl185Y5m8fuNAyxnFdvxicf5Ihah8OV7+r1sJJvt/TxQbBxQ
TEyzolY1J6wNLzhyE5fwlg58cpmtZTvfSMtD1LU/HOfG7Dlw4Uwf0KwAy2h0wSwXM5iEPekx9nOg
GxU0bRkRqzlKWwdThx1BUNOrn17Xr7BOKQwJ7569f2K85rsPzbS9VBxnnkwssAlUETyxtGhGXfwk
ZLbWbjfWDeRg7qDHc+cqeqa1bmeCtYrzFKTGycscrwhFNAFZaFEQdKkEeC+r5UJTQ9yZ05orZIBU
6j2mXbv5aZFKaaBfFbZR3ANXT1nDUVTTZxRsRUx0dkYZQ7Dfh5WVKw6ENxR7LOtcZiZvMFl3iXbT
E2Y5f5XTh3NMEyBUUJVWl/Qqa/sdeJrtzb2odtRE81Kcd1cKD0+DjFJIe4RO6OaPi268NUsxCC1f
nSQYoyPTFxoc4THgMRbVm1j0iul8o9tq3PHW0HzuP4hGnXA4HWy/GSn7ezelwyJYWDFZP48Hb+7F
PSXyvvAoWiVQe4oBsTKXtbvj6cb0cQ4SxCqe3LioieA1wEouvuFO038wcepwRCjZPOkxSvxUfDkv
O48DSQcMJyC88Mw8YtooxAVpE+ixLi9lHeyl6WrbOm95B2LfXstQtmoVVcLEqWx1dWDsA1RCvjKj
BwcIieaXhEDab1NYViN98wRwdLVALhpqcleAeKZ3MxSm+DXPA9Ktj8/arhln/UKMR7DEuROIYn/y
ayIddXGXeOeRo+Zn5YJVOrdYBxe0ouJBZW246kKMuKQaaBw7hA4qDj6PIotuindx7KwZ+pFTP29s
FTdavlxJE3llX9F0nFOPoERyOkRi7R9lgQgMQIZavyYEsJOG/MgYos5MVHKbBBT1JkzcVllcTBqh
I54c24+sfweCQvP/RNyCiKTTusQYJj9MXpDiv9T8G1gpW3oqcOy/eCFDUPccIvuDuiTIt/G/N/E1
NNI6Xuuh0wOIzoXhZKi40C0MKOnKFVi+0HyKQdL4AfnSZNd8JvPyEXjT5hGbkomp5s7KkNjfKK9A
nA8hAsh2DRECPQQ2F19pApy15LtZeOwONYdnZGmX3UL8e6/2lHF1rjLyPYZtiK8o0iE/trQHL4It
XNfXF0yo/4IEYYIjOzF4ldc/jKF9INlzbgnu4NQ9Rnelee8DkoczYZKPiLZfYuuDCYNqA4V201yE
KAqlARv29iIQJzpGV5SGHvKCt6fmcmUbWpxV4d3eMEOEe4Gms3mpMmovC8Vcl2jTeYDUncpc1lA6
pUwp1SlE/AChd6tCcWcnc4OTMDZXNt64zMx/xDy1sFqKJKhDbP9uATHNs+ZMbn1V6x7H6q/bIu+A
AvibN4vuBIJQX3ljYEa9nXTGBOV+jHE8RNkel+6Y00VmpC+PZNixtbHIJHFCeGsuGi4KNZ0UTKOm
3ZuNXav/4vrBK1IioujgvssnI2cDCew5AVUH9h09FkbPzKCBuj7pY7Y4e95coZMOeyN8BuDpcEFL
h+9Rtmft5X82d/TXTNWjhhnN9xvLPy0jJqA9vJlS/xpdJk9dxc//U+4QeFgdFwK3b44VKTfwbREY
MW8THJ7wvEc5hv6JPIe/IRFtid078lowzmN64Ziv5SCUbB8UdheajfeXpIvWioLcFtwDqA2ek/sm
0uwVZfP7oE80az2BoEMau+NGidHLUV78rjeCTURWe50GRrcydcUm5RvzUqD0+WNwF8xS4DxhTq+z
hKil01c3vbqHY7okFhH6AV0dS2PptWD3YswALUod+6bOgqvuDpvzzwOQc9lhU7MYyVgJndMzoCyZ
1vPpEWoxb5DpTOeSsp8h7oaXIbKBK4HnA/a/CkiWVLE0KTCC847ahclMpmf4096iJTusDT28t9lt
uwkxQM6V02+VbNmiSIjjy7MQQM/4kRqDx9Aej+x5jips1XmtQ25qncdQfztRMQUGCyA18zpQ2T4u
H00VuiOHfFdp/4u281WpU3+DK0OuOLWDC6BqvT0+FfiukMLxp2h0EJiVPzIe5DAop7QttFtaKvv1
pJRLHcFsHBX1/yzNFAWMv5BxeT6P8emOqJ8mI5zEMqBKv/RNzwTbjkm8GIMnMNlnpUnQEyqIMMEc
3ZF4mIq7dm/GgF8Dv0zjr47D5PF8Gvatlx0vzOJuGfVQc7WPYm2J96kxTSP0mS0fc5SPNguI9BoN
FrIdm6iF7d7rJOy2QZiKF8Ddk6zGMg75ln3rWB13ti4qTLxmNPZBnp6hdb9laxYj1VLfhY3mrPFu
HY3O/w/8pCU3h/uXaIj5w+uaIvYVTxpE6cBWkqy3TS2kkeSQGqJKtdP2HBFTSZcHcqlFuVrtfMtT
GDUko43nFsYP42+QrwX3F3O8If2F4f4/C1Kq7fQBeZbjkxDEzbt5HaV6ngrHLIB/z/Hi7jz4g7G0
YJqt1X2fkuMptJvTihk3zGBAUrgBZrDdgb+GF0TO7HHWehkeF2DOqtwxK6ryBTLoPCZu0w3ok9Hn
rEHhSF86tNmO0KX1xQE/uVnk6PIFq+8qIpTKXKit4QAbo5cIIAsoQy0RSlHPE3/zaxK11tYuA1ib
TXAiUOiQOz4XVFzHRIdWyoxgXjDMrikiiHZ+2sBkZOWD8/wAOt1yeSLfTY3RcKA6zGeOtqxU6mQu
w2p7wtcwi207s3gi8HKw5ZSM3kmzE80YqhyQmte35HeNn6S6S1U9CKvf4Rm1DpHLNoSkbA+w5dKi
aH8yn/n+n5rq4So5WUhhdzcaz92yK28X8sEFcN6/mjX/nM61Jtu5ewM/bJBBMKHkbX1tZnCnTcJK
G4je8a2/CmzTZSSGoTteQ+JzvfBpFSzMZ8G5dxtXE/UTvejYuN1fOPICSIjOxaxFK8XWwnlZ3Z0e
P+aQzxEP5cB4DVkioXCZycjBIuF5D5nPC7MDp/sQBXiSZjtPN+tllzNIHBe4zhyQdIcZ1O1PMUqA
u9jfqnV4six9CNwAUryiVCQsYdmFOXVEBTmOKJpQRYLwOUJ7eqJSKsXxo+L2h1798lArqTNEBwi9
+JV2/tOIGZCKctlJ1CWswqXb9O5os+IAsA+KDk7wRuRHdAqy+QfwiYDvMd8pE2syCZQEa7szpgwz
rRvieAM4wyv3YCFBxZvVpCiUZXfkyv+BdXlvkQ0dNpVeJPFJPSksIk34LKNtgu/G29eaaOUtF9fa
/PKI3INfR+X1RQnJC+wgvgdaTC6kEAMFueM4X/i2iDkFonobP32wx9xekH8eDyvHvXSZx7Voyigj
DFAlIIXb4PqGMn43t9KAZa6/PFdELA7iGod7U2DBCbtwa0UdF8cp+QUT7eCKTj4c1J8l+/3S3AAs
yPLam/tG/RpthFDsFNE+VwlCOOvkBeRafzHJUewgUy6HVxRy6jt4OvCX2WgzigrJiR55yrx6diqH
JmPZBobnM7f28eER+cD3gcB5Xjk9IUlR0bFiCoxmZAwXM9gANrokxPaT5z6a6PxVrIlHGydjRA/B
FbfdZ+kOnQeN41F6DaxyJbyB7anQMJ3Fped+ar6TMaYy0ZyVGbeknbsMCWInG1YQPs2zRfJAFRKm
nPMs0VvKExSGqGq3jECapaYjUnPyBfmeskIcJ43h/RRqGRZRyFVKrqMFXHAu9l1/e28suewEOxqp
TeJJmJi2VYFlN3a0qqjC4w8w1hAYZsqc9X55aAD8cS7ZdUuQtHgNTkfp+8UF6F7ifHce1DSMzsjn
MKFvwGEUnjH5xzY/MwAqoDtEOmAffzgshy8HmRQVI5G0zvhckx0QSMiegi5cgyEBntPSOiPjQD/x
bV0HY7HUFZku9KfsGziONd73ZTdUqBHPlYM+s3FyWg12w/ZckpcKn1pM0I6/rwrNa2rT6bWlGvrT
0GTZ7J5hnLQqPp9+Au+4ZXnLwiENVD8bcRhKOGvd2rwPdghwUIWYWEk4be/zzzSmaO3nq+LPmOOI
I41seMkB/pQ09InNob3zF4SsH75+3PSXZ93kVZHZjyXDgdOMeOMxpy9mCsYRmd7AHs2JKR88ap5l
ZD5fBSrk1Mh495hsV2U7AWpj0hNMuo7FaqAh3PJ679e0y7HmBZ0zujAbm2WMcsd/sDNo9wBq2nru
Fnp7KKQewON4MdltvnjbpMynF/1CYCDkJlD78f+JLcKsAg9um+1qXcY4rRPeRwgztyi7ea028x6L
6t453iGNcdXDQo00PtKlt6x1VeZPUwMh3w8si8h0mWmWQo/ABVbeyj6cnL5pPLjDHj6yW2zUhGII
u0ABsuTTXFIE8SriZC/GcWWAgHeXV01EmoNExvHzbqK37e6UDnPCkcWhsmYfIj1hsruFC1ZqEmXM
1OnzX/Q6V0Ms4Uf3LqEAKT9cbrnqE6nCAHXiWNUsL9W0lenkrO9BfuTD7fgReu0WMFLgm7sN1mDU
7PqjMjDjYOQJSgNQjla8mA5xhLv5AFb35Cme8qycLCtKvTtGNo/3MwkErj4ZKvj1cRDCE7Q+dCYy
JULC9K/FKRb4yHpGeOMp3eYYYU+/w6v6PHDi4lQ68LDmGIPkoTfbc3P/oSi0MctfldPAWh7Ax7yX
F7800MDkIEdofPpWLzAZFUzMUVLPmnm2TFDOkec/UmljlDLVTuCovv27pZlFv5IaAcgYFutH4jTq
Xfm/m1Bxlk2Wni9eCcWiATmiaoAUMu6rhj6VoNukQK1pdCLVk+jARNvHwJtCgHvT2iNqXdPXYDuT
MSuY29qRgTOcGd354WRqS1dDNStV/26ThVW4jbu59KVtL6DaflImmlcrAWnXHvKOygxQDPPR1+zD
GfVdV84p0e2qd5YfrmjnnE9U0wsu03EF/YAsoPu9eRqe0mIcCX8++kuMIFKzBDVUpFAgumtlzQm9
5JqV3tiM4i/w5XRPZhR9hbHEnt4WiNAiVAFHaAtQv2N8V83k9cua2D+KFsxPe3yGFZEIyV6vKE+4
8WadYMFsQBsNkPUYbVLWD7Ua2nO3kGb8jYlZb8Jbn0k/NFeyPlMA6NBFHK0g79ni3UB5gJj0sNA/
0x9SUQO1eioUldLy8tW+UX04dT/MpOGi0Mlb/ZB+vBPN3RGM4Z7EgoGs4uuyeeTGsavNvWAzaUJ7
k6gJvwrRqYSiSQrYN4x7Te/LFExM1AlTtHvGn5UKBsUAL72vY8M/gDGvBBJjg3cZr4mmDgezG3No
WDzg4Ur7IjoVAH69wb7C0UXzbleakZ1BQXdI6eybjTQObbQptV8HcuqVZgmM3uvYVYmHnpWhZklj
9QeD/fRejcpWYjujyc/Qb7Fc8sDbF9yX2bzHlXqdqRkzRBGZbj+QaNg8ZkohJ1PD5ypbtzZsKE7E
9bLUqL1qDOleHGXLHktV9Z2rfmFZmOsBv7v6r8e5Aj9bvA45VtfPiKvSZCsNvmZ06R+ZaCdlgKlW
0FY1qbQGFhq7+XkjT9a9NDwSiDasoeocqiyh/mMh1bkurW/6gjD6K2111JBGcoj/HZKojjQ3IiNo
FJ+ddawn+LXZfXL0JvMudXkZMCB0HlOFJftn6OhvZBebKLgysTcEuEMROwEXCfs9lx6OgWewjLmg
83h6K7Iy3Hohj1b1C0S3iyAGjKAfpsRpF6mSLNcOshcMrbYPXT3YhfE/teRMBXROE/RE2IkKgVAa
HeQOGdSc0DXKMIcIxqAv+Dp1lgU0wAAvg9vPie4vVLDqtPyjffRyhdZVgPX2i+Mz4mPaDJrPiXVg
FIN8EuOelTyKJ10G2u+9lEIeMm9siHKuHVvTonMWmVFFnLWitR1/cTsdC1cCPKVhyNL2XI7K4XYv
29AGfBnDIw2CQOf4nLhOABUvt3oZ0O/VS5O63lUxXNHExDej5KXr8u5Iol+6JdrBJNoGN+EXsai+
/u1GKkxeV5TT8TjCrTGegB9oE8TLq8aU9YaEAWBtuwzzGXTbsPwQg6aMEf9IVdvXU3Cmdur5tk5O
K9PKHUrpZTGhhiApJVCk8hQGsfxC0DFRdYb7r9xBPn0Y7iRAmFVVeinyBJ7xgZl46Y3/vuMRAvD0
rou9MN9WOCaOcAShhOcZMp0fpkj6aiNsoyN9GZ4Qe3iZEPCy7ZzUcKd/lUP97bLBE4vmUkkHS4jr
nJLE3R3/iHbG8go8VnSNRuA2fiB9kC05UUvo5Hsvbk6SqpEbnz57+Dd0IWynnKS06A6nzAMi3jcF
K8V7A2Cz2vWQm6j4bHi3KZaFqzyeODiSMKAXYEPLAESKXNvVtNEOP0tfgWIIMpREdvxuve+x/DuO
2xeoLUdlj8cN4EL2sbHZX/Kig9T/pzvvgkvzqFzV66cLKimZy565vxGq+UH+hb4XDs9YBFVpjQW7
NAAScyj7JYxoeoiiHAOjR3d7k8Iq96meeFJnkP98Mr33gT0i41YzBkqnO4OBt+WhP6K2Uzr1Pp9p
C6OWPMaL0Z1cx1qFs8QCVUx5esT0U30As170rH8elmk7YWld8KA0Qek2AzWcifmRH+3c/L2lglUm
DDxDTXKcBbLNLshRCszZ7Pjd6zoU6OAI0FsV+FQtGrbFUhCYZO/pfII0G+WHnrmI4lcaMtuf3zZT
RT3eLVrtHvdw86cXBw0LzqoJZVzEwC75PeOzXECvRb1bi/99xukGdaJ78MryaAw1AaqlXIpPpppb
7H96AGwhhBFcyVte48C+fLmlIJxeALEZPsvdPzgc0QWURUckxUYISePcdVyDdsmpYZ714OdvYMYo
j2OBPvpn6+07bezJk6xaZ00zcO3msLHUPjqeQdjbiXlvcJWVA+/MkYKMloEWQfCSNnjYj/+Bnbnx
WqEPUKONIe1KH9KQNHdbdO1c5yNr/9yBW4z5m8OUO4rOqytrPsfeT16oblOO5dd1NKGEYQAcJ7zP
7HsOOqTRCejIAY/idZQ0YcynfGASHQsoWeyTd0gUbKktMmUSKif3b7Uqfcg/bajLtIRpZcVPEeeZ
2cHAiItOG+7dqZcZ+Ji5/iYBWDK3zED+sGYEYrxVV8OBHcRF+HWpPbV9xUn9wmdQ5Zjq13MOGZjo
y3NZAZH0yNgU0R9CZSStat+DmCS/Cd41/tJNjGam1DvidSG7+Dah7tfMH9vfqon41Y2MNMwYxLY1
x7c1yTzxZDLfZ65kerAJOrYfHMxcMRc63toPp4DBRnUUSegOUt09Ff0/bGHk8MVtPxBHQ6vxs0HW
3UYbQ024rzrqYxvLJWkLmti/v2TYUjnbnjEiLqIvgXLcuBQY58PpEqo1rG9L4LEX387QuLO/FjpQ
bYLjKd7qhlfOZFjgCVi0VoUK7jJ7D4qLXK8hrNJyfLEKpZaUR52hNFTFi5Nz8LcLCeEtm07AQWQB
q6LGN0x45XSppx2JLuv78Oqqh6kOIqpfrJRPcF5YJnLJrO+mugGkqqkUOkJcU0RgqKz2tOQGs5UK
1JdaZALYDKGkHtqLBPY9JFqtsE8eMrMsGS/o13T3oNQZ9S3Gm7Bi4ib8L563+3O5gefZ6S1+uMqw
cFIsnucWxkwAKgumoZa6RuVyq/0jucLaG0X/oC5ZcK0YwkkIwjwnObBMGLybNeqmBlMJDqUHyMia
oht+xmlnIUMC/SFQg6dC39pmR/N64gb1l/KmVAh0B0JOnibwy1C9xchgIdRyiuPPtJMb9ZOMUeVG
JZE0C9x29P1PwSsb7xlqMm6eekaoUvgf/W9HS76s/8CK5hs8afJGmInJfLwIh2YVIetWZAlJ8Xjm
BAoVQJxv+WH/xnLo3PM8MvgJYUCarZiGutpRaItiQKVT/l59wsH5lB+m9V6jH1Tl8ljQjdrQSSqb
Zd5sUxHE4HGIAxNV9KWN8CsDopjDVPMzYXvx596jV5Md0cwD44T3gIKrraKqu+gkJ2Gw5GyTyNWP
Ae2JPRo6hie/0PkaaCRdb5kPYXxiozp3PA7ZmRW6+NTgpCNkhZKLLU1sgYy0f8FuChCwrE1S9/xG
jR4EJM57Q1zK8N/SG80FCM2B+MJkcLbux1mA8cyERFaHB56xPB8pLoAY3Ya+jFIJqebsgp6UK4+W
WQAVtHHTk8F1fMvJcd6uOs19JQLw9qHxWt1ZzmiffJSZPoRBLF10V9PX/+jcgjaKU41+lpgHXeT+
qNbPYVMLv8xveDpFWRvZCDH2uJUG0aKgMhAFea0nBYAWDew7TRz4ntbW/fBNkhQTMsgasYAPwq2V
CLIk+hUM7XP441+fYZtX/0fvYcp0SJMGxg1TgBlTqbSLIsEX2IKS11a/PHHkzqNmCx9+saHSPbzv
8d/SNz2Pr23l2M+YEsPux+uq6ambe2HFyTEKNYNvHNzyVfYH5B3W0LQT5SDn0qdB4we1JnOwoWVa
lX/e/ciGNDSFNrKxdxgUaqZ9ad72qGMJg2kMOs7lgm2eiPBC2abnJ85fr+8LTVjhFiCB01Ktr7av
DMXmneLvKpDYyBGj4wsS4s2V10KoiStoEV++9/ds4uConU8HqGGs8qjbsb58W+P6AliJ87wYwuAI
PVUiuPZFqU3tF0jfp7JT8LkdZp0TFjr6xyz1O5S/1DIrGl/yPeyhlbsP+D+ZdYzwTATbjDUz7l/A
2/H6GdmP+hTHU018Nan0XP0C+AbvjXithq8W7PPDGVgpJ9cInb3KE4PpJu5hOiqF6+tROWBbhlPs
ttXllIGDr3cswaTovSuf0sqwiSXLdqW0MutxEXXl0zH0Nql0NIETLpCHy6g9tzIXt9bbgvp2ydXa
ajdnZNpEMezp4SvcgGCPf0ut2I7NRRjvhtL3WSVUUtXY1F/QxmAuoKoI95eShRmqRc9ZMfpFNl7S
KrrViNpoBXch6uzHF72101NrP28uT6kKxeOVwjncvtpN7jcKqgGZJXcmfuY+Es0ldK7QeEd+i25i
bZcT82y99BjEqX9jOomGIkIYo9wR2vlj7GNIGmrj7Dn+3NMJvB4duLX4+jr7j9v0AguU5uu4ttO3
DaqxEMgI6/Db/WKf8EG7TW0smo8p2PNvHD40FSpf9Qoae2azYiv7F4meaMpEPW30/yzsEiKjgnst
KrafPmTd+nKQPUIx6mWde3WgvfXPuiyUjeT/NKOovRyp0tXkcBrJQbuMcVVOfwSAm4h4P93IIn/s
du4fNA0gmcrPZ7kGRMGmWq3w2mHok7QIHh7ETeSv5Si4sIFKelTx5nDP5sx0N2t9DskDa50Ri6K5
tbfbzX5Gqywh+MDMaxbvUQVW06xSdRbnXNCfISbezk4FXpDgEocC3N+HFh7Txj4KaIvjQnMALvJV
mmZ2dEm7SsEmHFQmJPL870nsiypqxBfIkqAtfdpLW9N1tNjAQVYd2CSuiXNnnnh8J/QeJtmXCP6w
7VVnk4Z06pbI7RR+hS1obustr9u+cY+GoDgFXLfxmpIOJiFkTh+p0aLiAuH/UqxON+saWrc1b7kY
3mM+g/U+q+2HbQSq/+6Et/Drcjjupy+1zUC8/zk3CYYXFM7SlvXu0u/ZK4Frpoj66oihPhdypQIL
o9T7yzakTZqAHwMJyY65ScwWBtaWnsvpXGX3vqZXnc82v6japcQtZMx3j6urHM7WuP/JxRklfeHG
wzBoEzJ2xWPctEbPSCwAZGq3WoCaQ09jcDnN5PYAX/NO6IWbA4nx90o7fHaCZA3NdwehEk3NFPd8
7ezr+BueeZAIL5vzKYadGK4DKTgb+gnzI70kv06ZVPNtOqUb8Y0ldI8saRZEswTWoWC9d++IEV2s
L57ftCnq3t2b0iuAj3FKKzs9tu4k5tzkRfcRc9ePEJg/eVNF5Ipvl7F4uyDwTMSNpfRGgGifmKuc
gUzIBr/eYZtPjlHPlZID3frhS/mD7LXdVQZNxucnFLjy7V+lEk/vmcG+iA3XEg9EjSUmfXb4hdcC
VYUMgvY31Eir5Fy06vYCapSz5NGT9BXWVrTiaTpIMvFi2khQwFHkDmp6IJTnfIop6HsQHqzGmSzp
aIEb7cYZEjLO9x1n3aIJ1b8DNOyRmtMp+usI1v9MSsh+1M36WTrp4ecyzxVgimQxelcdN6VAcvb+
rmtZ5GG7FireiHZ+lxY/ft+dJZ2vT4VgRtE1+o2sluUZlbEiwIdxuLpJ8vdPyrUZa5v9yUnnFkP9
fPfpESzUwKWus6xzPQwRJHXeDp/D8TU57z4w5NVsiAi2EbPUuWcOpViQsLHYnLn9DyJTJKzG1vij
yZ06XUZ1qgbgYeibMYRxTaM7yIJ1UULRI/wfNIeKAgp93jDwTFCcgrwv/nrkZY41nWyTRtyUXXWh
iSfwuqQU2rpf9T4/cqikndXOaC/CFRE0jzpZnIB3fhrT3TmPxKH2TKO98S9fNpI8RIx3jT7cGEvP
qEEm2JkxRHwUu13c3jQil2JxXzyOSzMP5R29NV1eurONG6CGVwrEkCNL2O+bwyqEUjajP2A3La2j
fLbXpxEoY2FrzTS7ZGGduEybFJ6HMNpz2sg7mOzG3zpstTIBA2LgVuFtWEGijnqNL5PSGddBUyLt
9fyj48BqdgMgBA6mRmS/hcFOJjuzkzxRFvEJqkBJ3J/+EkGYNzMxjC5wjfk+HZ/WMKXAmS21Niv2
n83YZh9vCRKAXXRKHWHOWYgT4gEZEv1+V8jmzctkSF8eMwIkHTTWyrKB2D/5Lz6igTk2I+B5jxO5
qLenYMI67npwQWHTxm3FytABB1VB50Sukz2/sUDHLGOSzl5JKx+JwV8JNTUVgMUr+zCZ/azoZrLd
JJofjYaBe/Mf71sN+IYk+FMhkmMpStjFvu21I5kqSyIGKUoI9mh2LI/Kvf9DVr3WYH0F0RzQe1T4
PFK9IUoUmdeSN7pXxvCGhsOzn5scjJ6binWkBSEm3xDzI0c6W4fTzYivJXFKc6YEi5WKrppXXp+c
BS4iWcrCarduGqV0H1vM6B78j3y1BOb4iK2O+s2qrsSAoHeRDc2yaMBGlAy2SGv5kZco1rHEBmVf
6RH2AbdM1x43FKc7Ers6STT06V963b7MN632jhv8tdTT8idPC1rxLwzUFlpJZS9DZYtPXiHe37bl
Qc+BHPIIYOp8c2TxpGAj1CyVyyhnR3o2Hh5nhiax4p+TWNAKx4lahJMBJWmUc5drXcAha/TtMfbV
EwzK3ZVEXGVmt+ql09gjLLi8K2AE7ttRIQ4V0pXGm9sjAiGP0n0gnALNgyfQp7hWpy9JjfvvCADV
xEM9RUw06oHit0EcfeWeCGm7rB2dnd3adxzrOZypTR1oYkqSd2++NV7WP31PQgIgPfH1hgcXdAE7
RKIsW5Ko2b9d4pDRQAeMkaX9JaoHbObwCQrwPtpPMj5Xfz4gYg0ksvuZmoLijErMP7KOPYHIxmJu
8ieCki86hOHwxE8BdKUPEUuKJ9xAeLnKkInaLAAd5J41nHgAuS8Urm5xk3WIWTS99mmjdtfy5sN+
SgTYRk7YCbxh7OR3/vMqfxva24Tn0dwoNGTWnO/VZaFqaEDWzHkXJNbUFjOo0MCSG5MDSnMF8r4o
M2IpV2KSeykTwsugqxz00UlQ2CS5I3TUFfJDPoAJSFEefI86Oj9xcuRZYGZXXS2NRodRf9u8jtSI
wBXfzfl0K5ouOrgopFdc3mnSADUHmQ0D/9w+35DkYOTU27JOxjNQn0Tb2eEZLLKUR25Q2um3Vvum
OcmfvnsaqHch7uMHIYWBZDEiHNV94DzhVCFfxx/RURctayZcQB4wDwhFt2jAH0AS+UNCxghUACzc
VMo07qQXeLSiXtBqFrdJPt1JPu3Qq56H6q6+bVxSpghG5oFrnkH1v/xPGCZ/l7r1POBVd6SJdUty
bo/i67sov2ShVH7rSnkW6hwsq5mCJUlLQDQWgyq/xTohJEHDd/WVZBeWfuclKrgB5ddZgvDnSCDI
NJUbAg6IBOag/dpbq2nnJiHnrMlSqxuxuD0ClVopWL5kLhG0Xl3PMcmGXEncustYXrRj2o/JCDgq
5frs/u9CSW5ws53sgvT52M48eMTthfMzRzyP+ZHyiQKtYIRSj9TEoFBCG3kxgQarSUktWW1WXsaa
dQ9UP/u412XwEXu9Z6yFcAkawCTN+aIXC6EH+XfAKR5xdNmxioF8mnekFW9B5nceQM8GT2g7N97K
+2IBWwG3KiOSZwP35/NER174ba/xyE8zCtWXfdqPzyeAyrZFDKdLShMGomO1nMq9XRC5LfkVz1L4
aQSAF9c+wzo/NVNPMk6ayJfOSZwyUiK4NbwsMtSsuJ0tvtvnTE/1ufswuBNA5gK9Cxd5mwTHYjX2
hRxyA0XDLMpmDdv8qwZCIOX3ZXSWMDj9+PK7VZnn1Bnuo4Hn+0HqW78GanV0KEXORKm/z1M9GVT7
cdu9HFEECiiuMFvKnnZUS23+hI0G6l0okhSi5sfiKjr0HW4Cq+7sEMuGFVOk3+2A1TMlUiDUncZv
meCEsujcv3l1vUcRZ/cv3h45GsrhGWeALghfdEJ2wrpZhdCu568Q+8+Mrg/esqPit2nh4a0WSAR+
zqO4XrbOv3QzJNvf4ndpftim9rgXw3aTVRv6KUe6e2iVLVpxwdT18PoF8ned/7jh0NuqzMvCMxm7
RmhDgoccua8z78qa/ozhbsfFi6/vDrokX6YnQTtZVJa/EDt4gNzQavHDCZXlvR5fSOStbrFOyfCV
0ZUiKI7yH4CvNUYo34ExQa6as0vnVUiL/7MXazTdowh9HCXAIimmaR7JcYn8SRiDjPjpzOXbuuL2
ETunNxtit1gsp2BzNmXPxq8su/o6+6S7UbLFHAqRIt3puQmOkiiXP7fAgdjJYHpZJ3eoStIl/ic3
ln79Auh4Zzps662XriReizOh/VmwHYqMmta30F+arCSJw+3mXBMJ6XI1IDfxERudK2oiCI2hw+wv
QUq83eWdmaZd6x+IOlKw6tVuA6COgDgnAX/qZQ5LwBuWVwVNNYpjWFKuObOC/ca/FFLSSgK+uW7F
Df1d/JWgOT0X8FwIjAt590hODP4Nv9yn02/utUYeGzIpW0H28Y6cSfCW1qufRgcZEjyvwUlVUXLo
oPRykE1BFaDNS+xWX/c43qNm/D2YH/G2bNgOugFkP96ioMs4kdG453EMsRlp16XJutXz6r5whi+U
t9/FOpY/wo12jDibdfG7Pjk8gJs8V+xktud+TyFGws2uB2d65CH17YyA+U9Aba4ZhwLf6cnnoKbP
n3zfsUmLfoJhWrcTYk13p7DvWtH/a0Xwa5VPpv15DYRe+lSYfKmYZezindAyXbGBWGRnR513u5Vh
Dhbwt1tkidcUGyOQnje+I/BKSs9WGQRRJ2L034VRPhMr7MwKglEP0NLhVyS1NTobsCkbaCYKv20N
331qnRUB5cXyVJtnTENZIzif1bIJ6L8Soiv6CkM5Cbb7B6NJk8JtNM6BfIvaSPpnNnqSBtG11YO8
M4GMXdN0sxPM5PNdj87hhyIkbmaq60PxMg64DSC+35Y72SZ1+sKJq3gqjJ3SZhQ0KAkqMIHfjEaH
v26zCNFqQ0yr5APtogDT4Z2KR1vKxHCGGcCWuPCeQCzMTsFwg/P9RWkNsFMJlKofSOHCsKB3/rJ6
yhcOplcSjfyGmDbnvXUzrxMdG/26zCXz1G13Wue0u0dh4pcbLuxdhB+vVLYONDxKHQ4xMZK12yGs
Hzfm1K9TJUoxYUNWG8c3vKd4viZlNSynBBTA9ui7luHFedUVg0ae7gwkH+o1XU0xN9sWeM66tC8o
8HIl1mZoPP2NZqDP9u2ErZtuETvUlnQRRMFcIv4TnfR1kqeaUjM7GomCEEk0aZJal3i3T5tkteSH
XTQ5bhgVYHUbt40dvbwvpBoiB2CvEG8yGXnHJiXq1b11GtMgeNLJiWFcztZwMzA2H1aZ9LrUa7I8
YihjKW2Mxb0GYuzIP/GyM3xykHEjvNT3OsGVm5/pw3PsEyQ7c/Houwwfpd2VQHhBJtJbYQA49cso
geyHwXZtQX53oT51nUfcbshxX8q9fO6FO+H4I01eierQ6p+aOrI7cV1xo3aXCff4yiCYXQBbKGOZ
dqr0NeeTUp9zlsYQDeZFb2RFZ08dgwMeFnizfNUEMZ1gRp0B8HYjNYe1VBXFwWOmu+z1olGxRNU7
izB8MbeCNOMFuoKaLabjdtIQsEtflsCAVZPG8/snaVRlCisyKasaPXPJcv3XXBO3utCOEoTnOlDU
ud8mH8LNrkNCqUAlXJLFEtJAN65JvhExkbeyu/Wgw92/460KE4VhD5iqtBNKjas28vRI8fsMymkl
CIpp7hOW77ceydfBY6TkCvDXS85m8og10erU6a//DESCgYN2YeJlqRnHESJcNjakTaXZ73mkT81x
rg6+R4P7kICxm5GfbEhPB59opn+wlM0x4bsVGjhx1ZCARTMSE4owSuty8vh1yhZ4Ctx6bRrxBL1f
AxV/ONO/qkL0tmzWAVhLbKIPeTCVaeSScCXq6gF8NcbJl5ZvDBQ1Jgr64IU9GvoH0UiouWo3yzwW
2137sp5s+Ar+Ig7fRrx4L4lMo2B41pIxxb3OSr14a6+2Io65DgCTPjMNZqKm3FTcSeXiSJVijB+i
W8diabRN7+TFwPs1wvUUxcOdMTfPk4hlEIWgUN3YihwbO7U4tULDHXWrffi85FsSy+KEeBqY/F6Y
pP6CDTcsZrdeZMJ5jUquN6lyz0+nqhsVQPc4rzLi+Z00z+aCN7CD6gpChlPPmVbw/RweiTh50hwq
VqjmWFA5qUN/98PUP2t4mLeJjgbK6380J4Rhv6huZrXhbU0jYwWCLsicVnoc7fgEasKH7PZ94xg1
FCXgVBJHL7Z+yAx0UmOIlKN0B4MwAoDe3zae8RHj0AcX+9P4DzURD1TB6JZ9Eqh29veFQ2Qz4C5C
TzExI28HO5cCNpXW4xGhSRX9w05qStmkSGosGl318U5IHSOL/mhNdj3YAtmNYims1NRsc3R0yLmB
rCWi5mpnEh2KLSzKr/NOI59zJDLqX5ApW2JJb41ZKagVX/MAGiowR+qjIh0iDkGBSMuO7K5FGZ6r
sBDg/w4Hw22croA1pYV9vStA3U8EzhQAawi2ao/7bMiwaRtE4gBWJbmFrMuqpIEYSXnLcWJNokCZ
GVyHQEBQyV0OgSlcRowh8nsrlNPssvwmHKeJjbagsRrKsNVVUYRpZrxm6g0VBQR0AUZUJXcBh9FF
bFZXhWNjB5si2fpum/5v9ymSkYdjrFtgt08aiSRpzpersrUQX2ygv+I2OgW/4CxW49bIZxJSfKDb
ciceDLu3kRG3LjrYXSabvGQ6PPc07p2mR2as1Fs6LSBkCX10C47FmDva8lcVB2JkAAarDwgSrmzz
499RvkmscR9h2RXooMZV6h4W4hrvp0LJKoOTTauqpliOnVzeInguXsRUWgOHztn4UhW77v4EBi9g
Ik9RznanH4OmDdz52GDVfomtk+2MRJlR9Bg3Sk7SCIpwQa7tYS2kLmZOLon/hSfXiyzdsr/5ofxM
CR1kDFr+vgXQEYvM8MndfYp31n8vMM5rJadvSGQyh14EMX8b4mD7r4IXpNSmZnuHLT8XENMW2Iki
pbRbXYRhXFfMNra4WdRa2fA94z2gy1eNFbHEu2cbtP6WjWi47GSDkj/vrUvAcGfGtDwDsTTirPR8
KqUJszOhWHj7213on5LHc3+CGOO1b4ppfPYD0WTGd5OuDpiu8xSIYxDiLjvHDdlVvsCF7t5dED31
7ZaGIX0zlkT00bnahtruxkNbgo9pqjj2Yx2HDcTf++wcdh0OvA89+Z43wh4Pae7F9gI0xsN3WYs7
6MDSd8lf6KTtdQC8UWFySQssyV+VWGv5KGS3IifZdgWwxNUZQnbOGIQth09+wWRRLTJ/xYMJK4wK
jAEeuXH/DGtv9C/bb+us4TjU4mCJ6zXA6kfdZtxMVLeVTeu5JEHqrfr+E62H16Txi5N6wMiR7hkk
0c7ChCsmMjy44Do8l+PJWb5Wmv8sxlO3hfPnSGdjnZBY3fQ/iqhXrtj/iO9HONCuSpgYpgM+cOUd
xGAi6XOcJ7ONsHJ8EYmW83sEs15vXJc0W1WvWQKcBP0ZE/mCnFXnxaWLVHc/6NXPH0nyzJPELl8c
MXOmODwkclfdMIvxL/sQBhiZPfmId+ZBJMeX7cg3NWampATxLYUvHvPmLcRP1ZCBWfUGrVjd6gnL
FNzamrA4t+G6z1fnwCNxiDMmNeDaGbGoIchxDgg2+4EanreueFYI4jozTlc9dpEOLW6q5sH6K0gU
3xxGzpuds7fTd1HIHonv8pSBAWsKV9Mxh4FuuI6A22xQlS+L0b81qkMyLoUZnFusySuKsy/+b489
5SBDwBilYw4Ir1x8nZ3Qc/rF3u+PA9CIl8hepVI5mqA3lPVSLiXUEb5pmFUM2tvSb5rkJzrKjR1D
s3nhkKW71Nrjko/13eNsW9gtlrCzro3qNVcCxCjv0uTtZEBvDjsnfmkrE8/ASrKXdULav1LBRxgR
UQ5VRQFoESRvsOW4dmT7F8wcghyHhN4IAwhN3+eTc2RjLpyC/rBseR4UwGpV2oGkKYwQWE9uG5Ie
K/2Do9VAEgeFKdfiy7Xr3UJVDNaSMEd2DXPJLuqHHKNnlwG0lIbNI+C/p2n1D4Vb+e4l99B4MtcJ
kb8oXZT13mQ1T2jCVC+CLjF9gTK+EDee9OIkWFy5QpJHV84Zpfpl2aKKW3aWA0ZW5YNvHaIl8Ff9
/GmRZEDSjdjQI6CufIZiTJNDBVlB8tbUZWCVAy2mBtCjxDP4kWle58JhijQXqAam9Gx76nRXkYvs
R/PlZl4yS0i7yFF8RFfPYLSeXulGshvNXLCSqornk+2OOV5RU2TGQ3F87dF6LD/HecrpVoH0ZsPd
pteTYd+rlJUCogi4QEidGAcqLPm2zue3qq0i7Q99Cf5x8nJhpbSoVmCCib56bGquM/pfeTSEHcuZ
e0ba1SDaB7PUp3qsek21fsaIu4FXEYD82VJsx7fagF1BHWIfI4Hg8kNT95z9W1Epl7OzYNc/PXEo
ubIQ5adVAohLCNoDzXxkfV9Ya/HjFfI86N/FerLoLWa5GAGSn4vNng4H5/v6e8Lp+8VtsEox8iyl
lVXIj1i5aDW5mCYg/3IBzTt0Ha7p2PRtfI8dvl0zPBLwYXeEhJdorh0DNWYqAN+UNxTdsq0Cu0v5
T1Az0TPlfKk5pKBMWwRjp2C+4tBJKM4qK4MD+D8Ol3jKvKngN6PVe4bzwJPlIAWRdQS++VAGc7bg
dbG5xy8r23NmsjttOnd+Z4zNx2fxzEhb9gnMIuz1TnM1j18KYekdWIahYcLaHE32fVXWDrjsjB8C
FiNWs6/MbumcNnkvkLY5rUbk5SZm36c7Xaa46WeuhLavcCiGaV4krnzhnujlE01T/kMhe7jtsgg4
z8htH93QposB0k/O+qZBu5NanVr9y6D/tJtXTjRCNZwbYglfRmceds2nKuDnoysUHOXbNh8w++bw
rR0y64X/ZcaNn03/J0LGRiCi9K1Y3EvP8qlOlgjCuJSfTG0f1aJ4wa43uUfLtGZ+Yme0HNdOmq5S
UHm/gNF3WAoJ7XnIk4laMBnBtp1lf8Y7pgMt7brsXATmcicqk/xpdVi4MZLgmoFnkeQcHdrf4MAM
1P8pc6R3fEfeoHLXuINkdOimQS1948nK27xc/ajmBumwjRXkM8v9H+droxsI/6nJ776MMiMrnN+w
CcYAvfiXhQcN3tzruDiGRPXjijcc1WfBtrfIk8XM66QMP/LuhYS33erpm+Yg400nesYHSPSZvnta
6Pc/6bQTz4du4tgZ2TfI2rnVc9/TrO3eqmr2CI5sk02KwOH+MsjKi03u8Q4EPZY+ni14arCG8rmk
rXbOJLpZls6m903NiFW9DBT4NRjRe5t1oZVRlHOM97p98fb+6sKp0CvUu1utgFf7FN9mEKOgfP0z
dziqCLL8YvGDlhfWdWHkWzZCflSJaDGI849BQZD7cpJ6q6KA4DUTYFAmHc1IaAS21ynZrWNEUnU2
FiDwNOGYT107pfUdlQZhfa9pTgWSeZvwNr+RBX4jEnngQQDefugzDIPaOBqy4E0Nz4lpFjy1Y/hO
i+xtsGdTl+Ae1bbXAwqZRv9/KkHz78924sE9dPpTjNqPR3sCkAta6+T3MBOPyRltsuYoPK6Fbq1F
aP8yEL61PDpx0DSrdSqoViTZBKPQ4cPMKeNA1G0TeGz4RFohdpAtbSM3SGzAWv7+P1AITJnLwz6K
7TpNMRdz7qrMVClqTXWyrPQIiu9zMTe2Sg7zyE1nLBCV+Wz6LKRU9V9rpcdX3+wO5PtZnAvpzuCR
nknEaWICYdE0BVTrjbTGqsvZgJOx84Y335ikeIH9dqj5xWZRyk+zQmtHcdAgivDMZEPomOqVH/2M
g4fLy22/pvF3PZ7M7Qg8dPX6L3X5FR1ZTU53DrtxtQ0lRzoPaFQYdftaXxPELC5EwKgTs6WFOAyn
UlBoVJ5Z4MFwr4B8/VZFOveMY9ipYiYiAtJM3DHfu0IQK/uKp0ED0AotmaP63OV57MlhL9BZDwtH
OMm9qkL35nsuaYZofrLVyPY6f80ZKvj9CC8aeMs8wasgtztqwj2oQe12zeTtHkErHaZtW3+r+Rl1
DYNXCc4/IqgyjzTiS64jTd0WXL8CIb5MYJIKES1hYmTQNWDl+MiI5UmelKEGOsPIH/ddgf6xUHOH
W88L6ybahq7KOjRGbnGOqXJzMx0iEwG2SJYOBaHG9lG8r/SrY9+kCGPtm8X0bBqoe2AVS5yuRG/e
tK8FTfIGIfOfO9SImRnTyxEG2erGPntf974UlZsFxN1GJ+aP5riLCizG1fJRYsp5YsQJYzbiU0Zd
cqwQbfuKgcgbKnlzKeumGD18/29yplxQ/axYqEK2Uv7K3lXAaP/kNbocmXTnoVLwxRvzXA7MXG2n
AvcGiQFjKEYyTBoKC9UcThNgXWBoaSyQI/LRJbCMNadyw8PJthdbr9iGYxBTP6ltc/Qw7+doY6CL
sYLTBDWPEbzkupjB+iPCnkNLq6KIEfS1zb7d8UQcBGz/dblaBxxTSxGU0qKAQq6C842DiG4TUdJK
/nQc0pShFP1Xh0gBntaI9x37fxVxcuH/qspt3ja7meBw+yLJTyca54O1lKs1acr5QOLfwtRtWdj4
1WWI5PmvNI+E0+WgRASqSK3vYiUKs7ZEBufFXT0AwAtyNLOlg8Cjq6L0/AwKWeYv646DWNL1OYnc
jvStEZC5FtF6I80vA8VcKeqYGnKK2q2uuAgvm1YliYVJErChBWW7YiUBZ7t71tEXAI/NU2ZF60pd
OzrxmR3bk86Y8Bdq8ZnsxKcigRQJgy2SRqunFD+hpMel9OVZzXxbRy4ZZu0n3XHdSUnvtp4JPB2G
ZYGQkfojXC6U2nmRwDXA39394k+FKx7QobeNb4DXlmEjKCu2dGfXGEYbnUnC2JvzbARZyd9x1vdP
XarERNGfOoCuc82dRuRWo0nDVhWm4Rj1QQpaz5HS2VVnlpAaC295k/CdZ9TChbex0VTpDdc4MR2Q
Ss9vGudryc+7tq81I4SpgW0gOfcNJu75wMORXec7QRZ/HEwDDHBAgPcGtXW8vY0dapYqASuxasyh
BcXTv9c+OxcUD9ZpYddIwfeOZmmDnzxlrTyz1rQAe8sHad5pJ+NZnm9GiAfILG1K9pt0FU7t7LGI
TmLY0HQ/qZRkFDMzcbroSv0x/Nx5jyqchnj+Xt2vrRXVjkV7wCW2JqSpv3stO21saujrGukzdyG+
ZorneP+OptF3P40lU6b4rSqt3dBLu59JLlJjwzNGc6n6Pe+UbG/aP8I+AFKqnWtKjSgyGh0sji4w
wmdNvdyQBr7tGYdtNMcFA+fNYWQH98ITCWjEnli57hl6dHsiYnQ0KjCbp27yaHlYrM9cLHBmLkue
aHAlMr+Ejaszt5kAX9Nusrh3pgBRiELWBl2bAzQJ6QiA/uxJIfKeNied8dt/rQG7nG70p7BkyJSo
ocMk9hL0n8GNpDzG1FW1j/CTvYX1FQLF1PvpEx4kgDYPxFbFVjf7fstcJ2HRFhZm9jMYpXla7ezc
m16Vl6DVt+No2nce/CWY4CtBxQ6GVg+qDOmksfpm1jH06CKSPtMMjPVpmusIa4Dnw3JME4LN+IvY
ikAGJNRLqpjkOgiI2GxykhNLAbkbA8kp10yCaXiUbrNyWwR7PblgrqwbLdHJtkePbKXpyfUsC8Zi
xVhJeSKSwpJzRpC93lYJ4S41Oa48W5hIAq/pH4Z9uI81RZgPWQgg5/vBvcEo08bVFm4COAHHV4pM
NeBXkOIuKK6idewU7dgtlBEUVaNRoa+wMKki595z6n0L21UYaQ9oICSaEthMHYR4b7+VjxK6/G5L
Ika2GBPD+WCzxKT5oCr7Qy10R0q6otOXmWZscwcWpdRrxxz0Rrvdkv3RVJfk8OPqN7exf5cW4uNR
xX87Hm4BvSrKtlkAd0vF0OPmBALOKvxASvORnh9kJ/6sSPFPn2MylbFWMAH9p/JMKx4XnjfGdcFb
PdG1FzyfMd5ra6O7bxVVjdTTbuCvoO50kGm6g6bnbIGgeBIjh1CAavNpDwxpx6x7/Nyc4+WPpvlu
90pVkcnmypeoeUFqzlULFfQBNrEYoJ9jZVe5qw8Aqq34P1I/SxOPUVQzVwGqyLsi7ayWD54ZZi/r
dCJHThmQ2GWa3CrvHVL0Dt9FuGB4c1Y7VlDNNMokRJFFvlE1Q0cC+7HnmNmLDfxjlYJYsMSNRyJL
CKoFhpK0OAYmKR575QOFa1AAEirb/HTN7oCQePfKTqoqcH5O7XPtmUL1bxLUoNIjdecYK4yE+GRy
TD834IwQAfna3nxSq/OvtXw6PUuB+KQmkH3Rm90CoYibb/azUUcOh9SNgEdZ09rcD8ZZHTQxyF2R
h4sRokgcyLJhzd+rSXOqDFUUMeUo6O8KWSN+JxgkbG8eR0mcyVJPgfDRJ+PP8+5YC1makLptiFO8
Pd1/FOlQWNsaWm6UeVSCAcBZ3HMzO4avJ5K3LBPLat9VqVIuFHw9+ZhaTl7WCntLBWXkRcIyZK91
d5nOgstGDoek1Cbrdn04FabagJZt1a66UxEn1u8Kt0CTudqUhPTL5xt1bHy16N+z4I7xAvdyOqNV
j0GLhw1jhgqmvRWbF2/zyRqIGCanDBlckCV048SZ0VqrVLta5xSilN4Gw4iR027qruSBljZhob5H
heGp46Vc/Ta/cA+8OmYYH9c8ByVE0Wt1wRkJ67rR9bP45KSmK8vGvvdtxp33Umv1l03SBAafFsYq
BBOn2EQjj+NAT1PDdFiVmk4Hpz29IC4By6UuO1ZClsiF8+5ahE1ESthXGfIPsM0mP+o++BmynkZb
YGAwPm9asfWkD+htXM9Jxnq2+AozhvKWlPn6IlZik5+Tbri4gONS9Qw6dAk/4a+JPrD6RelmKT8H
wVAn/Hw0VjEKkcZqinu+aAyQKDGWdl8eupBWCI78l2MstOdjfqcM4AzjgsUGve6LBJcEm7/Vppjq
zWPx1+y5G+49pAV25l7uWqrGPvEvt8qmZ9a2//iaP+gfzbBGbobWUFaWowR3YwJbciOJyGa4mtq1
BUSM1/+mRSYDPuIwryIf+UEK5qVkXgxrMXMtxRj0AVOPMbmMmlZVp66iq12mcYqAo2Ms45DUL2dq
P1h2GD/H+6V97AhXBDFAaKT6uNaTOZGrPx3dIS4RDJGBaKzJdkpLkuXrXOlkgI48X8XQT/j8lRz6
gT7lJFAbkWBAL6tKmSQ7lyU0qu/sBC2U+Im8TuigrHBR0PWNO2F4dgml3gDCVAkjJzySisKAqSO0
4pZUB44aHcSEX0KACqxEOmjDcT65aTF4M6Gc2QBMseq+3KDuLftirq0d7Fzjet+m+h2/ItfZVv4W
nPnpMPb6t01aB6U1osMI1vOAe4OwmLIEhbg5vduqPONdRfdkg8EaA9VqwMa1crV0hXOCISrJCPBM
0raxHGoWgOiLrhipyjkIwngJHHKhsk1uAR7iC0WESptxUZaoZrpwD6zH1AmRwVwOkHUAjGwqZL7c
TAXjXvJ5GYstH0VlN8jv4azoJCmU4puN6mei1sPWQbl4wIhkGoJyYQ0Sy90lRBnBwF9LKJrW9drj
2LGqZmoYkYTuOUgP1s20+XOtjUjJEc2hNOucGd0SGut8GR1ej/oHpx5JUGZAbzBS2VRRtkEH2wu3
mvv4rwxuYsF3dVIfd3B3kfuXquLfOU/TRVhYjD+zRSmDcxMfG5OEFTi2I6sgu8XAY+Pb95+MRsLl
HWjAqnQKOmpZE0Xyj2ppYOc/A571MkMV+VSNeUUW99Lyl7HX6zR6/BQdv4u5jlvCrwWaXIbK0jbB
baqd4Lk4+kF2Efl9SMrSIp0rYtdQPqjuW7AEuyCK1raB/mPCahuCOm/atJIwCsOd/uvirKOAa9CC
vbyX46jlLsn4owSwmb8XEG+0yx99Bkt//llLoWJ0Da0HO29R2VcCYmfB/vK+QQHkplsMcMDGP0ue
eURVc4uM4T1KTivIAAzVjYJcMspgL83MNhPwnIS5V173fz1m290YS2KLrWJQeWtlrRrQcLW5HBHM
tyCJWnRoOpBvj3SNAaMWCij4m/OLn+cV/DsRD/tykNnkdNOOxmP0eElcIGW7RYyjC4+CxIYvrSNJ
5vkgHyVyrUmGK2ohNTwsOyZx/EPI2FB365A4uFrm77FfqQDoG4+N7Rvv6YtW5fEcZJKuh/p3t2te
x7ohP/wrekSBUpiFqHuvt3aRCkWA652kkgiFf21oBCSfaZDzju553LfXufKkXgj6t8Un0B4IRBMx
vJHZc7OPlcvCJQTXfbQ2TsKw59D+rALFWoj89WJfiWVVfbyLKttsGNSYmQHNbcOmZka/LicQ/lGV
LOcdiCXMaArSYtBwyo1Km6ra5+QuocRQSbO6GbdLOAa3RDfu/Ju4UmsLvimFgumGdrUDRE6oPXsy
RhiKMO+XC8KyYq51Cd3YLifrWgLvy4Q/iy8OUuw7Q3p+91AyjQMIEyVdJyxHMgvZ58F/7dntQ/qv
Y6WvWyGDMWlPIBeqB0J+vh2xyuN/MXVaoiTyd+pt0bFA2oIsHhmtYCMJk8r+DI/R00AVnDOaNyIS
49imkRR3aZmtMryVQh6H9zrVXP9uH0BBDySCK+zKrpDmInYcE3EGfX8UAGdGpDf7WMV2tPI70SjU
GZf3wC/fb/KPMis+rHSnqTcqAABp8xRwVtRqOhq7SJxTOXDQo2eK1/35QvpoQskhHWBz4xo/CuqL
HMIC5OZkLQcVDjwCXWQ0LzQ6BiRh2AaUZvR85zdAfvNdIL79havubog7GownhF37/PiQZkPXzBq4
gp+uRM/zzkxNn+xXBNvBnZl73tj24KRDb1+Jy6ZG/VS8vBpzVSBjoqsauwzlZzM190MNiyZIRAjz
nrbqMoCYWAMMDxpazdyJ4xUAirLdM71wH+S1thH1DUxFrrsO/nhiyAfJgi+pY+wbNKZar8ddS6Gc
ZNRltZKS7LGzIdtnYME3QZ3YdzCJfDmrXCm3MOATyqERsLE3OinrSl9RiQYmYYXcud36po+SoCyE
cW4SNBtEtfgfWEY/6nAYPCYh6yKSDngnI6CyKFJCnlYVlm3jSwBcyw7YC+n3pKnjdODGx2zxPDAQ
oKIyd18uHh9a0A8MUtBktZz0X87uuZLfOaK5+wasYhBRZ7E4yO6DYkrP5EQEP2MJr9iKthGVAifI
KA5GVvQkxUlChtElRVvPgrp8pJAk/dTyWZ1tDWui4LsTVroIIiglyk1Uz6eX/JXIelZlN1MQHImP
M22+gdWx5dCshtdkNjeSofxGjV6Mlzmns8xumd2on9tL4khHoWnAP5Cqib7frKekFjoKKz0zJt4H
2Lp6rIyv8/VR97sqGUP5HYXExJrENO32XJ751M8rBkxXlmGlIRvwrpMWIhscgX5ZWPusOqPPCeWs
GEwU7gDmkn1R3qk63RphTeVyf3Wk10bJIpPLlmospI6LqH/lEoM2uIern05WgPw1ZZCtkAyZt8eR
bqtJgwF+R8e74wpU1NFHi8KTE2geD744kgclzxPIsuJqnx3f9Nw5KXrS2B4GsxKzQBMjtmf1zAbY
wiI7YsBa1vWbU+m9ExSxhE/xgBIqB14ZvHFqEthCPat6hfFhZzu6in/2xNGSfJvXlwT9FGufPlL6
Q9Fs/PCk48rcnzBRbQOP+DdsgOniHtGUUQ8OwyRBe2FCgZGsfnsOHV/IKVsXpPGGikk8CaRthspp
yEieshNOohoK6CJkdteEq9sQZRM7Ny4SyRJ6wHwqXBacfWL4bPDHMdLOY46NHtcKoVkClzXpY7o1
sy6jzM2YBcK8eqfK59rQmPL6tZusLPtkRQCvnumH0cyKVGE+cXyeyB1BPwXhWb5l/8sLxMcezmFd
+3Q0YKzC3AKM/xfleJrAGQr0iekg2/p+GYcEwZAy1+rzmAtHaG8aOhi+26682A6DwGU/yJ+Y7Cj4
Yx5HZ7/F0gQRC52eJIr04IUO+Q76g5M3CCdSPBpQiISsPrhwVfo88uOToVvTW96EIbNZWr9XYNtn
XOkWEygw5bIIHJIbNwhw1XApvNvLgUH/0383h/s3+e7tceC5VVMeLRLKq39R1EpTbmF0WqCLZABR
tzuwqg47T4H9k+YrcglRJuJdc/7F12C6mIAYI661dEUHB5MgxuEcFAInOPqM9QHTe+7G0n1Jvm2E
uwDjq1FFAvkvHO8gpfyIBQqmiGrCkpiHyXJ2IEw/0ldIuMiCpiNpTzepY616Mm6qoPcN0YcTYRYv
1su6B1wHHRi9fIzzFYxqf/cZDx71pTXQTwpMPVG8hbBh0nfHzQVndVsYQ+paLdUWm7sTFAtPxczi
GIchWzoSyomZwx0kJm1yFrGuLMzsCv66LFwc4YI8bl4cXptAMzv91Gr+n1Y4KUlvDEQ54uCc2nic
95uRRSjg5H/6ehfXG5v3JQzZggtEYpoDJhCYqUJ2/RyIFlKcr61JaleTC8kZadLS+WfpJqblKvXX
m6N70yCVJL7cKI6MZmQKYdSNrDOpTyrdsp64CJQDMzxAgJFegGE2Z2YAjDib9VquKJxdklwxBNe2
K/pyM4UyjWfDbZZ+jFCooo11In3Sj5vtN3FguvB/mue8MrVcc/r+wu9ORXym/hrGlFau7ww2oTWQ
hZSkBhTrv6vv75osM3H1xEpkUY04vqLYlk632iXbWCkoOvMUn7bZb51/y/fHmsrBRukyHPtb8Cii
u0nw9UrH7v76tfEgsgbXqE5diApgjA+Ii4iwGIYhlA7/kfKYg8um7cZY4bwteuoSwiLfSZjBoRIf
f9eV/RY4oNlbdYbBGthyR86nBxF3RbHlgTlxdySoUf2QHBbMVCGJKksmAcTMNcaFGZT8SpvYOxl+
gHsioJcIA2avLUnfUq/dEXgr0jz0FFVjj3eMR5saQAFo3XFCl42kwjw6KuBcV8ao+saNXKRf2dml
d2mkB4+70tpl+PyEFMz0ByFgcrAwM6a6CMgVKuJjI6Q4YPbUplHFC+TLw7Mj+VU/rYVISLbZmbTt
Vj4U5mwEm/e7f9ihqw/2Mk+VAThYa58o3eTptaXKb6VYO06TBojZOSN0c4/mM2jDIACqbnTBs/pJ
se9nNbWAxidH9KFT1pl0tKuph3VBcF0qREVyBZeOXWnmIfFIhiaTjimlirQzbA88/0XMz6TtHAEU
BQ+zckw/X8NFXg5CZzoeKf77azkMhpk19akQ9uaE02A4LrONORSOScYZFwYH7SOwjZwp3EuC8+nu
bP0Tyg808raurUlPIuLi5IEMDwyulodnADEttd2kl4AWysQUjvJTU4KATOjdXntcQVUsRCDoOkhK
IZQ02NL99p4s+ezF+oYmRmW/eqdlS/kCuBpl9IUoSdRv8UFanY5wuTWzczYqP85EkhdQMD+m4XzZ
mVnr5FfxDz8L4ryghPmLvxxCwR+/9M7qQNSImQWuZCxoaDt5Nr9gLqfKy00kgEb0NLIYReR+9Ord
nlS+X6G8xAaqwvKd0wCbbywx4zyq5BSwibSOQhVBt0+3ulwQ8bwITseq/v7TMNnMhDWws3y0Bifn
eVgZZ+zWNdZ+0vm/9hdA+MevZY8rNsO13WV8JCLLmknzBoCwLnsqIEmObHNVgsCn5M04iUnWkgkt
L/SwuVEMS6kn0oziD0xQwXJkygOKTmfSUbLGRvq5ae7jIjEgGeAjlMA83pPN8gvkPb9M6aliXB/V
tDs1jkL3cSwHYC6ArSLkdg8kMgAyo0mThSM/Lo+T2sapwsl0fN39/bW24olreyq43AeqpIybrthx
t3i8zC3DDgSYKlAIB0VVTxqY0YGdKlDBHI2jcl0WUHZJ43GnZyyACv5SPXvI8H3DFdzPWu4lVovw
pDxwrSXA0S+aXQC5xAbusnDEy2YB7CEAXILGSfXiAbXUaay/jtvryCxUe1YsVn4k5678BjcQgLyV
pS4VCeN5UjL6d9aonr26V5Ertr5oNYU3l3Y/+KgqObPpG0DZqgH0+O3IEqufq4fa3ZfumEw2yyaG
zMgMgRDaD1wXmbkWuIxpBnvHTM+rKd+ouKAXwQwKgEtLsX3s90BmgEglWYOEna9u5GJWVOYFlHmL
CaC/yY6EE1wef1iLgxQyCCSFREFpovR63SXc1cbm+3hpIJZcEpPdDHvdECUBSfEHPa87JDlA4cLP
IPiHJ2Zy7n2En3UT6MKsjMHSDFB1BOx2y/sf5ja5WP3h1B6uLAkqoyTb7ww6mmKc3Wf1SUFXuJW0
QUzxy+6wBQT0mytcpIV4cksDSlc+ovXvbq75nyqSpdAtOQ3t5s8hSrWskZVSUTQ8MQO1beouWaM3
Vc1yimJlh79zc18lV6//uH6tDhAKKUhwYBI4nI37qCAKaQxByCQQDr1L/jmR9U4HmhNZPJns6Rkn
bKkb3d1Mcoaa60/6wqAJdJVygPNDWb9v6JZX/rWk+rDcrl+dhuJ0M2gtiU1FGn9LKsFqRpTErciU
cmuWBVp0/CVasq1/YASaV52FoJ72B7/2mxwR9MNmo0ZdUA4xgpk1Zf0sOpzfziFDXSUt6qnHfRK/
m9obDaIl1QL8KKHbP/a74qrFPS4uoZcg5aVuoF5bbuN9teMOuZVgNbwb+elcTyccr+btfrXfrAxb
HVtbZXxNyIPRYPgXJD+B5Ww3/GYqtwwN6chPe4PJXpNMQpGG6AMx6cpX891eTCgDaeZwXMskW/cM
WQtmn4UQBLTnmbhBSoyuGR7IsnYqHy8L4iAeaQUNYjAI0LucgcAnOkAtea5YYWfILRART4CwlY4u
aYaVCsr2Ktf46fMrapWVbU3Uoga5p+GJPS3TRQx2KwtsUJ1wBoKhXzbIJSedljfXlph4/PWMaIRN
9i8LzO/PkG2tvYSRUrWauBWR4+HrRI9dbKQAuMcpR99bHBZPgoqSYGUV6SFPZz0YYlR8hBjfldCw
DeH45h5kPX1pNBLCoHu54+GAESU+r9HwB8lnseUep7//7CC2x5S94GNkSwY2uBWG73eg6At0NLWB
4Rqf6cbmdPSsk5kwDKY3+0jeWURpdy7RxnhxRgCDRna7XtEsCAH7ZJuBDbPCt/wm2Y7LElGRZ4I2
8EZ+oX3TGcSgmT+/FcLepe4gAvT5s4LCPP5wSXs+RE9r4GtUXvqkrDfuU5Bs4bmM3K5Xgg28yGi4
ynvQtIpa9sc6/O0iy+OAjBG8Y2aP8uKVN6nRAY2KQYAomYJZ5+CEmJwa22B20f1O1LMWyPhxRICP
eRrY28QmHoOvK08KUlA9QhNQVG/vPqmS028C1Brh2QFhYJDvMegudGO9Vv4whMenZtOFKP5Fub0f
FedqWxRlpmZIuBiUNTjbduEBAPqyH/KEuzswYqsVvJWXIGHDKdoTjGQgEAlpGLv8FlxQQhRD2xEv
/Ytz5iSOxuAxo5IEySl7ZwRO7j6WN3aajUru69stvAkCprQk04r6K85aZz7Mn0dlhDCBibtF2REp
ZG3S2u+Glk9TM751NPbAVh3TKc6NH8DAshJNExNHARsLIBy76OFNiV1QTvDSnDDHJuTmjxEqGX01
TZXmfOroumdEfnwjUQd06mRsb2xH1LgNxzBkrrbICllJA7U5UXC5XzMWqEl388ME2AvDHkpJtaB/
ZAdf5UWzMC8zsI/8eP9V2OiQpHZrAe60/4nnwSeRB7/XA/IJZ8BzbWA4vd4sstvsJlvSQIuHgMtU
Z3TIqyvi7AkRvYwsPgZn+YTD2p0Ck/dIqZ6sChZ9So9i56tQewhsN3m6OjA7A5wpixnue2TXdhO4
yEe/x6YnIyzrghoYJdFcGR1iaBN/inlszhtTRPGNYsh/7nAUW0z7H3iT+N0kEjdGgZUcBAgOdO/7
MJMI/eDpq/YlYNlOxSFKLLBiXhIhIxwM3HviI/sOPxribvwDehMLsOG5q6F9Plyu/6WPUdvMPGQZ
pXtB6e5jim90nNFr94sIkFjacthuY13CN18gM8ShlpdK64AH21EEpOZfAM2r7BNmRNUWmsWm0oZ/
BnGXKGPZllGATVtz12qkzdYi+acowrPlu8iWfImAW5bSRpWX5bumT/WAEIO1AwQBv/aplnQxwqNX
aTDF8KFey9kAF7Ryc3+dbg5FcrGPMF5UKRowraIw3GDcHc2eDCx3mvopkVAy2fjAq8uodRbqL9pS
evYbQRBTEXtVD6BRzRuZnhbK3hswrehscLpEtZl3I3Z7T0W9Ik5VWWX0FJHd9jmanMEvxkYvUt4S
sRKZEo+a4C40DxMDVyg9zr7CJ2A+ZaEhKB254Xo+S8KsFmDef/74eDPug1bUInhbyZn9RW/n2r/2
DV97qNMRZ9JbmX0eSSrIP9noPn9jeF2Ph46yEN/wZJprXKNuFkZnwqasb2/xpf7mOa33+2Y5+l0B
EfIBlt/vu/Zn5sxrdPYqez89X7myWbES2eCEEglYOyK8R7t7BSLu+16H5vS12btBy4tKX/lMO993
d7zAbSk2oklTB697CDlp9/ACZjccxPOMypfdB4FhM5+FkL1K9pOtDoKSCKa0DUx7/z4fX2gGVGG/
PlFltNEgXv/CckOSiOTVyMiWdr8K52xXh1JHhNgvn6isC/+/U+h3h0C1AJyhTH+N4DNfid7wnU9h
xPBP8jbgjvBENtsC5zmyf6WCcHxlmzta1g6D5e/sU0Kfxfdo3FSqqB12TdXRCZ8ePssSD/UgksVl
Llm1WVn1b8qoUgVElwvVizyV6hGNxgvnTZhJaCiL3vpvIVInUO6l4Leh/01myJYAkWFHti49Yd+U
TkfNontJg68RSo08wmQzV0/TWelEqXoCI0i1YGWIwbBuPUr+ARj20A296YGr5acYschAEnoN3sdb
sfwR+Z5DrZTRCPymZep9DvirdHZON4VvGkmUZt0+148DD1oBhJaCWzJTbXvtd0jCGUKpGBDcov4s
G/gplVb2hWO3PUWipKOkV64w6ww9EU0dw5UVtLJm9s0kl4EAt1En7q4DvXKzqM0HUvABwEV1ucve
2Ec0YpwkeUTU74Ogx6CUcYKJWCNOztQWUH1Ti25gWq1h+G5032NpQ4uRf1C/O4lLlxmlorU3Q66/
bnXCuQRfW+gg9EekDfI82zRW099RtIiYYfurVI8knQlvqTK0jXfcSvA2XaYZ6ChlAa0fck/AajwS
EDm1MrMLa9MMDJh7eG0mk7Yirku9BDbatQIQ2uGK2/FGT6TrVw1MMJAX1KoiltzYz75bXqW9xbpY
yUEke8nadqcZRW1sO4x6Lw5EBM4iPXcTtEcPQ2iDPu6Ceu8CPAdow4NUxB8YgI6gTteWRgRVFCWs
JPmFkRpJGZF7WRVaApTdLDAE2RrbcOBdyMmC8RJA/V9eRxEkzn9xVYpaiYrOGqPbHap31qfDiwoE
HIPoMR6H0o1JiYi4P9DFDEjqfYcOHqwnvnDwJf0AWy8mwU1VLGebJ37FUYHE25vXZC7okt8bU3Ca
Yed6457gaxD/fp769RzdqK7ML6MPY/BjWN369cn728KsOa57QQJA+m7KWmEamPGFo3Z600XgUfL1
UXkV9S0JGWLAiM2uMkmqw3yWcv8267psXVLo40B4va/m9u2kttyMbwtkEbny8RpT7T+9/hPKLAGd
ThTdDTq9tEaIQkp52K/YI+Zb0HnNep51y2mQZDtEgHCJE5eud1EiHnCcfprlp+1EmZJqLD5TJzUp
WZkKjdRha5OW3EjK9lw7SW1JXUK3i8eOiBJQbe8QUievfSvMxoezO/wrXyHSKLa/cAoE2PilDy7E
a+QLU0R1NiptXy5cx+fUM+rLPUCEeqmMULxUnu+ClTi7Znl0g/upU8shE/WCAmSEFaQLstn0uBOr
W0oCo0a/YBNxE59x29eDui3sg+n2Q1gjQomY7XRAmMkqtdOesxd4mMB39XyBlCt9DiErvAOvFpoq
kzRviDPDTe2qsNBuu/noy30wsOiS+qBEYE619gX5l8tpMFXJF3lbivAvOgYKlCUXvsyrQpmhsRNv
a7/85RuViI2iMWHlyF59TiH9hssB+0OYVaRFUsf1UgCOPiy7upq0qx4dfB1l/181Sw4J5QZ3GWK5
Nd9Tj9rWc8OIMfBXdv3XmQQXJxEhncYwnQ7LK/pZES48M53Q0EbnrVEIF6ty5m0WqHS6NVe/aJFD
zrHsTGCNCFp/6Ks/q/zegVWv+O4nIKZmGQl+GMS/Kj6/4hNToV5jbzYWfvUVU7/zbSyeuA3sVC+7
UReSx2gIn62FB9Lec2JRypI722m988bkC725qpNWNQWGTv9k/JgmTqvlKcu53cNXl1MoJjbK4OiJ
YfocYOTpjuw3pvXQcWJs4PXQHBb6KlmdDEDLf7ltx5DC8MjJBlZsL9kBS0srPoqtB+PWIlabWrHw
0QCCWIJ9oHYtBFikxy/dcYV4gZiMx4xBS7pRnb+jUrUj0+4g9oMlRgAKaQcqgQhw8EWIAcj8uFU/
qMg9BdeLNJJRuaKhErnAsVnpMzPgUH31k2vVg6RL/+FUGJBAHZBlytvO/Wb99GCumYSud3uzN2Bl
7NM1Z8mXcU7PJWWNgKwYd7Y5zkT1OFSUhwB3GSOk54ovEJn6yTcA/9pOkQvijaI0WkR1kcx+fga7
OgcGEulL4wkvnCZGeBodEL5xfDULQvwXO0q9JfZg0Om3e/EGQPC/iHl4fmVwc9o3SQGFQKW9bpB7
mCak5owx2mboRhA2iBEBqksvtKr2TGkzwK6bDvP2wZMclbewz5vUtuN8HHRgJuYvsOtW1+q0ZXsH
K12mJJNPZ8o1jtRZMeErkrAM/x1hYf5ZwZCVZDDHLWx9bgly/jwb//OgPDIScIYjthD5s0QDIiju
9Gd5D9deQ5WyifG7IIL0fR1extqlI2ON+Dd3RYs//Ft9+ObsaZrEJDXlA2HdzgWhVxGd3Mh5FTnn
eyDSQex/9vMa7mubtwHdpIsrEqpTK8lUJbdLaeAr8c4F8D4c3ycIX+G4d6R5fMiRrbXA3kXjgUjc
nw5qMCl+EXsZB7wrn9QL9WuYIgaQSSMlws6iM+RPqeQdhBVvM6BaADQvLB73GSeIbJUm283+NvAC
o9uXH9kct0nUO37zlUDUzW3ngJuUJk6JjYHiN5I3VsKUaLMgFd8R0kS5dcQ33dY+V6Q5HxXoNklW
OBC/KxHZZdaZZ/5XQVw2Kdl1ETpBUcC2NjYbLWtLZR2HMtTi/oKvo9uRxHl2OpbkVGrhUnw9wmhi
DY3eIawtEJdtOKxMMPhe/zXj62Hr08JOOK0a+3L3Y68rutwGarJ0TrvsAcJKZvcLzL85eF68KM+0
+2GbeQvkNWggIyMDLCnQy1nSnywvS+cgK9zxUMs3thDFJBPcMrGmkxSsNv5bBtADbMsUXnMJcznv
/bUxadvSI3SIJ34tslCvWTDVr5OY4/iKYEa6w2Wen9FZszTEGuv+GH92hmHxQ7iiuHf3RJRyInc9
ymQjMQVHoCtQWjVA0nAJpzit07osXM/5jtbqdM0c13G7Ni4mg8kHLe0fDrpuEHRfvQ8zVhc4pica
bOqZzd+5Mn/dbpkQfVA2Gxutk7FuU1heoBJ84s2ouVp7QipHtaoOMzCMpFMozXtH8RjZsKvLIPRO
TbvQlKeuGgPjPHJPUHja/qT7nHdf7SneTl1tu2LxmwQZhEeDvQrtXpgbx1gpa1PFqR8ylRznmpL5
bNkCnGYlD4f3zwR85oXnW2MpyEWVN0q3FPtutL3RIW2R1JnzlZpfjSdjvyF+l+nrGuXJ26QJPP33
g/6G2DgtpVovgBa5hHFm/VNRBWJ9bbNz1nOPvdDVJwYU+7hIX1YyQd7zxHvTrV9MGBoEmMSknQVo
c+ZP6L0d65FvupV+jMG7pNXmkqCzdHVAwx88FejLvfPFUKG3TBcKIsrecHy9JYKrV2kM0JDAp8mu
HUIIJvNbtcgN91UUwd4MVudyYc96KkAQrSpeNSgv6FyOOMqppKHcYlIoKP2JTpvweX/lq7kWawny
Qci4cYZXgt4ouyAhFzD9nTuUR8juUWSMeP7u1klQCdiyZkpCRhnmg/TgIOBEl9DnJlintnCcr3N6
oM/kDmRshvEwQYHaFPK7tNib3aq/X5fn8A4jH3JCJgZo0dLkHenTIrHivOQmj4jV+zzAvGxPU9Jw
81aJGwUVE7SBockYAuUEU7opL5uK2h1RqEeHYLbaqtAseQ6ln1+KNisGJppwEQYXOIqh+NQQke0i
aGs3mxCi2jmtGyE5mgyM2ETkRZRD2BgPmd3iEv+UCh/INHG6Vzl5xUZUyknkzKixauuYRBOsSu5x
qQjAdnwRwUaLDpbRY/yQTJQXaYo53unX3vinO312mkc7FHbdn/2QIEMMT7Uxjvnnk8TPA880i4qZ
IFzcmEqHuUftOzUrtL23ef1Q9f3lgah+7Si3tPuaZ6fj8IESrXwBi9ROiglNEtQxIV38JfCO/lnC
CUYMsOmaFGkL7shhjOOrZ4lSBbRns1fxKJsl0JFtXFBJENKDZO/6hOhWuEVoTWA88T5NntcUFkAc
DhGpJQmPSpl0dNlJuYBE2Yu2t+uywAevwXSv7Itj8TprYKwsFAhnFeYwVV6q0oVh1ozopih6nnzH
sGHZHEOhuz/Eu9qmLsrYQyZy4gkYqG3cAwqrf7FyGmba1uKEU4J3+wm0vTZevX0mMYEViH116khb
9D5q7pMJ8AOoaJvbIfqineU+N25jtoPhb+Z/Y1URbRGQlIqEB5iHpzOFkkt3HVV28VftTROxTfOz
es8885aDJlZt0uxz1dFNwFGjqmjh6h5qf3ABKmh4JY1GCkpF0AN8wM9hh5Jc78n3oaYp/lvZt+Y/
saXaHrZ5SUP9OLjn30aVIzLtcGLdNUYR53gfzF4SJ42J6fIqNXyjujxNVa9KDoYtyl0PUQHjOUt4
qLewd1q8DnEbzB+g4NUgcyDXFqgZ0Ucy91+k+Ui9j2LTiOzR8e4orHuOp8BGHidQV2Hf6EJ0AgX7
iFBynZ2t149yZEW7h/Emtu5LNgEcnQx0vS3XUSLMw3NaRFw7AIpKJdDker7yxcUCSKP/uctTadtR
q5RkpRrXKLGLbb8VkpOrooxE9kToAICVFXwoprhERXAGMpaI4thdEsXUH9sxYEtw9czKyyE304mw
yFe1xnpi14+kGFHO/u+uXIssWvMO1Kp6ruzwKO7e287hSwPxhD/dlnP8oks+9rWtIuLoGbRsYSfY
jIYWSl757uNInf06WfYeI8/xD7nimSlzBmUbsX5OYpc3RnJbAO91wzV8ch2kszLE8iBjxdElX0gn
J3sD0jILvHmDVHX0z5gFgbUhzHRV02fHJ8zH4gGVC5hs22or9dsaAPqkRAkQh8frDNpl25lhm64M
1ZE6Y+1TfhMlaWEspzAam8yQNLgYcjcJjmZCXJkA21VPf9dlyGJPV2gS2u8/FA07d6uhb7qlU8nc
QoUKOI2APn4IZbchXrhqCDPlPt2UNhjR+1ng8w3+kOVkLy+jS4Aljm7snc1carz+AKSP/CYLtSXD
xI+qjaPzjVdeHRDzoWUEFIOj038p0tdeZuAWs888/Ivfxh3mrz2IgFefC4JAv/jJQRy3fLFIa44r
aO3HRfMXs2m6Rq+Cu085KO4FVsbxj7noN6Mp2hiarhAoFoyZoADUbOaophKVUE5kTDPDlo8EEgJn
VLiKyxLjX1qJ4ZmfLBNISBuxEglZyYP4XFBBKPQubIdNPj1P/KGdpvNiXWsTkaqT7nt69nKAW+KG
coURtkp618W3VWNGlnYpVWzzBLSRzG/99rLxQsRfd6PdKnXIijNOxJ5DvH++5QiY563Qqid3apJf
B5MS28MVvDPscQkd5CmPI4uWodaGVYR1mhE+hLDEda2TUGW2mnL2jga+KmkgvjqZDT9nB7QQNgAW
lvQClxXZ6dz859bn2IvnGFHN1uZeKLVA9bbxPFefGQq75+682Z4AjhvYPycaUwuiAUa4N0SR36zm
L3Ixv7ZZGmNGfhDrvvDdzgpNKZh4NPPXdHnDretyONi6qEOioo6YOwdQOYhzFq2qPJIU7q2RvZPQ
o2IkhsyeOaNUSAPFU3vu7LbtpiWrF0Widqv6SrqbCIVmU73Wn2A9h8GKDQXb8N+Ou6GX33Kvr0hi
e53zf5+UCb3dOWov4kvA4CFSmvv+pb4XmVvUGE3yom5LhKfsp5UH6J19MFfzpNRL1wCMOemM2Ii2
wYEYU1mEOd7kzVBWFqOl7Y+MjxITqnYz4pCQ2bcBRlrCRePDdu5corwXfseTV8afmq/lL4djXz2L
eWPL/U9gvN63JFUukVzBEg3rb7vEO7sskLfLNwJWeGI+fzkIFUxnypKmOSiQxBbN+rt1YX3FfNB6
REQsSADhdXcU2AcOfcR++WTVutpPaRhKARt7Z89uziNyYRMxb/vv65m1TKjMpYIBz+8C98S4Hi10
xLH2ldpZYdb66jE8JMh6bIhAsHI/zAUTva6zTkIhAbXH6gnBuaKwSWHGRKqkasde7HgKPsqNBwX3
s8XYr3FnsZuZPMWX9yBA/bDu7y71GOXUGTe/yULhS5PImIlyP6BcMpZr8DU4MqBFVs9d6rWrhPPd
XDUrvMySxYSQp800pQ6d1lDPw56Oxhx6biuL/zzbB3Te77S5XJFYwKG3S6033ccw6w+Yb+ZzO3/o
Zvd7YQK8/hXv6rv2lxsuVHfYmqMSB9BGnktKWqKYhEGej+Es2R3CME85rDL1+Z24TBxzCQmgt5xt
Gl5+fV2+7+Qxi1unVIKzdW13jSXKZ0xkq+wM6x1j2iaMz10Dvs/TxoSxvldLA08Plrcv1ciSRuP9
l2Cr/Fz3P419vv5VnHc+De66gLSy21PuNYqf8bYeMQKXFswolKyXD9mzPC04b9ihL3E947ONMsco
C5WUbRwzJUzSnQA5DNckrJ9ffxSaM9X24LOvBUdl7bGDo+46yklHVQemuuN8vygc5qjZFhIWcwTK
bG4hck5nKPcsjyYORifM0sCBiNfrroQqj8M/wGKI3e2wTbrGfgzBuIAzkK23rPO2RL6JouuOSviY
5whYIyssFSuyNJ03tHRKA+12rovil82y5h0QP7VyhqTwE6ifi8UrIG1q8KrZUWNWe7wd+kTT/WmO
xCKCl+JCv1fUbcRQsOxZGmH1DwD46NFTtiz/0yBebHOXu572/oMfYNtJGcNT+aEvsvMAc4+WQjmC
SyLjvCS80sc0vXiO08Z15aAYr9UdKDp3ycaQBUBcee9uGw/4olUZiDfVo6YmI50kLAN5OGNcbcs0
tf+15QVjVKklyea80NKaiswThnXjryRHNv8ApsxxUJssP4q8fXYaFpPm8EtBAQHDuoVasz/V4J0m
XI1pGo8csmQbhH4PrBuFhRr9h+ouLW4D3rkTM/Qyw0C7EV4vz79kWhwX4WVIgB20bPTPMQ4TMgzz
MRGJSOyLaM0pyjBM6j48XLLqJVs+LOmRHtBLksnp+yXigMUmasA2WseRLpVRqf9XOMetZhHcvMBW
CLaQW2WgslxOGgZM+UCHFA0Am/BKxAaSqDlpSnOLP01SIVH1kswn7QwBnjLI7mGdVYl556SRVI43
NkN1STaUz+QQL2F/tsRlN+FfR+KgfTAQL1g7V2r236kCjmtNf97HN2SyQ+uoyXsO8VDuBekPsCkI
7tlK3ejvRRK3Gy+EuB54bUsSfTH1eySGaXyG4GxYZlocMbsTREUKeK2ucFpJa3L7HqVO2+N2fA+N
WWH4d5HhKfOhbzcXtqSqCpzNx3VQGhD/ylGVFlBIhoaPOg05ICBHBr8t3X/J5b7ncKsmEGJU1N/g
STCLgz7pfvcxIADaR1F5CXoSvIWJUISXlGzeygrdelD3eFMjm6OjIYJnpTI3b1XA6/KfVxYtJSHA
L7piYiCgkT1QpEPJOXEdGU7toGTaqX5PGe62Iy+ETwMkBRWnihO5K3g9vNydoM5+/29fuc4wTVn+
KqqKG7O/tRLueltLMzPRX5EoGnJZXEJJRRp9vD51UgWzEPGpN5zT5czBRckExzubeEeEzIHKRsZU
KLaXY1/FxYhf37amc2yjkVTYKsxNbF+r8xC4EeD+9FQxjY7QRQt/FVP/1NDLCxIjsmVbYsTtmsOq
JqK/gi1pU7E1D4koVv36nQGbWrUq2H5ieePPmGxN8VPZl5x3f2OTXYiEkp51DvrbntVbSL4ARqrn
fgbfH8ny2diuMOxx8VwwSLX7gRLIgwAnvFq9pW4hvReG+Ce5BOhr8LCOqDnsw4l98vBds9JPgst4
YiJzsYTih4rB+O25WgMxe1T0V94S0aoDIyilKslHZKJKjMySQ8PMervyoWHnOAb6Qme4JkksTGDk
RIsv6cbKyJv1hFfvuNSM3C3e17uxAeEuvRpdWiVX6/O2BqfOkmo/UdIFIf8axh0M2F8S7fk3pQ56
w4fvpchCbWng3o011jEQNMIse3EObcSfWHYqZd0B8aWd8sYnJu2hMQurZ93ei4QDfEuBOgriKFQv
9IQMcBxhQt9dHLwlkw+wwyhEVVYeZaRHqsMM9/DWAV990t7IBUYUOHeIO/Zw05uf/kqX2ND4oAtP
noVv28h9UWAo5WyT0h2bwAMHNyZ3YISBiWpjiEvqK0Z0gx9l30fARPJO2DkAZEWaDPbfG6byxZ6i
Ypy1yxrqD6GAL1VZvwYLwj1ZY9SsoO6Tkc9QJ5QGwaTyqXoetFV+AMbCRUSojwdG6B86vzbF9OMF
svyOHQpyn34mSayJHm7cKrHpvcA7hSQpR41Bm70KoDI3Vgk3iORfYKreeJEmpWl+60iEd52nkHcc
T8HzfsCM7jTdMdM5HIQPhBjUTiDq5RDfi+pqSWkxTSdP6GQ4P0H/vdQDBg56VBTHc7PLI6eI17k2
CQCK1vlN2m9bx96xZ575oatindZjy+kuCtrdzYDwLG2IVZO63BQ1b/vYY5bVNFKnffkGVNMdom3v
eAcqG3ezHVoC1LxsZ6RdD0k82hBXpDx+XP+/UtcS3dkmo5dH1dhQi3XrHI6tX5bWj5MHDc2fC1as
r05ZwODlwhCwGLh352kZQLx/D8/zfGzjXKJwZZ441bmnp4pKSizcmne6Q65lEYgi487D6wEiQiiB
oPDPlGAXoOaRYknryZq2icezT/IkYbINE0jMneZxa/YhD20+SakOkoLABPpKFyJivoo+9QovGjM9
pBRZezMEJnnYueTGgy1XFMQ+RrAB7Kmbmep8gjQqycTw1wgOo7Ba396o5mpMgaMlCpfh6N7+3AD3
3VhOQG7LpaKNe2vcOPkLabcRuVLOd7xcaudI09SQ4W/w9RnDg+5uQ/RL287qLeO+yeMdEJuoh3Ez
Ubkn54J6A+Vjc7ZNpA1r8l6P9PldKNfuURftz3AUPA51Rsv9mPid9sRolpxjzhx8fmCxGdgcsrW6
znSpQgZsy6bMAaZLs61BujkBmHS2HO7gOEQFtkP7V2geabxBcK/SWj3x0mbfvAC7id9c3wYvaYv/
egqy6ZLOafuAnCVP7a4IjPbn6nKGuIEIa96wVO7oqkHARoE0cerMVRPVWcOkPOWxjdBs9DLlNrrk
MxtoGn0JMTYN19tJnie6cyHLxgW+5YSWZPT1fqCBkzdgJL4FuCP/x1SRtYAcyx83XTr1tNXtde4g
tIWrmsnD0Xp8S57htZj5qIgPSQ0OpKPe4IYpTWaLmGtxf8ROGsipBAY/UCFBhmuXrQs9LqbA5nCa
/tGQdU3LOQrBHAUkvGvwc0gN8cRIiRVbp5NYmXrYeBq0Vw/oisYY5FrH3yahRePLFIJMnyD23nZa
+yDq7mFy2hVst1aBHQH2wSPFJiIBOCHzPR/et1P5cAd0AVZae34e1nGT1Dd8iVUO67CzM8kLU3jP
5bP0ug3zIeaAVZu5Yd0Rmjgvdnx1F0tUmXVGOozXohjiqgytfh7ZdAlzGYqM6nNOIatb93S4O/dx
Ce/CKdHoSjIeaedOySiyt76ACVeHaa2ElpumhfBuiEX7D2IB2h9cnVy/AMaJI129DtjupV/nk8Vo
fQeU77j17dAJM86Y4SqsiQPOfHBIgriogWS15uWwXgnT7cO/XlwPEZFWpYTQQjaUUhXF3Oap4ayC
x/NbWPA528060SH+v71yid2hRohlNmFtrSXQVOKOwGvkGhiPEEK+vnIUSlICIIgUqcLR41keqcwr
/Hc4Pju9PZankUemtdA4IxqOyHy8n7duqJ5/Sa3+JOfkVBQfBSblRMY7ayc1wCoWewdQcfhru+/K
eFICr8805OawxSxF/tyOdClWzRGKpg+ci6E9yLKHiV7AjYI+AO2B0niOkuy5H9zvNje0aBZ/WMc4
6D3aTWhJO/+P3ddY1hrVzm9Q/dRdzxsbFKkh/sJzIYWffGI8aDAxDkyNpggs8sbbrguXFpm+Y0GY
hZR5sKv+jsAYUEvDe/GTHNtbFjlMB4XMBqwiA1VElHROVkQX1oFsf9J+MrOwmI7MruJTGzv1S1lo
e7DszjImT5wKGoV+k1j6e4Vz5X6OoT8pPVWfdXQgsGV3deDllobZUy9utKhnCJpp/RUz43YHQYfx
GLNUrvommfuSEafwFOTeL4O2M/+5qhSsb3ZQ60kS0BPwxvPiaioAX/t9AVU5vWOaUBfKz2AHvLxp
02d/VnH6xUdTpsD83Fv3uUx2PFZ41p3As55vqesId738QaDbFHkkOQA/UjM+tPd0ZYdtG9VoDR11
WtsYZg4zU97C/pffYqbzh4C4Qf3rhS7c8d5s844xGdE+0KTW/kheBksb1HU8wEgIT7YIOIMNkbiO
phZwRMSGGNigeIJ6iQs3RiJRMzmldjhRB1eM+0s8YjtctLWNKsR1QbG5KL83ukEqtospYRXuhbhU
/TiYNVWhuCNZjfA7ZY5JmLCZm26S3yikqM1JUe+9u48Bbl6mmcH2IyAZfqHjDBL1MoAFPHNffMb2
c5S/Ge1xtCiVreC4JZiklIJaQNnQelyDJYwkz+LNH0aqRDCMIzkOijQEG6HrOb1l2G/2c28yxRsp
B7dp15bqw+CZVA9VmB4v0dYmRQQtj/k+6iS7MiNGj8HT7+i9HJpCMWYtiQ4wrtWgkj3aHwHBbhoX
ha/T6jiBNYzszF74PB6ek0RQg7LTmNXH0wrJS9yhGWAAIqv8c9CgUZPt7Vy7jhp19yMUWZbSEHCr
RgSyZj8kjl4DDA0+3+jyWu/CcfQiGvhpU4zshyNMTWRGPG6g+DschYC4n8WJWdhlHF+RNw3T+Xyv
Q1mWODeNci0GYwggbysESz/sMGR3RvqUwhQay1ZLURXqu1VxKHy/qIGXJW3GicHTg0iSvbgEYOZE
qM0dU6DImn5i2IIo59xqU/vf0/NsuygZnj8pGyjvQ9ZIAvkDOlHX8P7Sm/fkye98DePogugGgEOV
zpsFQ7XHKAoW5J/5G1xR+Jpcd/H7Cs52rGht9X3DgM0C/C+bsX/2fW2vl/rT23cJmTcnwVYPBVT1
YmWp10QoMxV6VEyHLxhUV0TV7Z4191u6FhjZKZ+yrxHmBpJNNZO9TEOoiQvR5H7H4PNt5hpq+gFJ
uwHuFGpTqodtCBa7NKu2PrY1OEm6VUYAJ1b0FkXK8RZraeJYhLj/emmHJQiLyhefe3cIVEXhRhgm
HY69FMC8k/Y/vkHV4jZ4f4AVFR+bGIMlRz4LB8OKpQzDCGBvviHS06JkZH5vvk4JkfG8CaU7luTB
Qq0JY1FoHaIwYTWD3ATfqOz2yYz/4K1m1hAp8amd9YB8WjxBKrMLlu6HHn+ARI/Ybb+XWrqHaHQf
xaN5acpzibHYup0fTMf+dGkzenWoY9tMXQMdfttegx4keI2MQpwMhrYOJqE/pvgABeM6v4XRSEry
Pg0b+Z/u+lXH+fTRC4zvcVKN7KksZHhU626or6y5EMzCy26wfwTemP8Y9W3zHwN/JE7rJvNIwVit
2ngOFaARSpJFMhvpuYiqI3pVDpJYZp2m/ab5tjZPMr4S6u54KXBfzwbeMjmlCy59csrS0jJDnFTt
9Hhy6NGL6XpbJcEJ4ZRelESQaJL8E17sFWszv3kVUtjorsac7vs7fa8ihDBBI6dswAFNzwZcCQyS
uMbzaqSQ1rkvP5/zWmKlg/1c6M9Z/NXUJKm0E1oidCKlnd0Il5DNaQokq5kI/e/PxylB1JO3e7bL
9WjXWA3Q4xyFWZ97PfGT+JowWAk/q8zWL+gK0qG/yaLG24+hFZt22ifj68wdHYLzyVQwVxl/PTz7
eDFBi/X93puoc7BBvsk6XM+yCd+764vjlEu09fuZGlkhu1GAa+N6FtWZTNj7S//2sK2Qsp9HH8LS
1B7v/G0IDTuXjdhUUrhgKXf/ddLdTp4fcq3AQ8HEYAfyqRCRZTPAteJB7h2nCBRElbLxE8em6QKN
xs2BU/NpxOyc8+ew+AV6avEBoxknLi+y8NOmDxgX1DGzDgXDHVAfdOxT2X/NxPdbsYgjzZ2101mz
ZX2bW4p+t9qWUHtyh8o4516VN102Z2PTQ5tZObiie5tWeV7ezcWwoT7tVcR4irdr6TPSFQnpgo46
U5nl5W82e0JZvPbJJZyjHqmxXLZkuWvlPwUhfv+inZUi/j8c4P57nPEIpO9ziALwQqj8Thl7XSu+
RW/eLdgTzZNowRw/Y9h6xkS0c96E9jjLsbuuvvgVumIF+Yh+1Yi59k4NJ1+wUmXe+flOvbL8UJCs
/B6lo4GAJ4mJlqwxEmZkgqW9kWNGYLdQwaQ6Sxtus47vrsl2aj4WAktTV3wnlToPAj8qiaFR0WoM
tw5iA7LZmjLM/4yOCGSAJvPvj+g0p+624icRAk8uwjrz21GgKeWgg/FD0WUv/f0QIs/Ady+L+Jg5
7qCMmvDH2wtCTbQ4PuGQwz4mP3WSi8QnTvfrbNQS7nq7/QiDuollLdg6s3h6ood0zr6606PtEhpr
2kQ2FhU3qZ04abYJutDHEMcL2Mtvk7XmLmYImgdXBKs+eF2V/5l+IFd23FcriAbKLntdexbrQOAL
tSMJ6VpqwM55j71TG3kIKlYv3Ff4iA3nLrKMpjTf8fXppgiA20yoUAbaKS1IKoS36uEJghc17TzX
EC6t96uJKWZINollIftN0gphgQK75+Jds7C6ym1GQe1x/utm2M6RMLIBl71QLq23iv2Kw60qRhbD
mW6EReg3Lo43JF5k8GkicNZ3QUIQyCtS9FllbUb2zaYMecZXe3ZdzWv7nhGSTMoHnimztciIizS5
1YhJ1JhhOPZQ+wa4kW6cB7IroPtaRsFMKI23UmQaqKFnt8wx1kgnGKwt9hFPL5XZnTRK+xOtTDAB
Nxch+Y7FRmFWn58laUPJ3QZkKGGDAYqqpD2JTrA5+KLeyn9TF28Nff2W2eZwFPKHgzhBexrcRnrN
TzgDjg0u4sNdNdf26dBPXa4TPjywALHxApowV1Wc9ISnNtmtDsrXMYZXWe5zLMPZwZg+fBkbAZJn
kfXxG+hI+pYlgYsvdde20iaTFPHsCjFkfIpflmg1mC6Gu5Cc2F9z3wGbIVXU888V2dGhr+OYN+Jw
1PEnwsazULWLaI3oVJn28FhBWKwHAZM/hIUi+0e+t01U6ZnodgPqFlyuW6Dg2GZreq3vxzaGlI8l
cBjNwmdcomF3Keask6TRgOu8c7A/67xdx6mabxB1YtU7DUtXmnDvS3vxizQYW90O+ORqwO37VlU3
96lkgHsdeNfa3+58GwDWR67XMhApPM0idhezhXNIgUPyuNRbMOnlL1XbMcwoz6tHC3K7OXldd9Kj
WKZ3mFCgP+bbU6jQFacbe5ArPpduehG/x+O4m5O4rm2UVS7cg/I5yQEmtxorZBv2O4kb0qaLrg0i
/qF+c8nGLgMnNzuNKUXWEP4NU8zPasXRgE9n80nvZs3Emhzoj+GueEJhlMWvWFBGrKbWCFJ4IEXd
MnCKoCBxpXFiAiqHTjBwKkk52+4IoXdScsJiZqr02Cbpr1loH0/NYVNEe0bc/GZCbrUrgTxPmT8E
rmDFeQVKIyubwHRjs2e4cOy3e5bzg/BpF3qHMXIO5hpE97AWOz6qNjWf0W6IJDPvZk8tPOmh3r8V
ZOXZPMeakUta0UcYiEvmnOUicmSA8BKOakTrPUJOoS6ZG0eDlq4w8z6p+VBHW25Q6+lTaq9LkUiy
vILnNpHm5MFKd6r3GCw/3RMZnus73QiYhP3PznNjhI+4cfnRXsaZ8Tn3Nyn9FQAkAPvXjEPQfEED
Pn3w9AzBYMZa5+WWvcvotBD4EimZ31NH6hi+di+2kafgWDcsv0iO7nlo+Wv/zOrJunAxRPVtTSBE
3q3qObVQMUncclymWKKw+B1aWqMcovo2kMLoKVJHhxRv9+OQE4QHkm1NOWSvJnMSSWUSRASsbjuM
rZQtvRK/70hclkhjbp78EjcnlrSWo8skwmSF1FK7Sz52sNPjlslbfqzXVLxFWHCGrl7BdPWmwTNa
jSyuJcq083mghRQwEklEtlfbJ1xZdoq4Vtd/PnG3sKqjdXpcwcvm7938YHu647NSyIpL0dtN7zNb
2o1iQicteUshQLwQ/eL8zHuno6JO78qdyp3ea4RzDIOUdc2iK7lcUMYkC0s/zhEh/dgkdTaDQW89
Neh38juUJd62myWPJUwyUbXcERKgO4qywb4aMv5ttyskcWvGYheksxkbTNSD6Czb+VJnDafITIb1
EC5WX2mV4z5X8b+U0BjgULceIQ/JUHM2KRtZkpKWa6p9wtTGjrjXXMQ+9Nb6eu9tOMd0EjTOfu1U
ap+Gjr8vCMUERgVC2GE8GFx92pz0rMNDRumGN+JdPl6eQGuZWAxAVvDObb+TQlok3LMcyWz7V9So
ZLtYMlkA6FzqPrWytXTGLCBxrsx5JEf4U9hbPlDaEbpvnau12iGNA8uWyPzodWFD0ha9ApMHMKrC
jHm+diL9IP+kqQqy/5MO6YsAE0ELQI8e1NnAeU7+GygQe7L/YOG+l1GxIzGwnTLK2dXNFHPg3omm
v++hZJq6eEibBRJQs4t9U6BmSvkCbWppswqXK8i6OqUVWYeqLi2IAWSLUTtTQx0AEWEtx6wn4Cj8
oShxuTIbEqRjqu/klKnfHEn/dC/c8vxaFr4gO/kaeO7At8lntMz8Av8hQ3UlBd5VMYxNM7X+uFLb
fyK8J4DoCm6Wawm04RzZ8M4xHuWhv4aMSYU3OcJrRUrg6T3+Q/tWvhF8G2E1446Nwh672c4leJa+
RPu1oW2MwGwyvABzVCgQD5CxsFtVaPKa2NzPDYB+pzooHz9WJIIVGbh0iX66CcE8K8CoPX2FnjFx
MJKbgOL9Dh7Wkn41W9GPBJRDAV7h4tABxn2U/myjFKOBkZ4F2KTdTqGMA4CSb8OUu3nL/1e6jCD/
MyEb4+Vmx8+zoerEKaaz/volD/b8s8V4wSuYZwhEYBL5oStJqkJz8E4xWVIXVg5AZBalOvlsLtY9
tg2m+Kkl4HygKLCLCauKA1LfbDLPcEsVGY/nBOSPRDjd08Gr+cykKkovqwmjJ/xNUguyOiKLoiwu
8vSzwn7tjRkKotVDNnYyWyUK98AcWpQG01zGFedW7qn9EKyYrTn5vMmMl/JgnbHOXXRwxHAkhqmy
fztAYt4tI3ZvoCJ7HM3DXlBn6QH4yejaWRWa+kayakdDFoD/4EPvS/zjVE2cR/kKoKRrtwRbJZwK
PloWFUH8Mx08LC5vZ5hpj6J0Q35cReBSwYFpIhTw5G3uPWtQ4F8iziRmUdp/5S9pCdEUvzjqeDnB
Y3TtzzO1zbepldT06m4DouRWr9wW4tp2G256FjaDk/SmLEXwQMXbIt2BNO05Lgij1ggsKwK395AP
UFe5jF26da4yqxCIq3zUNxY0bI9uRzTS2/c/9wGSsndU0PE7j/ILIVLJxUxCKTciRdbZnOlaOVmR
3I/BkMeXffY7/Pfm0oLXGU7wqSxd62W2mLKfV0JcoqzliqiAta/qr6Od+HXSkVkouT2TvApEd1uF
MdCFpQra1AyzFg2/KK9N5+HIFkt0ia31ZrH9ZKxVbHCiKzZnkgde372wj3ziAw7qps2spRlDMEh3
6722618F+X35FL7U9DPaSHC1kwmmShq/pJLcR2mc6/nPxNGaXncgywP/EmeK4CmlhPxDi6AB5lPC
y2ZnCV/HMkg3MLDRwTXvRdZYdjUIRgUAx1DnnbU6MkJBsVAW6gnb8bh7dcEbl3WTGdTpVtBDzQXX
uF+/HdE1ZXtxXcSy/vd6kIkRDDrWe4pXFRVzH0GN0CLem26iP+9EsIPupT2hWJeAHrS++as6/Z8m
zD5PT8VTp3Y476eYeu+Ay4B2RD9t+h7xH2UjZ/EdJAUMTcCvR6YQt7F+XUNIQ31xhGiyuwNTUMaZ
KCmpbaYuPz0pstbJ+Zr7IPcisf1YnmABDKwBWs+KmZdT/YFh1RctDdA1xR2yrApyd94PoRtyoLlG
/TNJQdODARDRmpM9FcRI8WCwBoRSnP93khrvr1z5rH++4fCi/d2eUQ6IPUyNiGAXFDaxYqNZftvQ
tqXZf6JL2AjLGKkyg0hWiozH7tQvi7j6BfjRBZS9PyCvhYej+IHrwQqtB/ebrAeM+4pyxIXF9z6V
FD8T6UyNer3RrAPYRHx4LkxXzOekfX/mwdMFM5bjYaV80XS8kNS/02F8cJCr7jP9z0pWtGySLOUO
Or/YDU8nxrwAfy3clRKgusGWxCF+M3NrKct+lmtPrZ+81RPLI2EcE4Bm+C+ZYdf1FUM/lEKky4cQ
sYElHfUywjNFxXmSBLEMbc7HFhSYKioxL2P1/aADjPJuTq4cJyBEmVjPduSaTFu+6ctnDE2SOZlg
i9EMBumPIwHDaRDc39w3zQx23kJM7J8+aP/zqD7cyisfhmb8p5mp1h7Z7fW4hXs0/SJMBpF0tFvU
rGrrgzIqAo1BBnAPreh86Jsb5gQsugsKq6cnJbnsKvKPTIEeK+GnN0v6PyNGTsv6pPTwv/j1l10U
hk3z9XloS1wuY0CAZz0kzhVVvaKhltf8HACavWF6hGkmhos6zHNzLEQZCoEjw1X9qzneIHe/PbnL
yUwrIMIl/cY7gd4Vd8GU12/2FhA1yF9U1L1yuEwLMqwe2MWLrLCgrZAVFApQHv17lITz/wG4h5Ye
96AV+Dnny0owIdWAjO2VcFaU856nFuHQYKwYaP3KjtJYHs3+3ju1ttSnklP9c4cKmkFBGcZRA/rj
/vuz2AEjJFdLxP2Qtt5FukBBz7ySBEW21L6BkXoxRhPUcGLk644x+Wmq9E9/OFTBz0CD/D9vxYNw
LD2nOpt8QW2nXi/kmNT820G6PXny8F82J2g7a/M01JANyrflD05ejjZ4c77An1qIG4KbZ7PU9fEn
70RpzsFD+wdcJYjFLlmDpw9LzHAYFBOWaewwGF9G0Zf1hIe8AZq07tBBYUehn85JRgdfuOsJcjP/
4wjLc1XOC0Xqm55CQ/LEK7mzzYDROzjkoYJQqcFnIQ6J3znd/V56X7uiThFg5VsLVu5rP5hKH5Bk
57LfAQMzfeEQggnOfwxwGmrKvuph0/B8YebGw4p//GuiTvallCUyTAGk4X6Mg2rOvAmjJILmgPS1
8ERa0xVN/iqCMs6UrfDgRLpqrCiWtaDbf1pVexwp6ULbBEfDsszVcfh/e3BN5Sx9/emkIin0Xwn/
J8nal8eShiWEgnXvs04C6WUH/cCPKWr7lOKqw3moQpgalh3vPtUU5IGfcb18yhSZq8Ifdx3LtNQK
WcXDRq4HeuLbrYB3SM5eXXC3WnnxBOyXiSwdAYDFwXc8YVg7Swt15+kivruTmVVwF324aBnNhbgz
mq+KCU/wrlP/wotNa8WKyI/IoUCP8mfMsEEFktaGxsOpIp+CjLb415yUWLh2BveHcnRWaILksKoX
Qxw0hJD+4knPkLXXcGntVKvVrMQhDIMOWN/qXn8QrIoBbkmuMfMpVmLg4aGsanQv8ZUCG1nomPU/
saUEGoGLpmhtMOq0nqp3u3xGG1SIPchMo9azmJdVBo6+TYhZo2DJ+9eTAdOj2dD29HNjvSFhZ1R6
xc17B5M4b4/eFXLjEgLH99/XwV2KDoFZHv/8DIAS0WI+Slwox7+XC2H/rEXz6eiCWhxCjB4mqO4N
vMRF5vE6Nmd/MDLyYxmnt0bkmY6YJTNTHbmNyz6q4Y3Bg18C2U+HO7cRuMRb0Z79DzUxO3/htSN4
wcO61zgWm3hh8smS29aOssVrwaXMeXnRgY7WuKCUjPpDa1qUXRgMxL+XmcR/NR/UaPwdx8NB+bxw
ctvOkytyZaZF6lHgTwOl6H5c6vLoj9T1818zGjuxsP1v4fTsZmAEOW5DRutdW2YAZyHO+HsBLbMp
lLl+yE1R0Yn8jlXWR+pIy8r5VEAyon5lIFu5Z7pKP6JKevFb0vvpH97AlfBt1yGqbK5uNlMflJYW
p2e7czNqPVhRpaOBt54bzgAlHL5d3RHXjtiOm9dE4HEAfEsTonb4wM7cKa/LWoV6j06KNoF1maq3
vZxPC3cD8eCDl6n4sHP0p3NCWHMnKZ68HoePcTYckggGG+WK9jwqCsiTD2ds+lod0vvoLbYJC+3v
OH3wjksxlhgl4tY7sKStzk6A7XXAvT/oWeUeIISDHReOEYW2Zx8WMPtYFG+5Oq1zGZzeo0bGSsg/
NYyplPO9gCodCKQQvq02xEcB6JVbsq9v96GRDAjvDh0qRTz5gG01ZnphSQL9Yuvn0dWGIZmvQIAh
/tNnxhiEC4w1CCIMeHqe5BMFQOiKEmNfs1F4bAXorevMi2dmOFM2Pq+edbokadib+WzQg/CSsBpB
1mU8uG702/TWMWCyEY3fzwQOZd5DsBuCyaJiNglfGMZtGBZfjK2DZTMtAByGphwOEdMhJrpZ5vY8
WpstL7aHAUJRsC/2aLdxtRN+J3oANWO0cOgzigPm30hv7IZXAwUlE57X9ofoXQGJvNC0edasbInO
N417VBWaWOXJBNouyVB4xkRsYb+tgTmYWfOKX61hxbM70AK9ynMDtCv6p+VU+uGGPEiO+aauhrHV
hiSjgPxq7KQSHu9Wa6ZX6RX23fH4g87maDaRTawBmBEEbthHjiuN956FxmhTBgUcAKOmBBqquSOx
8VA/wG/knrQFUUpeZMINelvnB5w6xuFfoDKLXtwwF90yNmXNLsTudONwxu272UiD4oFtRv/bG+H7
NsFWyID6joeNZUO5ikVNfdz0UQHI+GJ9/miQaPa4Sipwdm/pqz+T1h6/vIsFb6hNMnAZRKS2iMOW
uoMF8ZjBu/XnDKQ5c8+AhcUY7QVdhMHAPw1UuMisd92dwhXqdy3UT06llGyqaeBxbmuGOzADnnEa
fpyRAzBpCkAtCizFk/m3rQUet5xQYRsYmZrYvsYOBxXT1WqWcr6ukO26vEw1REqDdra+3UFN1EZt
t758t1v6l92YCJ+7UQWgbjS/8fdSWhUcPasz36ByeHiXU6nr/QblmAw5Ii9Ci2W+3JtmO1SXm0jo
OHwFgQkWaERa3FH1orE3NfHQQO9U4Qs/b1gmxSz48cNYAY2vFgTGcU/2bnr0uunwr8jiv2WtEDQJ
tCfPnpY5xqv77zIEv6u74sAwH/NvgO0A7b/MKi6NdBjHVbUlLayWrM5fI90CtXvx3yF9fyak9Zxl
kXC5tl74lDbJ5xX28/7HQOGjjs7mWevx3uOSlIZx879wA2sQy08xJxIN1/C9hhDZiF6zxxLbR9Pp
REmUZSXfL8TLOfffWu+1Fi0eocfjsZiIC2k90nvwFYktF/vCVmq16acyclihVSKCSWA2BZJvNIX+
yuCNBt1h57NhZhE9EkSBra66pgtXqwCN+9Dh6FFJxq/ZlViObBIZDHUtYaHcKWROEAt+tzVnvPgF
XJgB3LlPbgn63kC2er6pLraX4hYWw/230Bd347/wncqszjoq6Oa7ZFesaJoHF9PEShbgoDSGnFV/
c2NFgy9WuxmMsXEiGih5MlaCoqNKjR1NdYp8lRt0pqBRacW6xyQRIr7Hz8g/w8eD504O79Ua8TiS
7jA+1vcbgyEqyTgAXCLnOjKE0hM12BvSjUV/+v90tgzbX9830XuDBk7zRKzfr1y4ZK7EoRYWhE4f
x8JMqe0Po2ETSQPtb7lGblETp/AVZiAWK6+YzEDHAdRLVy5EmNYiLBMfHjTam5BUK2xJCGEwA90i
HqSYhReaiGnvBQfFeUGXN+ntvZ7/Kqd/d2SJFScBViI40i7ihjlCrjRrOCbQID5aBgylebATlWiY
8JPI4gJ6CyYs7XWkUqaB8fa/flxJoWpeg24iW3YfUuZDT7qDa7v+6vTdYM5ziZ79b3HfLMfjJXFQ
iX44rF1NZfaN/FVmusvwey9wiub/qk0a8nU8J2PtUDbZXeWxNHhVWb7fDJWeakpuvJiu3LT9vlsU
LTMwZVX+SAp3gGcVWcT/93cd4v8zf0YsQybrZEbL9AcIiVZoKoSf8wsc0gpnRDewb4JBGZ78z09p
RhfQ7MsvumM++p67tUi5JMiBUWQYlOTNl2phJsBfmV9Tu+Y3qsJ/+DX7qeC8wanQWyY2m+jauW0s
Xr7MJjfneOhi6KI7YBLv22ga3G7kBSQT8VqwxK53KOWDkiZcuCeuhCVn6EVPszn+od9qz9Xp/d9t
dMMqzv+tzCrDCxSHtp/nE7noSzzehd2EzQDuWRC19r58nvlOPK8TRCKbqNmY9w11njgz+CZKuY+M
hUTjJO9n38pbugQDQLfCI9VxmOCT7jtkGMiI8WeHvr66ICWP5HMXyI3u3S/pH3uKdnZpG9CPvgV6
f4k6iO32y7vGdMXIUilFA38EhODoBjuMsm3anzk740FGqN0hqsiU5NwpuCMom3t/FTPPXCx+nCCK
84SIQOuMpyLi/zY9KY/wBpT4NePHa/eVit5Rx+n2+SlrFhgWV4P8DH9cCso6Jn4QbgGVMro8cpa7
ntY3SObvGICB3rheQsfzdj7CJ5OZl9a0PvW6uENYzS7JCptHdiw9+lifqZsVcjXSaH2v8uOWG7qy
mofeKeSwoW/3sOLXztk6wgqtheJ64U5ocTV0tpurmSHusjmeDyng9aFG2nFyzIfTrC6fwlb0lLr/
SNe986M4BzpiQ2qQAkCnZRNefIxAY+F5g9DJUXV6vUs55z8kmwBLXXrs9ZozXhi207pioVR2IqWk
lykgdYTrWE0Gap4WkgT/Q8iFB/S08Nn9CF9S5FUtKE4xFKJCUEV5ZmF2Eoy4wO99ScaJUkE4rbRN
AKpXqwKhipdYSFuHNO98P/d85U696s9xt7MTjOm1KoceVJ2wA+rs8tdAepokKF4pvEXISzBPjVbe
mgPiLylZ2t7RGfdEcKHFO7cimgI98/MaeZWissse0QQir0F0eop7dwtu76cqCasLxcr7JR/+RqZl
Y4Msjboqy3P84n1XATed4acfd601wF616WsH5e44IwgnsS6HIJ4lAFULJPMljSHdXW7cJI3vF0S7
5hdtb08ZUZJRantqD7o0QIAxOvnFGdNVtUNdM9M69JmFrM0pul0A4NIhKjAV8WX3xgNqOhLVrVV7
Pa3WM6cz4PAJ9JAdExH9wtlev6qv05NXFOvTf9QFzSdaa5or0vSqxmTOIWaeLPfF352VSHWqK4vb
o/aGG+Frspq9ajn3vM1HhzmV5vpzFRDoCAgaF1dkB5pRN/VK1Gu8eNrJ99lgVkCKbLo8/YdOUgCg
ltnhH1zbnwkED00v4Zflw9EpvkIeLaBPtsSUbM0nilZc/sHTvuwGVGNvea4AkszvPv9wSH6MXzCQ
tFNsEBtevVlFXV7JrWE+IIw8Oyy0o+Fx+Xkf9GuazRFFDf1Yywkvkqb/kr/w1R4SpUU75Rcmh5Oa
VL+txjOlkm1x+JplnayPf/62ndPD2+GzqAMYTMY5Auq3k0njdP4g9UQ+nxhnTQDinHLeEWtNQiH5
xyY4saMUnLuJTCWuv1k6VWywuUtT6UsGTVM/okwEN8pmERiTywzfVCJxfIdJ7FXWWXzSeLXHM67i
Goxvi70x7acOe9E4nIPBlSsf55c8jM4/cnoiz3jOq04flxWc/ic4BtCIxR0BROOl1e6Vw1RkELkc
YKDikJlVHbSojgPrxg5kZet5AFdySMp3e7PruVAEZF2aQqoSQwG/JiGwiR+7HDVQHBwpqo4CjsEC
CHmnhdpfFWpax7ICSnxHdWjpJppPTR+io/f2+qRBRKp2Dvdf+gWmhHsnfyFIXLGd2f76AUUT66vp
+99EPaWjaMGmxBLoYxpvq7fv6vULxbVLMy1W4PC7aKw6I54do7zu/K6/xF3cp7cct9+H4z3KfKBR
qPGs9zLl4HaQZxyOG8g2xeBcFsuU0SnoUaMj0JEQtuX8BGR/HuEBlsYyIisxfV8K6YbfCNMtn9yj
8ULCYouScPcQvpFJpWeH9040GUmS35gtclZ+za9umtf5hxRzlPU3AvY6J35CCzUv3am1F1lsgyiq
+2zMK9NkGxJuPTpFRPyDUNTDzz9891NayF1HOJOPKlg3dqEkReInnoOSb8foiL72XmEE85lfctme
NPWCTKWQ8KfnG4qR1+kGhz/Xce0IVX+Um4JWVBfn9po2hdpLluIakqf8C19ndFUHnkzuK5MxOTwN
nZNGnD5qS6IsbOYq7Q3UF0gKpkimlTDd+nl7pPdNE3Fv0fPnVVkEKs2CujyKEyR0oDvzzqmZlk9K
voZQ64MPiMfAK14nunaeHaQrZ837/8iPFJn6rapD1a7ZMXQDkKKCBQAg0qyGvQMcEDuqy50K0CQE
W4Fg4EWOfV/G9oMgaNpS5sbgfAHh3ujeoWHl78Qa2sxx8Wf3fPhh8eWQzakXDDoIFXmWbolSSTm8
bLRrUNTB+svOCK1mDnCvdlnXSpU1s4Sfys0q8DwhjW5RGeBjVW7bmVv0SEOjoMGw2pr7bRNsPA3a
9uhTusG2jYtaS3ZrCkxbvKb/9BSkhjlHhKYzYvTKKEThY2pW5NYFCmTsj6jB0ESbYidmyeeMJWmC
FogVJBmRlTvLC/R9sRuxlrzwVjqE9irHFO2a/xblp5R1tsh6gZlZ2XKHluxWPDMp9SO9PCDz6VSU
3VxwyrwZS6ObjKbYTrfQhKy+kSlKp/JP7HqDVBd6a00IJVFQ2waUpYD11gRPkF7iI1ATKNcg6YDb
RnPEfCDm6e8xbIs693RmIU2DcHro5e9NYfZxiqbDbNaSY4TF790aqVI+eXeMvqxMDIyqvrptxymp
YQbU6jxmGBmfPzf5D4gXKZHaSN1ngjfxsdjy4gTqLu8erpgTyLhaxJFX+4Wocy0BByoon0AkrDaP
zUtaYu8f85zE+PrHdzX4Bbvn98bm4o0G92Ew3DYdvYu3Zm0l5R+E2ojCwRzExG8RPNPb9/tenyF6
1etlY9IsiXd+Sy3gICFpBbxoZYtXnAXFtelKpBk0d+liEAY5XyeNOwaHEYdxJLwySfvjhoNDleio
aLeS2fOXXfspERM6Y5OBLRwRg2LKlqyY/tddZnaSfUUh/N3/vk/Ec6fiE3n353lxvf0kGmERwfkb
hShkbiMbTMTzq3zVizpmcVDtCX0FOnb+c/WwdhSWQe3OLfxa8jv53PVghkdWUyViLEyi2wKZm1Th
13H/lQV68aYgwYbM2dQZRXNcu9xvvERV4DH2MFo17USi8XC/rI+QaTkVkb+DBfkR3Fnb7PAmEHX0
asVAXebpUfGA3+/M+Xik7E41P7sstbLLmTWNhLIlRDQdwlTmw11ApDtpsr3Rp/T/Ev/3dbF9twkW
QRTkZH+xOxWhjso0fOlqnEWgQZn/VIWFMplIkBub5QeYQ2ZKs3JmetUmK6GSd30ygOYrynBEXq3k
0hYcFVnyzQrPC8o4Gl10PMARMV3BhActWWTkpZnpMS2RPMOymNhhBErJ/LcSHx8s8cYzqkmEohJD
+dXQ3z5ywJNYiNWbbVwy1nUJe8Ov/sYDyYQE1GX3uHfByIhUQjLg+bOisZsCnZHVNpAxluw/aHR0
26WwtcD+kA5URksZVyw3+70ytsMwu7vlOk3VRsGYOULBT9UJ7BWGJLaQvh7HjHyauwOoWczAiTkU
VRY4rOeYGMYqq/VS15jad82hEZbRSh/kN+2pwMrxm6a5Aw2VSGgG+MKtDZL3aYxaMkg9zwH+P30R
fwDbXgZNCVmwf8oWOma4NJnrWEV9BUM4ViY+d7Hj1pa2Ode1kCviJ7kznGw8A/oUfznD/d0j38vf
xl2r8y0QFgZHaEeSQLC9uSzC8Bkc8IgG6OLbvCr8wWTaheyK6lvcsOscgRb4NlXjQYF8qp+dmO0x
UnUwVDxokoVH/ErcoU9qquD+c/eyVhhBe2OlkLkJJ0MF1QaIYNmMbe9dbGPEmH0rWIPOMX57m+Ib
+3AFQ2RUUteQtJeNw1higbO40OiOjxQodi0lUWpcKZVOa26y9t0alyphuu55T6QQbtWokPtLM0Eo
UVjGMtrN6aPe1LqoVYq66mxbZ4GECmuK1zXacITJoiXw9ptaTV3VNv5cPXBTOZctcYo7toR/juW+
SgY2cVZ0B664iBxb8zhXlSjLfzxyv6wPNPXLjsmHEREKIDP6vx9F9L1JFx9BkeLhy43UEFWscYwk
5pDUnMjJIQ0LDPO2QHKEFhKwdnBdBimKRACFcR6INEXNmvBjN3p9IbyMs1GJgfwZJs1CWJIZlKuu
qwX0xnvlOUO4hhg1rWLtfyo3Nyscr5a9sIxuOKcC8l11s38NDsjIBGKFRXTvFwGimIUGo/8g97TQ
trRW0grPbHamgbreCym3E6opoYGn6AVxq8AVedAcG12n6fxox4xIADHaAdekuzWxiTQnbeDTzb2m
5RTqGrkj/Aw5YHva86KG6Xu9TzR4h1F1Bkq49F3u3czUl0sJ4Lhm28QjktJnDvtvvSFYrz2AzvcQ
Q5MtNThddthSIUoO7WsgnYHXlyVudfhOg5Ojnm/DDdoGZ+/vx/vsd/865H0wR3nhELM/TWN3yj1K
zMrm5UdaHeovXTWCNsf28wLefcLaMYgRmpjYPuZQ/Nnn5YiAZiMKcPXuc6o+kxIf0maYv27fqi7r
erPohf64uY7D6NGL7hGFVdIGDdh5Sbcvf3HkGF/Ep/K/yTtD7iViiGKW1GvWs/b83Lssohhlk+6B
/WJHaXYMvzB3g+dRB6QcOy115utztFGqmMb3yp1+TE5jckPXOFJs0wgU9Atw5xXb0MXA9z++yV9w
/H+Mpsyokj2pD/jta+W1hrDd87wiWie1I9P73XTkOT80Z50v8Lo7LkGS5xzs8C8fCRqgKIX0y0QE
7iI3wr9/f06ZPIFN5IWkCBmio0Ss1HkX2P88s1ecP+Cd3y/CdEMC4DIW6s05fQU7vwP1CKzGHZ6S
C8aopEyGyn4cHIIJp0cjEG2I/9DtCcGjim6DkDMrQgD6crCfCrj0y0gbrA3fbvJe6tGyx2IC/8EO
aXBWb5c6I3kfp+InINZvHYFkfDshgoOseUSoAbcFytVLNQ9+fDR4n0AscHWyaYI0TzOca+oMXMYb
w4Hq6qtULt5NDlC+vgMTqvrhgAd0BeVmR83T6wI+sJjdn7r+OMJpWKwhkwOpd3fNL2h9N0UMh5NC
906iWT/Tt/tr4MmditGSFv04/yPd8U7TQh+7fUkU3/JzfdOsirAKGQ2iuNWXLchN5KN6rtNBk6aa
16nAuWIJO/lP0lzDXLrJypHf1wQDVzL/EBWQLTOPHJGb7fMKJ/Cfwk31s5xdSODc/pdEg1Sx7KZu
IimyRkkde/mnzcKskMb5EWYFqIdlQpI0e+/IscoMvD6CGYHaTiX4OMdJWIGjYOIiH9+rqiGBl0NK
ApARUbPTXf/HwTpcYm8e73cHcTBC9VVdxa66vUP45KnMyz/2mxNhI28TqatE41tC/4NbX+5VUlOD
UUsxKmhURcqC7tuPStTLYCTwP0JWX6Ct5ahsGh09svj08WDG10zf6PanwnP7mDWmKjVHJJPjAHmW
25M7omAZHF7fxZIjwuiq3VvMWfumfUIKp7i6G2/bHQXli2WHdDZ1DtynqvqZiCAUP92DvKQsCfLV
0W5DNglWVjTUBvDW6D2vVpboExEgFnNRWHuwnCJTGDVUPXBB3RFp0iwRmzi7nV1y+3Uf5L+sDoQE
f+zkF4RBYVhphDlX7n0idN3tiZwKW2Te2tfPVmLI+67MDdvESmJM6Fl5C8uF9vjx4B6f7agcB0YH
7b2dmYCQHBu63LFj469ta0JFLM1kOiCS6Qyl7P279OVPOY9YYmMYLPySXHOck6FleKqGHL30l7I0
X3LatAslSdOtp25xh0aaGME9Nvq0nCGzuY5FKQlEFDNxBlGvMf//Poais8603vRrIDohwwkjYdTf
1VxqjQcNYUiPY1y6oK39Rv0n4NtdeNz0pEfsWsg4/5eKLSvxCWVBqKw4/RXMbvOmt/15+sbvzFNA
3OdgleiAjbIeL9Xx6HzgO75TyRHuuqoG8XNhHolG/6oy479D5yMcgckEI/PPWOpctqm1yrftBOoB
mu/0Z3c2KllyVxlSGkkdwjfxB54NkJm2FAapXWHinx/q9+iyFaTFHFkNEPjzU93jQdcKjedWdrv/
KuTRRplm1dS8/JkNqJG2HNwzSdLFGciycG+ISQGyIYEefNCftHrQU5Tmg6MIZ2EX+6JKU7yW5otw
eV4WOdQ7yzauUm+3Izgi6pFczgnQouML/b74cDnT8GN8m7Iz/mN+F4W7Y64k0w9gQTuEtVR15Cgc
s8EC1YjuO4e7F7ZR3iIr1gqxpLxC5CyI59287L9nw3G7MfA3ASkBI/UqmXA/1jXNQVuvTjRVks1j
JfymTyZWsrYQ82oBcnb+Cm0QjTxLei/2FK5i1rJTjxEQAyvWow/NR9GT/HwOg/1WySfgtEvTwCy/
4ZeH3WkoRArLDsjPwL7iAvJJ7zERsDWEOKVNzH9bld7UtzvTfl4+GoawuiTbfREhQ/876GP8qhTQ
oxWBxrhuUy2VmS8T26YjfGbSCSO158cPJWfe4WdY0yknMBslJsT6HDeh9qxalgnHYwFGcabh3xki
g5itW5Ee6/TN5r7ntar1Q0GB2kk6lC/kKckXZUVWWTWc1Eyxa980t+qz39ayf8W5y1v0LFuADPt7
/MG+FoEXSOJhZsbMFchZVGfSRpwDjCgSpt2vaxHI9Qkpq1062ZXkfoE2yb0zg0IvUoho0PCLx5J6
lWAaSrdVcR1oot0vgmlx8fS5oOLPYtpayn9Ke9jHmMTqvmY+d32HUQYVK34Axu+VWeZIPUR4lM1j
vEf/7yBej0JoWbaRXEVChsFc0EwgAFP1lF/8b8ZdsGl3DyWa60zs4S/TdavJXEd92HAm5hDmu+pF
e/GOzJX7R0CCQY3r3nK2/KyHXcFfJw7VwIOH499aDN4NsbySjzaUQX3MIC/su9rpGdTK5qszzehG
43u36txDPOmqfSvfjIa84j5DLiZDBGytH/oSK9dwR8fXLnSKv7wxSkocMihcuKaWwXzKxeejJSGq
GhLQ329IS7zFnB89DXVtE8nLkwruy1q9s4rsoZDZ+xCli13t5/ECvaRQiqVJQjH+pfLYuUR5syWO
sUtzu85fdTBejniTaSumcY7kzZiuWZMDgjzmkPAvldOttXB9rDHFyzv/04x5+l3G8hRrocTYAIJ+
Y4K5CsUFyDc/ozH6a6MP2/5JgvsxPZUsOOWLat9/LG0K1cMYzehcR8dQXyEcmzlLPjeYFP8q7UrG
uO0Mz4WN4zOSjUcGPe9OGufCb0RNHMh4Fm6Ng6Q8tbh/rV6ZQHiJj/QW0wwDDlFAC6CS2ajBTtKD
UK2Tsk9JndpXkxvqXzp5+/vOt68XTOa0cnzMgmHhviOSffDXzFYr4SL7G168pAH0cSMmKhDXccyr
a6ElakVfj0Ijs0Cv3ZgtWigwtSgRGMHRbVVEUkKbE/STMF3CXd53Z/CtPxaiifTD+NIKZOvYxqbc
NMpJCCXtPEn9BnYR3TbEyyuC3O2WG4dNq89dEmlYb3WOu9sjdGuNaMQ5qZyvasu3s33pTWlODEMi
XdNxF/GOmBxBXqUepTT/kj6nJ3yaW6rb77zPe1j+Iau5A26YmWMo5+PIME2HeHQZoN3ZBI9yFD83
CY2D980ap17dNuZI9HkipcxLIRFaBIB/qnBXu+bAGCxAjlH+KqnEg5v4tOIbu0HeC+r33f2EhVgI
6p1aX8UguK8WxzD2EXeGMUrT1IkX8NZPoQmV6F6tlP/5wE6BMzpvD3sFZ7STMysDWYFghuDMV2PI
ahq89rs69bxqcLF/uKaMSjrfc1mWYi0jMUDp+MCVGYEgfCEGTk89Drq78Hv8s0A/7Cbw93KtBK/P
9WUcCt2iHh+koHqNVYfXjzHDIBgg/M3/wGxE6rlPymUhLnx0GSYyFExbg/D6Td8oinNxdqV6lKqv
I8CmRyDTfTS/kHap7hFWY2L/s6rEeMcdJqF5aYdOdpulRWITOUKnogsl8Kzm2hyb2cg6nTOK/HtE
gwIKT87IIAs4B0Y7o/8RGAnTx1pkFgbyJS9sRWmcEsW3/FQkWnLEr9t7HoYQy6GobE4b+bvtk1zD
Ad6yF2sC9DSy6mVXjO4F5vchQe/+y53R1wHf8/2iF4bge8bi/j1NLrfOxv8TN+QfhMI3dNr6x51H
faggICCUCynoV2254tgzR1VMeHFrv4awOZW2YMzc/i5YeJt0qz3NCf9mx1TYCTQJLMyQvEnDAN5j
RZ+1xTbObVjvgAtYNepJBpYCPSnm7OkYZFi01A4++WOE9NGkByTUWBvBhOiS+PWzmXLp6p4p52wz
00fQeAgkcbdUIZSxYSGaxeNsdF27gB6LfbeykbLVNuyvjbhfaq3rC6Si2X8pmAaxXDPvM10YJXia
NFTN+T13wnREi99X5UJDbLQBaaDYX7XgWbtooYmKErnfA47h5Gorcf1xvV7FjkKYyf0C4FPKwrjE
CrevOr5UKNa8Y/PJgNj3dd5z+YlqE5tcYlI28YklQSkEHfdfcqHxKoq1BOqUHW4JkoX+bCWkj8x0
RvNnnWQYssaC8g7V2WptUOtwC9EEPqMmpUHIn6cfQGkmnU4DfPz/nkFAojW/gS3v4EtLUQHllb8w
vTx68kplSaY9txw5HRv5NWwjRsuYamCtNLoeaN5TWlhX1482cWMq1teoBL9yyTCFnOyblCONFv/n
xkz1HFIBnQtVeQTiJd4dvmF24MtxTKvV4QPJJHqzNm4uM5htUHW1CmuYjQYXnIwVT/q3QbHhTTPi
woE5B1HOjQCV5Ywne6/FV/aCfAU8Ik1nwWSCs7XO2xWYRqeejScVYvX7Uzq3Kf3VD41/wiWgcxkQ
l2BCs0gO48BABJQo/17Kwx3RwMVnQKRfISm0M+QHbk1BnQvVEnWRWUCtiUU9PVmBeb8jrYr+d5UF
KWZqEWExyAXEXVC+4DWiW7bSph86QsD+cXd/qH8lvgVW6V+lasxE9FRfTfFVw4sYfG+cwsRkkhVi
LnYggs63hrEgJRTOkq5Y0CjQ5l1xyRD6CYDnzWGUYQM5Gj9ZTQdugYtfg395NXoE3SkIrnTFswOQ
n7AJbeLp9l9bEkhT+43Jg/NKz5xaK/iT7UU+UoJHSiRXwvUoa0lq4fvHxa4TmHFQ0gKDED7f47z/
i6zDv2TfEujfuaSqdSRd675F7107UbowyiwvJ1UQn6OePKftldjQKUClqSQ5XTboWQLkyIXcFGwn
TnJy3orDJ0MphtpgQfkRkQNpx8isx95It0XpzfqeIl8xxt5Gr5G7jNW706D/+OfEzUV19b/w3JhK
uGHVqW/LGhEJeniB4X7bAEe3VkEJsfysk0BeCJOxY8jEI7QB4qOcaREd256LI3QQa9l5+R5O6F23
vAgm7jnqsEIyG2kjDI4fzu9I+JdfzIYNB8GEwrSWT550Twz2gjJ7HBrcWAFh4ZJnd66UxMGCbkqj
YY+lK47Sg3GcAgqLx+VrrdhpXnDAjIaBcqFjeJA3+4pK1032AJB1hUNJcoa/zz+2PH/lC123v7xO
NtlRwpOq7zDLTX28VBzsCKyD3fnjl1Z3563ioFXH3ccs0T0z7qru9gTGXG64rVcQ5ZVzrcciQ5tG
ZrE4oA10xpeQl0dIkbRbeTejj128DpGRfkJEkSevY/foeKmea69KaTtotFd5nTsDaj+ksLbeZIZ5
daXSEHpHGbcvO8RxZyFijd3ki5zeccdz1X4FMAqhWdN2ZjLQ6hFQgROxK1k7PAS7MctywA8M2Mrf
JdqWJ9pBoAmBiNW4qEG/6clvkC1KbcJMMauSlEYeSwug+Bad2OWPXX3xZKF2sttC3QBU+66Mc/1G
cDKN+dT3ktfIm//Cf1bXt1wP+S7WI5xiv7fDkubqKIOPAlrGJYvCWoQzbh+n3ya3Y5GdCVE1HiXq
4SotNZ2d+hO2my7LMqumwYnwAwW4NC7qeup65upMyUYl6pqp2nGk+ermqNCpvm8AMsI64KQHgzDP
f3jd4eCenqw45xVRUFvfojiQjSNB1ly3tn0EVCMQquOf3QIutpappTykxd1j78Vdv8wNFakoSr9t
yLAYq/7aIm7oX6u4NLvyDpU7PFcz8haaghEbeqY9l+B81EFg4MOSLEJsBtXv7sVknRhOhJ2/MhsL
LqaeJQ0DfRJxY6jkhtciLBY+gK90IJhqtCmR3BJgUmMfNPxLwvP7ARG5MDEHxMZ/R11kTkUiH230
LeftJnxSSkzaJK+rY7lK9czY1XFuG6PDf86s1hePrt1bCvov0ndgj68pdmO5HVLNeNrWI3EYlzJZ
RSpTU6q+XuY278Ympbh5D8KSzN9u7H3d44IKZoUIUc+Wdz671T/HUUSXLgXDskkabOgeGXVZF6sy
C5oiNoWatnn1Rb0LbeoDCxSs5jR99RRDla2SlI06kT4X1xrd83MXXMrm6JU2xumwzlUy8wSyiQkw
o4su04SAWDLLlKbyqxy22mx1Eq17/YRWQB5Aoeh1oQAaxpZkhCqic+r9UEiSW3INpZgr4zeAVJ/w
7HAuU8hB+ytUWyAbT3RHBjYmrcUezGyU+HGQVH2ka0jNEQ3/KKGgZ9Xxx2S8tohUSUpytqisv63u
QNp+VHXqaTLfjplZJuyqqjGX5Sk8gOKoy0t5J12KXINRIGmuWe9xGFsoFFCnZE+1OVytiS+h4OnH
iKcsUGGZ0W+hUOiYH5PKKfJO4tZLLhyNG+pFHyH3eKaKnW8ceQ0ucWL05Tho1tMHyJAUzYiAzicg
QjQQiIruj3+1nTuFcRYNN+X+ifVhVYEz+CuWfSOt7IkmIuoK+SNurFqMWuhboTiYpvcuygq1uCZO
xiJYLqaW/CXXULYXtrhtKLGmmpsCVyF5Yd2UqGqOv0ZwhvYPm7B7nNuRWJQMoK6mDObjfhLk9cjq
dCAmaMp8MKXcjlBBZlW/NEH1+E54z0q57WY+fixqnmlyCX+Qh9kj15FpmegqzbVcUAuopWklhh44
5SzSnaWahQDS4cv952moHBABxpumIApaCcJFGx1o3Q08ZFygCaQcLbcRAP4nDTfVdhv0jM3HhhCq
06i1Pr/JMAgSncy1RowNFsPJWiPh4bvCVmbCgRH/rYLpFrLsGZZ+4t83vdT2/lb02OWgM5kvWG5B
QjjE7edpH6zS3qbu8oMWkfFufUzeVcgbPSHb4BdMc4ySPQWFwlSne3R40RalcUu2fiqtriMXXER+
xbNIpYQ47cVPLd95TUT34RneuNvRQ3I+kIMwfe1Y0i61QjLIjKkG8XOIgF6I7T49eoXCNDCo45PV
wKzoxYjDJHQtpznRiKcouUykLOIT9Mc0UumQslK+UBtnspgEcJprEwxcJ6f3bUml1SkAA+Yh1x5R
V/PDydBNagPrCAcDgatSQb4/HSNwTqhRGgXqROyHxBLy2db+wPAVnrhajh0AV6GXU110CHqAfhS8
3WeTrj0vzPsvd3JKbfAuWU7kWyprmRcrIfaeIKi7GU2J18LMsu67NtIYQH8CQP79zUEeFsieoScL
YOfziKTpoOX8p2ACn/5GVdi1eims5mkhO5EvzaX/HQaV9TJSxMp+TfVhQ0dWUi1bJxhrUcGjvspi
qLm8k8cm2fd54tFLzKYuM1kjzBCuf62PghzBCgsOFQg0pwUTDjl9awApaKbXWVA/RYTqGBQr2Llt
n4IRcj1aVRG8WBljelUpn2a3KKAbiK1L6bG8yr5mQv9/V3KsykzzE8nmuiLVMMr1LsxPAwjPWSkS
rjTsR5Bat7MP2Y4tzYZhcs8hydXD8Pcyl4VDCnURsW6XYKFZHcr4DWihjS3cNRg0P5rUAZzByldP
zL9ywQF+Ukyo2j8iIME0renJrmI0InCPUywvpugcH0u1pn8qDemdpfjNG/z02/s/1imOBadnkSPL
Sn0rrMIU6XXMQ2rQ5nZSbNViPSiq6izOwXT452o26pscHvntbGpLRrYP+5DJhSV5oVRdisnV3BDc
GhwEq4wD1iXn2b/0LAIEfj4YPrB89IIl01FnRt1by0xKv4T2bmgN2mb5Pkud2pEnlamzyjs3IQ6T
dMEZDjMRzdEWF0qU9tCTXOaDZL+YKJ+F08oJPmaD4rXJDIupfbZ1bcwBmM1dvKGh39WykhMD0X/R
GsI/iI4saZqOk+casK11S/NxOE9+U8OudVyH97sTFgmhg1i/TKoCdNVS10LcN2k0fj+exoprf7Be
+mWDezdpD8egtPMplH4PR9TzbaaSHdFYbRtCn+uO9PHuyuwub7+60jfN6AoorIf4on23CtTwRj6n
z1GGhJWLu/dntzpLwVfTl7HOaFFs35dkEUND8HO5/0BMUfWc8lqw2r7zCSW4iskZ1vHG0GloQ73U
A4V0vyzUl+f8AFt4/TajLSZzG08M+lPbw42GkpLlmscYx8Gl0pcPn3Zznq+G53BGkRXpqIPiHaMB
4fPVZ8/Jzwai6H1eJOl1hgaImY1NuQARvyuFD6Dkt/nz3b0z654hmDw1i1tE350sw2JJHVtn9xe3
5Av17wDse+0cLC/fZdFZKpahZXYr/mUZ+K8mvDGTjZHrmypk1Ud+//9FZPqdqZE2DgUeuAv+VQcZ
khPxLIQY+AYGpOZ/vuEDwA+m7QAJxx0cr2WmivlvOLkgNNz5uefazxqT5NlwR+7fTZnRwPViVFPs
YEHNWBw4rq26ZAA6CbFp7MD0i247WKuaIfo6yOK2Gd/2Bgg5q27UwbLc5oOIGu3N1gReQyrOPgjX
N2zAEQq+qvDjWW02iEfShH9+FaOkmVPf3yr5bmCfWf5xKk0SeHnFPV5lgVp/kJ0yhZZF2CFAjzYp
GZMvrEqHL0kyuq0DCS/GlLVMz74GgohDZoGGnKkRFV1yZFOG/CekIewexYmHaX1jb9BXM6h4BDpk
6Ddh5LZbsvdW31GnXvJaV2esF+nc+tVYZyfYEb3kCzGqb5gc7n+k0VxAsc0wJjRcd1/AtFGob+RW
rsdlNVeIsKDPoarP4zUdT9l+VUa2JjJsXrRZKz1QKdHN0BzZOoZzVjOiahwQN0XANEcnLnkTPvv6
+vU4/gWXE4fFHRdQl0T6MJwcNcJKVv2OdILLOOoSvzKjey1GfVxCB5xbrwrL2PhRNqfV78dkJvQ0
oudcnw/yc7PtUYZKWskHQTVIAzY5bUWdeWIoPc2WOJ7TQb7nn7x29JBxiALv0/h5CD3IEJsVTZWy
sdUxa6qPieGS8535NUnpaQQFLnthay9QYoC+KdEz8Jol6d11bkPT0L9GfWq+7nQlPk8+mB8Mwrn9
1F5pflDkIYyd1L3HiKVHdkDAgWoI9Nh2jdx36NosSVU3H+niA1RS2bT/1+Y+GcD0v6LzCA80233x
31cN4klDJ/MwQEH78Y+MMjlFN8amTs4EeH3d3rKEefhtcXfvAQrmPHzNX7HZK4w/QWOi93KbA+xr
wi7h+jpYtrFsuC8fMd8vfdfX8PioObczIlrmewKpfRafAxvbQaebROE62IarSffQNC9N+pPCPMK/
KObIR3HLJkk3Lw5EeANAoylv49+YycfnwjAXYuwlbEpZjZgbPvmT68kHVCEhy7rGe37LtP0V7EyA
on37RV9mL29XPRb47QGy0dNI/q/E+S30oACeeZp4ocX284z9hUCsWnSR0Ci7TleWWhX1FWfBLSE6
3DNdFCbjRn9eIG7vP1EQ5q8O1z4jcLTcgaygPsDtITGiS/HRXw5wK3VL2xOAXA6nukj2P9BVewCe
nNBgJAuP6jkRpiEfD/MjIUaX1CaD8XThBdW+8N7/O4FXaQ4J8QEMN6iKraHpR303nNVXLUK3QJ43
JoKM/lydhOy0mPjF/XuFQh5YK3cKp3v5EcBIyW0LmpkZHwtIiekq+v6pijO5x/syQRn6ifxnpPkA
nAPv0w908yzcMZrn3X03w5GY/iFkyE1ZK09EBYCQm7ZYZG0i5MzIy+U5bOCF/P2lI8hljbydTMHE
id+WEVFBUCw8oYtm24t5oItlveofFdmJp7YluU4hle7P3o/pvb4Xs8JyBFUQNtR3i7j5iT3TCuUx
e/oyT5V96bbYJmxXHyl3l1gZA2dQXd0exESlQce7ycckBti5hDKN8XmMGUqha397KZ6mfDD85XoP
7klPfr1UCjw9Yx5478+v7lLRDosiboOAUt+wVgsc6nKBtVTfAg4iQ3qPk7nu0nRu7dlk1nnC7l/J
cTgv+N6eLU8Ei5blX3BcNZsPFXb1/IfVwO39rkkj6J/tsOdcp3mWQzffdQpuGEcy4G0RRjyxlMHd
FMlLZlzFqF8u4sNC+6qqZXz9j9qy2+Z3A475CCuxgtRYdcJWV+vAlYG1+Lvb+RTVSrcBv9xrhA3U
spzPtUqJOCzE78uzkx5y6Ztwn2c9QH0bmYGzUT2obIO5HqNjkHwuf9zgGGnYaQEfAdAyF3Y2obZM
3XY9i2SRM1+ZyvL4YyPFM/GQfLFS8f0B2W7XDrCqB1Psfkq4aZT/soNu/F3eS6xoeg5sB6Z3dAFr
UmkUioxDLqNFEMpFDp6zk2xvztDKWCiucxU1yxu/nW7WM9Y4XS0Jh34gKLhgK+9ksFqQKJl4MFU8
+y4PNoC+nqrGxa0qlXvooEX8vrgwcJzMGiy6MTllTfPM/LYAObe1dIGlio4zWhNOF/IdDuBUqdNA
L4MIe0hHFZDPC92QrKxZzVGi8RtE0wQfIVJlPS9Q142MOPPFhpgwmD/v0FSfgfipE+ZCGIOahAmG
sFd7jdixlztAeMaUK2ZeLeiVeT8ceW1LBnUg0HEGvtJ6lW+Sw9Q7zMcrptLg+IFKaSw0zbBrPE7O
oPiwQxH6ZOQt9g/gpEuvHwz5CmYt1TSmqUwblt7ktf5Y82dNT8iKP0vuGeEJvzcUpKUxywIDOlLR
QHZnDsSbBWRerFF2hEDMoX+j/MycciuHIPlxB+SlK/TSQpfDo0KeKAF6TttnUUcmHlK07YgwRVj7
wr95n3+RTq5kYa3pk1FiN6I4t8+RAyrXwL7CX4h0M4RooIL3L0av/mPUaOaveaMDkGEMDnw0tKgL
gqcuzGyGTNm1dh/krADV25Aw8Z3s+dBVhGEuc8e9r6MUSL7BPJgz2ch8Tk7XRy78GW2AGtYbKCdZ
nBum5j2gX+jrUemCI85q8QUI5jvPy01fQJSz0EO5lQNgzLt4w+TYDCJmE8sBUoBpmxbpCbCp7x25
mJT/B3jk/0GoUARarZGTidxvJP8bL7RNo4RCAjUUtpd1qVUlr0KpJt9VHXS/Jyrc4HJIloSjf05m
tY+MLWh7M40fg2Q1mjQ0JdIcnY3VSkDqRyhGTJrW+ymRZJB2HgNzyPngKlatV2MwsawSONXvvW53
EmcQjvQ8zDZuwS52+tharic5vnlLW99YSFrmT/BzCs0E0idV7SYEj8n880yXgbEwGIxcr9W8cG4X
u841atLCaHs56c3kMjs1xh9JUIhQqn1WwkkIvEohxvidEoXT07wd5Gk1sK45Ihp0HWOR63JoVklQ
XSIrC3b8kNxAv3m/fMYqDUyIvxeN+S//UhvQNdYNFpZ8Te2Krr11fxWUbd5XoXpX9Mt21gFag78R
gopaNx1iR18erc8RbcreYE4idg778nh1LLY/oZ6Q24oO6drKtVXWGCOKUUfNXPv++52MZ2a/XIYi
vK2EZ5QAyVOO0aeXH+dZwe/pkj0xkiTT1TOzuPxW9xfGU0d11VO1w17tPaAh7hheaBAz2kN6gD6O
BhtPE4nOJNOyHyV01mZcBvtHkkxsce97AeKGnoMuGP2UPb1SLyzA1+W49C7KbnpyFe3+wsnDjpPp
AN/f1NEnuS7rOOybc5KGGjI61gFpBotzDyGw17+SaIWhJv+/GmlPUq98h5UBhZZeFeG6uqjo09fH
MdTAnj9Mcb89z9LinrAOQmcEUsCanLyw8LPNRN4iAXWkdB47ANV3OG+jyJFiyUS6Eg/oOfLrkLcK
OtI9sxc8Dm9/YBxpUluS6irPAj7EVH0nICl1jA70wgPOmBjjUEZ6AwX+2dnbtBPyUWZJkuK6LN4c
mdeJtaHMFap/XmF0tYUNg5++hU1BhSgbKC63+B2k7TV+N+sXMKWMO05ga6YcvU2scpMkcKyvuUaE
WMpoTzQZ/4xTz05wctJzHVaw8Z8zVkLpam3m9mTbdVW6Ztp1wRXPvY3mmAeuuBo9a04iVGmfLrku
LzCNhmWaa7nJFK05Acv7fw59Uf55Gh33o0IF+Sv7I6Lf9gLjvF+aAj4QRHZprlTMvOJcNN96CUls
8XYn37YcWow3POJYo/eQ8bJ38+0/0Jyy4uOFt7T8u138hdCDZjc/oeoLQkL4KysS7yAl4prLJ1ka
wlwCgL8xuZA3fTbtjBXbj7afY5ceqz2zSoIzoQSR8NpT8hnivcBiUe1hDiqp2y7NOnGlcsHle1Lk
VsIrOfcoZ+HaJk0wAJ81vfJkQEegKTuJRjy79MG8BA0PmHOiAyfwnVBf1yQreRln9UJg5YQ5sdLM
HTCrv3HPqsBlSGojqWOCA9GNCPOUVC9Rimd5dC+Wdn6b7T4jvsOpBktNIf61LSYstCi+RJcq/NmU
1Shrzh8FZp0L6QV0/WjzKsdsSJau+74IYUrTPaUM252cqm9mo4uqqAFDbwnNrmsoqwMtmB6d1RaM
m4KkMk8Un9JMbxFEYU3NT70v/MlY3FEV4zrGz1qMmxuO+wgXsIrhL5Y7iNNXHb/Blege2WCnoGH1
XB08uxZA64nxsIyynJi/gmCdM1MyeqvxJx6TP2YspPMsb97/z7Pci260AVcRGYnSUpaDTQb/0WYQ
S0JAKMK4wPfoTbz1sZsXwevCViqvhL5zUwCRswq/OFSbs/aFgYgLU6J2SNrV+HLIDIAuHjP8mx0t
3V4HtZiUUnlHTbB84rd2qortmfszXTK/XVZg1zHDgd0MhEhWTG1d7FRNe6aikZS0GskhXSZXF9tN
GGk4xj3vnVUqVToMjCHAf2VnV9+VR5DsnP98OUO70bNYehuzl71U+ZBOHzK21wrcQDHybIpte6ac
JQMemRibLyfMH1jXtsBtGIYzB+LGzNvI3fvIkpXs/KiWQg5iRMKjO5+ttPBr2B7zzN/HgakIj8Ky
ZtlZu2hWDCVBqIYJR9j0s9PTXjHK6tVUJOi5y/yzDmv95cuK/T+o5CUF3QTi0a3DiFP3gs/ZYGCw
3ANhPHP3LgQJeT758keO2wikbUbaNCtoUHZYIVMSIuLceBi777RyQT+bxw/F1KyW6xS/scoxB8cS
1zwzyJe/QjGdwAbJeB9LCo6+y0FXRMktCDe2+Pbvt1voF5GLmBCoR4foywAE+R67nFWV6XYIGVjU
xcwjQ5Dhwfih6uJkp6MEW4zwQ4g+T161oNGyyh56Op26nmurkQqJH/uy20/9zrGesYaUR6II4HQh
AdN86h9aZ2Wq5OHeJnmPlMW35ul8AxAf4hdTU79Be+LA9LpChqiCUz/Kg1ekbarzsOkLGFFXNYlz
f7GlPPjkkz7VzrxBN4gPz0sx16E/SpB9j3LtK+1uu+ID1U7hHZc3fQzwkG8jMLgLQjSLj/+hTElb
BMIaHPpF42riMx/Kowyl60PshUYEYlKiLf2Df4uSFAQMxAF+Nnpewyj00nwUDJlfWp1LI1ft0EmO
fOC8/nw237/0HfVrMpBmY9YHLgxeDtsCHGe59KO6A7tdWZX4kkRj2B82YOhOXGQYz9fHuVeKaxDf
59i1g9CuwddvAfAJIeyIXoiFF/C1pX2boyuKWoqO5nn9nkr77gV4Idblh3cO5qEuXB1k8nxDXGbZ
WoIZ2/YnjAYZn2R9/gDInLdUXYEnrUQZOgqMMA66SSwOJ33+pcbJN6L6p77O/Up4XAtNk8LPGpsr
oErn4DOQTpbRll6OZHgLr1nUZuRU9dH/p8eINabikpIVSutakDLkzOpvAJCd4ifNp8gaHfVYf2gw
FA6tYZPEi9RgU16xGXVCni5kZJdhaSxWjYrJRW1185sJ1tRx11MZbX0uBqH3Q4dhU78Ap61qVVoG
nvwvQyRA9StUcSQ/c21pVhUfwzeCjmJ3tGyyxNlJYHsNIUHR8AaRyfmnlCpQUKchg2i41aHZZW/t
N7A40z9zPB0b9bVoXXSvu8owcX2CUf/JHEVY+jTyzwv1N6Z+BmEkYgi4RO2Y68tCh5Mb3g4YqgcY
PhilwV+zUktnr21yZLKJkWYl7BG3BrrpZ20x6LdYsDUMmQHgrFeLrfuq7tlwOEMzU3kWrLLPCrdh
1Onyb8S15sUUdI8vJjN//IXs0MWMT9pSWAUtjNdR7r4SoEbFxMm1FJavFKcsnmfB8+tvstDW051w
gtVYnCJG/E7n71J5ms1X55HFsA/zGbL+Mu0idw4yF5/DdLyx30J3H4RnPtjhG0eBWEfG5SK5GsVg
dNzrtGFscFpg4UPw9nWB6QlifXZn+EYGbqi/z1c1EtNthWwEq5LYkC0pyMIp4E/b8tMd+U6MVYMc
eCSd0hP7R9JFD12sZt14WbpIhxtRorQu84Jp++iFSs2c8x+l8dxBFJX0D4GBxgTylfMgkidvL1X9
KHnkl1UqFHSVoGVstNqQTKuwWQe0PcbPEL0yYQsfQzc1maZWBXz3+NDyd+r5XEZjA9Re/ne0Bxys
vrmpwAiZPG2386COEj4vtHn+qYUfqRBNa1Jfz1EGK3l7a+lESZoOrHtbdJVwnGappBpgw6uLLxI9
WMG4DLkCme1Mby5NF0lz9R77Vygt5U5eelffHA6Fi5l0N5ZcGJ1WKFDgpBBxXZhITLN1sthngyk9
vxevtFwaBLduHdVe/vTwfwWWvntqQjFe2vOP4+igZMcgZyOZEXIlKnb+8uzwymeyAqokRiHpeDW7
qAJSsf83Qt243TenETTaisKl0Ib7ZXjxwegb7Maypu0nHRIPEtffNNnwMqkaAuyHH/4DGDzd4TdT
Z+40TACTN336E/k6FWHK2X/bA1XVvIZkVbTSz17FwaooHoVQx451jaGuvyA6EK1PkZzCragGIUd0
T9o5UgQOgEPGf9UN/GMBToJuK65zfapgBVUwmBAWb+qkhN2cHg1ng2ilAcoU6llgUqnQttFAvmel
5JfyogBGSfU8+ALzouy6vIjEPB3/iEwR1tJTCVminfOmJWDE9Mg2gR0c1aySjjH65JHgh3cYyuSI
MgR12J/pixXSJ2Aqr1FVPxZ+MmAc8rjEmCS4ZxOZlBCsg2Qama/zy/QhtCmWS9JL42O5BS3LzPOQ
wkcqe7Mw/xppT/CT1bVPV9zL2reYdyW6NZZH5P11jaXjw9tSDtyOv1DZNyvNvdQqEzrt8UTMMpZK
wTotRsjyqA8fApYwl7kdrynRxlmfikEtmGFyVftsWiC75yxLShr2VlinCZp3DD0Es32f4HnLY5lk
KxA6vqalY9WsOkyKmM4E36eQowTdFEbVNtqkI0HbTzRiJ4ErarpWvV7Vu3LQkDvWlumvUp7vTxL8
gCb/3dh6mxgO8a19M+vrxH2z46Heb2BbW41e17QZuXyHaxV93tkYR9alSfIy1GyTB1lewRV3UplJ
E9937etib1OKvgW2slnU0vwAyb3TfY+UCTt1xKMAGo9QLzsk0PXFxU7Y9kOr06BP9HrOLhjYAXgO
2IXvBrx8trB3Ztme7BnuebqD8+clabOJggDEYQFsvINHmQU2JJLQ1G6HUz4WhyOv5Lstg7QdSJ+T
I3zsMPPVMTzGNmVIcetenVJc+AuJFweh9WdgM+BCozxRHavEdjhgpp2bAsXRB15JlZeRonhMbYYN
7hsSB2KnNWCFSQueO+hT+lNWrR4yeDvK08oufxRBVlb4g9iaWSoW74th5FDljlfW8HEbT2WkiA+B
jbCZuEqWu5/sDyl86QIIeLx+yVYXj+sxg5NRacS7Dr7ZOjCW8O3vC/00eDaSM6b+QuYyFHzN10v4
693WvWW6cm0Gyv8FPOLDqH0i/ZMy6pCEJoUdm0lLeeM7yJYFA/Xc9Wd7s3XQd2+D7K5+z+mWgO9o
+0Bug5YaaI3LCozcG2WA3B91OGff/9ydWACILCKs9UTLbY0C5K8QWyvTRKBXHyamSv7QbQ+KYjVe
R9FR6ZcjmO+idSIMyQxMMY3rdqrhcFL40lQ6CUg5j4P6/A5XltIVtZYRiUm2Qcyj7YHVkVUs96IL
PmNSgm8OYDR2CKHn4xHNS0qb4aHyFPHH80E8R1uDaWc8upYrrLHMM4srFzj2euESMVQlwEZ+KwiO
hLX3t+/9nE2+SKlWLJMdY0waNs6x635PfPwKuB2GA/0DddARTi9oi2SUMt3amKvofhhokX8I1gN6
6EiIlKNupy5pvDrwH3I2udrpbNwUg9rLpsfcEsqG6RCYSny7VEkLcqJySoBvWZE6ttXWVX8tL+oD
8kQHRhAgXZQR6/IayNyV7aO8NI2iWx58xG+S5yfKSej2vN0DcBSgnzIEiExz1gWxnfUZGlfHsPYl
9ED+KT+HIERz5VWECJKBLXJJ62Z+M749gCoKrHddLnLz7HLG9K2qNzD0Dq/EqpmZhoqyhqa+Ew2+
pMOtLRn32coEMEg55btI+ahG7HxW1h/tsMGuEafqE1k/jgZcAlOKQ/lPEYW9HiWelyIo0Fj4vunv
kq3hOKFE2S7nFNEqn0BA2fdX1iq4swgaJcCUfKP82z2lw1F7+o9exM4m2Jq80xCFQY07R7iKzk60
ofXqGbrOrKQ4hIvikckFR6qDm657nIXr49SJsEK8Duc8XIQwC01n7Js7Rw6jBygCzBKkrJB5x12q
nyDkuKnwXz5ygM1ithXJxs31Cc6/IPL8dQc9FCz5Df4T7i+O/a7LEVVaxHIIkqcTHnCx1HsBm/Jk
MyllM2U72aV6EY0KPfcd4/sGSQMkrHBHHyFbDbeJjhsG3RrrL496aNcZb3cfrDnQWJxOxu5HMc0e
Y0o0aNR11jKIt8NYjdDdRqFoeZik2g+5FPxXRY1SKljGe1GTg+l7Bmd7K0Kv9tIs8W/R2d0U4OWj
lQUkvNbFcb3+h9UgAxJl0kBJ16AbJZjriyIbEzsG6tPPJujpT60Vw7mVHcL1pWBY78bb2MufCB0p
cEblk8v9GwFyDuM4AK0prVvi7cs1ILH3VMF102+k7aEvAivs83HOAXNcruEi4KF4QLx2oLmq3X9/
3VrmM4ZNSVMcKmOmyv6tKQOB/qhu/bTk18amXB2pLiJa2SJFrlMB7EUokzqyO7lyyc3iIp33o4ts
J6H+n+T2/Z7W4NFpRQXMoWlEbpiM4NXxDwaNOiyByt1gniD3GZIjvUQuWr3gTYFrYE09KKhq9hLY
adDMlo6q1qwg3KSlJeFp6H5pjJw4b8ctHRcdZE3CnjguKktPdjqbaxQtUXPYCUUppwhram//Lofu
WgXRH7zgW7+r/lzEWjQgqrFkeD7jWrSS8Ry28PiatmMZ7NxH0kBaYhKVTvpsbhKPYbSV8A0Kda3a
AEK2t8rezoKYjhwPqmtrQOezRpTn6wZxGeZvQgNGZ94P+igncm8cUU3lnU8ci6g+pqwN4QdyOTw5
aC+Z1vdAAcZsfwSFKPiC+urq0mRQDu725imf9/A23guN7QEbhTqIgcU0FB3AJiYN2cOzhLmguNOF
SXwpivEXFvgaOU3sQzN9HpPQf30yofwWWIOVzydx7IG877VP3siZmtOD8p4UQtxUTmsM6zS4bJnx
bXQPYwZ+VRs6E0Iq/MwtWSPxPvmyVfgDO+sSr3KD6GyiK7NTUC13ZvENaLyEr8s/utr5clFZpK2u
2uYs9nHhC3Lhy5gm0SO+7z5+kfSpVGtwoI8maEvOGL3hBXVqAvYeZ5peM4O65EZ9TCKOKwgtRQTI
SpOkTFxNxWRTU8NMmVrn4OJbuFVGFu3aSWQHXeZh4XPvp4mKTEfTml9Wqu55355ATJqzT0SvSCak
CmNV/xjPgRdQX9EY0Un29cBcX3JuN2eX9om68WwO6+oW5FVo8z48PyjEJiKr/KouYtLMwLPQy7cr
FW7wfvUjV+sH+Ppr0c+6Uslc7NOMbYrxRmAN88W0VN9/mWK9jZ73stoJ1xALZj23pe5V1vdzL+XO
sBN0fi2PfiUMwEwcfbQ0sxs+3iCTnKVHPbp9+6T+oUDXsTjtQT9qXVffwYN+5mw9Z3lJ6JwV7tli
EAs/2sXccMH/RxMqQ/uKZTJArrxdbe1oR555RiDtOEowwPvvN4alrvIpwffpXbE+7vk2ntEpcXaS
AXl0H4VYu4brPJqKA0Arc78N5yw+XXjARR3i4sKCgr1CX+oLIXcNdrqWrPT+TGZiwRJ3XfcgLXOy
5fIy4F0IcMEs6qKZVhBW6FbDNdn1peXkoioexOjZGcwhfgikf0MGjrVknWlThd/Qu4mx8uyTXbpE
dxri5wefpg2kTwNbcYI2QypER05uAxk9lcICp1Y0oqOEVnxLZk9BUufRBkhcaemifKFSaRaJrfuJ
UBIOVZRsrFla1hii3FpB8aBpjAEclBNhZ5sr23NYBuyJw+S69LgZIzefQU824mcBCg1QIq2Lq2Gm
mOTbOVF1wSoLIh3YnoB6Sh6QUZFTNSGGS6KkzXdKVjl2dBYz+1HiqqdwreWRQrHh6eiFxjkWiI9R
I9u47azH2ipYR3mt6KZ1KaYA73HB2WeFSADMRY/l6fP9iNbYsmuZ5eVPIZTFDdAcErH8pE+aVGQR
6s6baHg1u45fGfGFilgeD6pgetjDE0kHqmcItIHYw5tDaasGFcodF0bBEZCZiXlqhWq/WhgWvcG2
+MI0VqWm6b8edAimvSH7EuDGbBbxPZ2X+ovX4wmFsF73EsPedbzuzlcIE4a9SNoLp3H+G5mGOeBv
TmqITi/HDDzm8eteMoGRYqpjNusUjRNncQr/MmXu969nZBtrY/2Hfc8Lj6+58oaU/2YCa/PL+BiK
KI7T8a4USCd0Alutz81PikH76XmVC3aVrWIjhwn2wm6+yh81TFBDRNoo0ISBAoqXVcKmCNPbPj3O
XQfPGM7mWdD0TQfyO3bpbgl92YEG9J0QPVvBZJHlPDZmKbKApSvvrbGtF8Gt/GsL1wLcVsDvUbot
YEhftFnTA2D8sC74uhFYN73ZRdUeP6qf1pGw67xuRdc//LIFMLv4pSI8Psb7ihAlErNmRWIWsTQa
9vrPOfLS2o+dZg6PvApBJ960tD14MKvxmv3ekqCDWh3lt5w5BVT8eLtBx2LqYB2VgN6r6UR3z38o
cIL0V869VO1z0UX+7KyIeKYYCYw6FC3tvg8oHUXehKhg/X3t8rGU+99ZxbjXE3JF6l6vtY9eh/Lr
r1kgPbvTXjT6c8G6at0wBVWwoR3Rew1ibAsi7Dg2zAQM2TZAS5Vz0qqdgKgIcF5KRmzYcRX7lOhw
ExIbcUzpy2vhP2YXAeL6omlMn34OQ5s6TGRT/VyZ2dUXSetOX/Xz+IG1PFcencTczoNoEh2xgnoa
IhhICyCgHrl0IDfMN/1pfTES1Gaiv2uQ+e+RRD7zXOW/U9nVevzFICGYgAgF2dbBwnc6NVkAvxsN
/E1bMMxJBukoBfC82GozyiQ95L4Hz2WjwVhF2kVZthx257vgNuk+KQPHT6lB2XtKIAPXyl2owWzz
C8unJCjcDubfpYel/X35HBWaalU/N+hSxcNJHpNFFZUgmPxXILQOr+CCUB2B5fn9xhz0eNh4S7AR
jy9DN2Ewo7VkOxYw5QxyLg1bnwyPholYid7x4zfJntq4bUe3wVM3ESKE1LHLvFX7omZpNm8nh2Uu
3NduAC91sKsN1cfRJszGswAk97Z3UtInt+wtNsBnanX+owXkBMB376Sh5hkw2uuGVLtBJMpq0lpG
eEyYp9nqWAGsceQhfJ3lYuG1d6cHfcoIUqIYZMwwLV/QaUh7StdAsoycXucY53F/YB+Rkcw7hCK9
tQ4d19sj7hcTjKOupqkTl4lqCnEdPFbZc5p3PVrxocRIaivhaR2rvLJ40UBl8A7j8VYSpTXrGBi9
PmS05RhfzQHBDuL8q8fVl1B7fUKqGhOrnYbNWoP+GgopqhmcUmz1c1H1h/qTiV0rUJPLS2xV3df6
YFnOA0XVow8DVEDa10OevfXKFhNBTrNB9v/fzcpqZNvlOAH5Lp5o7oc6aV6aEgm1rz6iBl7oQ8DG
ysQcR6oJEGFyimSpQ5tOJi7CMNW9QhbrleKjnVlwZIVjpmhGZ+o6UNmeqHLkyutbtK5DiwuKoaGj
H2P7a8d41PYxGE6MstnxSBner7Cnn7Ue776JHKuDzbHRjCt8+pc74C2q/Sgr6HN+BZZuWLcsz8LV
y75RnGucLxGak6GWGZkXUBWtaGRi2dMLrzuXCsYLAHoNFzS7VNqojEm3bTxsuaSL/6vIGOGTVd8G
54zdYuuZGQfRdijvxX4WrnPxRRKKCUv9HJDpkUVCfzZ1W8UXCuXyIiEvJdk8y8wo8x6o/QsnqxRW
VJEwenoyzaTiUXclneawvAICpITRvOmVzL8OYHBMPKZl+CyImn8bDZUfW4j5ERLJkeTa8z3o1uAY
eCF391XsT7rLtZD8A4frmTg1euQ01U2hAO7H656rA4GJmNut/97JS6K5O3pt22Rmtf2CZSxq7KB9
6o47dH7Bv9aM16hFcssT9q9r+WSb9EaeV3S7FS025GS/o7riVzcCcnQrQJXWeOiciXaHsezeAu5N
AQXYjAXqF51L7HXSZxPJYsH7pan0ZPwHEySA1JNQBnhcVekBzhv3rrR8XXz+FCmqH1pjlGabdojM
BLbWtrEzLP6UoPSe0iKlGlrHwtrVVcWcpYR7qAd4tBmNE06Z2yCht/4uRbvUugX8CMF1UtcZf74V
rHHYwqhrt6IGTYnypj0kKaFZhcgZ68lIT6PXNyveaw1nuyb+9pVrSkdOQa4bMptVqiGSa6itbHVL
5gZ2cfXPDMVcC1ZcgK291wbI236T70XvQLh3Iss2uBiuk62hLQ2n3Ccljh0XCSjkI3/DGsiLENrt
D3Dz+Xs5H8nFs770SYSniaBskFdi0hlGpULlwJ759Sg2QK4PcejaYz/VgLBEh1hXz1GSaqErH5W2
xH3+xVd2bE2tGQz4E55EWHJ9XiRlSEVlgKejdx10WPezcv48/R4Jqx0UTHpE+a41GWW9ok6HN4oU
wRBF6BePeGGDaI48tJlGWg4lqTI479Lwy6Lklg9n4Ycp/Y/9F+Q+00yQIkIZoRoDbM519Atr4plr
CQT1dSg2316zkIhZyU+lMJevCetRghVySuGdJ/AENN82Jlhlq6WyuZOD6djgHCmrDTOx1+PmKm0R
ydgWPBOF1ZO4KO8TQHpvt4yyE4KIxyXp3uqOv8rMU1tRAaqTmUlqR6EZ26VU3rLt0fhItWyDuGq2
doXGpRjvkXBXnZHV+SLSfHBj6accs7mcwBEhy9CxH/V27yVHhlvwKkow7lZvBnLGsDFkd8ffCFoW
guCbdhUCMo1C2Opdc2vWiroLCN4dMct4pwZnOlbNlMHFKf6lNBD+CB6tLpKirujp8idlf/dpl7sJ
76Hde0RNJsYgXUOJD9y4l/pLDiZh+akHsdoK0HSdxfbnuJ9ozg9sm6JuPtl4E1wC3Xi6LlfJ1z3I
cKrSSNmak3NS/e7U2recw5o/pM7zONJnCP4RQIKa6tRbT1pfQyNmKBhd0HHhgJ6B4jmDU9GMviM8
1TN1hXpsNgc4IyKyzRPmgwjGbFQ7fGS2jLg4XY98iJz3YCA8LJ8gpRuPQODsAUNNAPACqninETmt
LCsO3csbXef3FIXkum4yozLhdGDlmttR7i0egvqj+59RkSF2wtcIrmKJUX7Ji/cuYyg1tdwzl1/m
sttqhD4DjnpZdd9wsx1vA+7iTfnx2PvXvsTy0yLQvdCM+4urYkBXzXcdXPDAfs7tUOz2q+XWatNj
tkTzlTIa++kxj7MhiO1D0oAEHdCGNfkWQyjJKq69loLQKfdAPeJNnFE1iaZp4l4SUAa4+i268kVJ
JTmaPRtH6SvChndrlW0xiRGvIF08B9ZrudOmVaNUlXnLeIJgqm1oKLtuIqxk+Dh6QuIElj1wENp1
4Fwqt8SmQiaFdJL73+/XsT3xP67i0pD9oASOIMmMdLwXFSaPaQ/NH37DecSNSMCX8wD6cpK2jcJJ
dukt314kKEhtcSdLQJnUiMeU7wh+XE/0tk+DP/v7u/U0N77U7JGfiDGiLVgD4UY4UyG+5X/iOFNo
jZud1KwQlbTQHSvOI7GLrrXZuQLHvTgWIpOQ/a4gnfJKVT1EZOLOj5EwIPQmm4ib+NMuiCPs7mqd
ROigEUoIvzdWaTqO6CQ3aVa8KVgP0NeBvgQSDyaZwxHKg40Lyb538aR+W9iF1esxz/O+SjGhuvJf
haof5Nq1Bax0T0+GwcPbcLQ0E+4va0QcYdUsm6sLdAHyfnN883BnKa8sC3vehWXyZSlDojDdtE77
6KM8ZVnT9wFaS11XF18Z9RP5M0K1dcYCxWvKe1LPEryvOY9lJUoJIz3ESIOKRyuLHujRFKXYyO1U
fXupekQ2nz5R4ejduIVS7U0G16h8Ui+pmH+/v5szXY01zamsDja/8UDgCh0V7rpwHGGP557HJGnH
Uf88Ki9pYhZ0/neWohr8VkRTuJBZRqo8lLKrfQ2q5F0DP3pZT5Y2W8JIbqzpRpk+LE18EH7xOL7K
bxk4kEv1AkGdghRVe8GMO1iXSmmnCri1O2Q0IgvQQr3v3pCc1nAV4mIKUdUN0DLEaybPEAz+Ma+H
8RwlhJnWzCnIHiG9YlACaMf2PmirtwuiMFsp1crGQVMcjyq+QVmr4XfJZeRa+wBe1EKAStgS5PFC
F64RjQ98OCY3yygDYxHE74G/aTaQbqhJuyLfEHMHi/T/nPNtKeMqjwoeyLtYAcIn/H+oPnnffNw1
IG2Dh+Ce8lGlMdgLNpd56h2EtCAAjWUMwkxIiPYwVH1Cd3nt/D6+2sGkvBy5OaTg9CdQ9pRA67Zi
YBF8uwcfMy4i8Te6ocybf2NrM+X8EiVT7PSSxNya+Njd6Oxi22pXChBteyOep9YHsKoDzsDD1P8H
vM/uYNYhZWo4n2Bgw3/MFB7Ih4WX4o0J6TnZyUTq+Z8tEDikKJK5HBwD4JeGIGy+jWJzAsO2VPnm
h8u4k9IC0zISAS0tIf1T/bIrDZumMBTwQExoveczmKqnYdC3U23bsd+YbM3Sbu9lvJMp4XUpll4M
rMhRqeeWvQfrpcMLmIibFnQ6iZ78M9uKRgqq6sNMLUAOUG+dQDcU0hqIpILmkCYyy0aQYRScD+NO
+moT8H9Gck5Sj7OwfeMrTeSkpRrhjZr3ABsjA8EvM/hN5e5EWZ67GftVAWFAgD8P5QcleQDfI2+G
cXoOPwJneetQo1tFHFK3/SjObfSiI9WXHLBH8NWT6gyrGUrrkfmItWP7Z1ebHE3cfRATWtS+iWbY
wD3F42+rqStX0cWTJrKb7mPhmJH86XdoiRif0lRCnJvoxOEXjpGzN9vnl7JrgjgokoYVz9oomcZN
2u7fh8tuI3aZd7sIDzN3HLxcTbrCoUAqw6hR+P/EfROOyKcvFo/D2r3fMW9BWbJbslIlKM/2wrWE
c+u9WHjbjqqqNGg5qsgg6plHrA5lpnL9oUs2xf9buS1BLpYhO+S5H3TXNNILeiSMl4kxB8/hEl1n
vlOkb4IdXOVRY8WsJHDLV4Xh3H2NBPK8jsmaxWUDlSUb7vufMdFQl3E8D1FPOO1oazNqNRJdBgIa
2SpOghSr8FBwnJibERAUaUNV6N6RR6YtCZrODJilyHZNUHEi4u8UqHN8c+LAaUPifUL3Pm1t0AaQ
Ey3eJ42WbFy5oovJhPSImUvp3bvbrXj/fyKQR3wfbpSTpYBFB0xMtKwwuRC6yJyXXMisL9XxWsax
gqT+5UFk0HcoCdYGA7zeo7sb2AtWhVBUMauU37HbV5oUuTnORM6+6OKJ9rfjan7fpEuAWJahqCTJ
xjGbkTJetK/ey1NsHeOp+M8suIPB19Z9SbHGBeMG0cD0Ohob2C20t7/fXgXGrLlD4fj+6o+hYy/9
3t6debTd3kEYrThek1ZKyf/glnGcyRPrdfWSrVzjfgfMv12iijhMZTZURb+9rCIS+7gaIRwtK5mS
KqkYe3K14WnOSvWwD2rISbOL4AtRRLlWW7+8eRmiqsG33RR676nQWbzP4Pm5yA22jPgnJChCJ7++
DUFU0eO8POIQd4e6sjTOFOKJDOjj7zc4BS4JNPh2qXXXEhSogrhvSYKWsQRis0mqHERqOJulmPOk
eLPAkJ7nsKut6aNrZLP2YmOo5VsGB3rJa9q71+gvtZxs8Lfxh8WiH+HSDcEDDP2VMJyDWBI/eUDj
kThcsExlV+XxcFm2slTUKpZ/Re9dcmcZAheuD5lNRlWzzMj7jCvzUCbQNWnZjD1Y0sxzvgsZGPRD
Pzr1dlPFDpLWAW6c791pOhH9A6J6RZvcolaBH4peefKkjWZIGLR5yjCIaVrqxxgfZDCXO8W7xfhi
7/WlyOn/IUAPDGmoADRJq7wtpnzoNllRg4MTnVAXheA01CPzKS5VSdyn57F+5yc0IOfF+vicTj4W
3QowEjQ9795sIbvo4QHq7cVlJa7hBJokbYaFnTbU0uhDh3Q9j5oQnUwt8bH0O+iHCxRf5CoT3+72
BCGPiMdf/mHVQy93JiccHYZ+Y+ExnxS6BvixXkqSRVAGJ7y99GGykey3/zRirv5YFkTgFcrtkBht
66Gjnse/wU5bpxyXyyiR45Rnrl44NXGwHF9LvidHORxLlQtFqdC53wdT9WVowK9zF4W7p+Z6UpyK
JvbJoDU0Cd/YJRyWk41YwSMpdm9zz3z0dKH1NN7OoYpCOghLDBxhTGnE8qzJ+GZ612WkUpdMoPep
0Rm5EERvNwrHqz35cnFN4I+sgLv2A9DYsvuZVLu8y6uwjOdENXd2m2mgU63b4cxrw/tC5sBlYw/N
51kBnTdtTSkLEeVV49oasZZ7gIDe4JCVPcO9S03W+VgR2//c8B8j3SkKbz1VtVdtIUn5GWgVLJxT
JSudrSl1DXQ34cjhDCP9Pu7l8rIOhqtvAkm0xIyXYLZ98wHSzTZ2mVG7htuj+FLoVRGQhrfGiILP
eo0BGltJA8hE6jRjmCuHWp08QD0Rz1TsX5Mb9y/C5kVRZPas6obV/51otp/qpbMxBTLo2hUTbMBu
k53kFsxuWJNOB4kvRokCQrTvNXBr9r3pyJLBni55MnwfpSmB8VAecTRoEC2lSUSMfOnvpiSz45vB
VXTuZOh2//btS5Smeya8DH+PxSR2Yt4M4GCCuE4tr4FQcqGikFyAK1fQLxp9bafXewwEBMapIYkz
P2HL2PQnEAmP7N29kiYN7sHrvv45jF4f66rYvUdxNy1Br3YMSv9/bvShxWfs4AcdlhDMyhGpI0h3
nx80Jk8JUYS8unuD77TA63GSYaGWG+EIr0af8M1XkAoXle/lIP+aAnQrIV82RWdLk3wts7WOeQu9
l01qJ7PSgwGq3eOoVGLIowOjRVoi741yO2DiQ7Fw9qS5OG+6n6uvn6AzlkrZnOSIiOwPZrqdNK/1
DWCRMdOtH3Q78HeCno4jNGwVArV3hWEQEto5EXPaiqxR3ypsm1zmkwVKw/xTxtHEFuKB7Ut9ahsX
HiQ3p29DEDtwOjeISGJxkCXBZYOv+ZX7ERS/9OsTGs/dgx4L4oN8pC+vTlMXIPv7/c1UFFtniwuJ
NDIdgFjKGQ1DA8Aj9kmsutw/IWfvCnuBiPQ3IhZ3eyUph/zEJCZ8gtpWog5QAFXMWjuwvo9wvmJP
7O3a6/dthceyjDOpnOTf6aHaF8W2owP97h5JqHEYPneXhWtaR4igZ9b7ZiIQN1mClUd5wNG1jPJr
bQ8xInOVWdjo4HPzovMR4hdC5aF7wnKqFYSJhQgR6jePiYAtwvSFCgNA3Rzi9jWB34qQ7R0VIJge
w5bXhxJjTv911fSzWcfbdgjnIL2eVAW8tUnTjsGxDo+kx6E/YklDXmCY8jHaURJ59hymRAe+II30
qCfXzTizyYnAQfMrALcglQOFRZRlo6dVPRdymPvkRSrdXNz3pCQUnb0w7qRKrI+KE3dd1ND2S1k+
b461PiE4me066j093IDJoLXtAx/DjZUxiuC6ICrcjGUTYJZ61TedASOxBYGWFkP1Zcti0RwlEBGX
YRhy9ufBmBXfhk6wuL1YSYqCiBfccFdySI0dnYTBmUBdNHcRKDSIu9pgS8t5+TYEy1lMeJYS56hv
YQE75CflvHRcbBhPB6arvJ4ZDy2kiz8pm3foPkxvZAypFenGkox36P4RsTvRtgSiaa2pc1IXI5z8
qkPbg8+Rk9afXzg22AX6joGAzF6f3MW3KntZmKVktHmQCxN5+zYeS0xyMyP67IGp2b014okt2Rxn
TxauwkPEIskcS4EHChJTUuXsmLD4/3aqUPVE9Tz5rFdO+JEHxIDXxTbfW0DwpObKvXuANJ9lIUba
gY0VD2jcnIWSaG2UBnWisSll9bTxy3+HD/+wUS/SaUZpdM5KrVWv08xNW2FBvQTwAOh6nIu0Nmae
YAu/df9Yb5qxjHmPSEhHOSDjmWYFWi4jYiVn8Sh33M6bdNUDjc5XNE2/ofirbD0LOTzd8IZ1i1/4
/fquoSb547pYs4D/KEmyeU4MiGcY5+voTsnwG6B/zLtBe6pFWl1ZaaoFDISOz/XpF5qLxjGIujK3
Sw4Gi/nH4SfxmqSC6qbwXJ2fqr0NI1yROgc2VEZrm8GyPDYmo9xEFWLSXyYyuwyLjqUUr/mMDT5z
oYrKjV1NxQ7WnvzkMP45Ty8m0k3iJ4DSdoD+bKYXBZt/Xp2koaPmVjRkWALbKa8fmHHWYdA6vUqO
9hBv3kIW9FA45RIrCH3T8xO17+JD3vQZuqKaIwODUkC1BkIbpY1Cq/N+83ecr6XZroPuv225er3a
AUiP5Dnikqn4AujFlfR8ED5uQ50DahYMClr39d9Ux/RDbb5UuoJNFPwgCckPDA9ifNCbBGWaVciF
p9hj7gVSdgsjQ1iNr1AGoC/LUml4a72mO3AWO9hwqkZFR8MdCgdbFQt68vRnfjSHsuDfAZ5+oiiV
9GmTZW/XCe3K0JfapbwYjPVCkNDIE30mu3NrNtVcHRRgGFxsYwxxq+BFOaMU27mb3BL7o6jfq8EE
k6ZXmnTYbfQgL5rl3JGaEK2R4tXAmO73mkmiWjFxKNNpXITBIExpAya4KWedYUYJJpWZfMp5GDHg
2ft0KCwPfxhkz9XNkn5TK9QCwywSOnReMLoLAYAzfjq6tzr8d2DbpyC3+1mYyVN/7Topc0znomkD
BZVfqCySiHGASYkPk9Fq/deRlpF9bqavG9jpup3g8qJy2Uu+H5BJyrSJMkaOm22S951XKtl8ybHW
+Cu5euh92zDuhZf4gldq5+2kUYkz+4xoWlWs6UOOPFd93/h7wXp1ll2DbdKbDPUXRgxfvQXz9ulI
Q5+WJG/XLS5VEXJ0Fw5hxpCNrPZ8E+phrUylBCFtD60QczLJ8550yHmfXA1+88QWWVTkotwheU19
M8HszjeUZipKur0WlwPRZOlswNt1bVqakH/SrLtvI/CndB7wI5/D7xrPoHlKTHwVajZwpNGVks/B
OwA3qLHrVA5m+q4hFOi77u46vnlHBmRSJGEArWsI2YjCApAt5D3yuXAWSX4Jdjt/yQMyqic7+F7O
VQSJgQ43c1EqnLfz4avr7vKNKYULvbP7WkTvEHFMrPjR1BekwkJ7/bGaJYRyz271jOpTG0YrBnf+
y+/DuoZ1B27r8OB5mahb5BIYYOKKHRv34wAntL7sno8gKIOy/EhHpIJbH3l//199FpZS4U+pTqZU
G0nirGjVh0laK6zt3B3G/P+CyCrSV3Oncytq3xWaHZAF8lUBgAok63lTYR5yZWiuNiQEP92CsUE6
IqLpTZipFhNT6rb0u1OLYUdPoEO+OoHdT5GMw3hOmvjvQSH31r1SK+bWObSxK/52buxIL43fF9/l
nPMKyQg/MibQr6aTbDzWZ1ccmjEoDds3Wlll2FE18zP6bpYUzir1j8IAu8KKGyZbbDUYFg0+XLeE
Dwi8gsK0sQ+Suwr05QLFi3IdIAQWHKuYaSF6qQlEv8xMCvL/cW8MlPD3yjWd8OqqwFqD4LidB1uS
QNGIKsmd4oCzbKKxDkL6lRzhHvesSEOsHF8MbYCVfxBf7B08PF+e+a0P3AjlH8b8VKdOf2sabhvR
DvUY2cZLqjg77rmvCUYN/HEvRq2U0B4DCQFRik/bDeg8LmfqzcDTYUbQoAz7pV7uEeBF6mYqm3sr
fne/X+eDq2PC0liTgYL1/CadrjBOQ1r3qKyLQ+2WBy18IGmY1CzpUj803ZClh2IM+WSi4zDET/z6
+/jFD5+N/6jvsoZLAKGrYTYQj1eJakrLBM4YCC7Gxm8YD0PeUTmcJBS7L/zQuWNe+JFxzAajw2nD
xOpXF+cb+sMpJj2saUOAztOjxm6AkEhoUmZMPoPHtuTW3o2KqZm46NJg6cV2VXZz6juP80pk2jph
b46i8L7dBq7ufuscGCm+XHQrLmRn+XQNOMZRo5A0JZbUqm69cDJHZ5y8uz5snIoInWxk0h2+vOxR
Q75b6kdqFZV5XwZTgKPWVcml9Rz2+pjUyHryIJFHFSIKTF7i171C4nrutMUtRwz48npoIZ0SAUkY
VBPnhChsMtDS3FmhXDDS15w/GiViWfvRnf237PJ8XgRAEyjwlcvjz1j6eES+oirNezyJMr1aHe8V
j+CyKDp/LZfcThdwDMkuiJ/9zjuMa9HdRNNAU6Zg0xIlK21vu9w2nwcJx8PI2rOhLoXROdxfHRs5
NucPn3K+JRsKSXOsYL0LtX9dXqTAgugXrMb7nJkvCV7r9SXScYZin0Gnz89bntDYfMvCniZ4GS54
j/umsghEHz27qDckYQcgd8gL6C8LK6rCFOXMIkbzbds8dunp3G4F4YLV+yr6I0XNy55CvXdPYMDy
ZzsAUqEwnjbWO+j6v9Un3Qg/LV+vtNaC8DHYR8c6pm0jOEnnpspgXs5W3GaJN8kSFOFfou8TigKO
XwPbTKqokpbrMrqOSfX5JoHFEC7xey5T2gBZX+Yr4ODd9oGxOH2Ayn7FgoV70e3Uw30E882X0Zc+
SAbyUeM2xwkPV4ofrkuSovzefwCBTQqM9pwGv/aTOwQdPvAlLtiRBzYowpbLSCWRSuLlw+KSwOrg
X7z+GUM2743KFkBUcFQOJ3Ynw2KuUwxuswp05Mz8AKb5zz+Jrq9TNM3yqpKCeIF0FFq0UzWxgtCu
NVDbPhnEwdiAzC0NURIChrJ8PxP4lh2CtE+vtJ0Da+NAWdjM8EQQBzEdxmp1fveTjmjYNA9vWeU4
JyAYsEc3HrNGR19WYHdbk/Ynjg9hsU/0aEKirvksLHeuLloLJMlMAZCS1lvLoPUyJHpq2uTIxJRa
tdmAEoBlOhjh4vnrh3TQhzBjrU5uJRhKKtD4f4Z3uZegUjLnzRcRgO4Nk20iQt6ktNa1D6FjzNsO
eoDCgZl0JMs1p3zhuJCSTtWwvGVUdwwihz1uofn245vnHjKVjnrQ9m7CtmY21hadzWfTi4B6XxWP
7DOTCcpR8/iugDvGRr89cA0prELaYDN0HlfKnLYFAeMc7atr9isaxaTRxlDyAYErPQYNnjJUzBhf
mmf6xIyqvLEQc8+ptumiteyRChLU/wjt1CWKEtjdh7SoTKIhCxw7sXKe7EGS42HFVH6DO2N3eLJs
hKeURmKPcktUZLAnAxNE8HXxUUXhdcAx1QLi9hsSrJ314anzy+6DtvL/SWP37CyD+2WI3AJ1XB7v
EoeI4eXRijAotMVpQ/yrIFlZUCpgs+FzR9TBDEG4mqeyykyYrmK5/2bP6rxUMX+/EGU/QiRA6V2q
wDBvcwYMMRok8N1ovbgUQlPVVyZzescWL39PpbOdhhJpiVUNi326jLXVWW2oG+TI9iNZ+I0Vb+83
eLZxWcIC5uar1JhOXoUOt8Wmr8DEkRPZpw3UtSXrcZv/9C6ECvMsmkzFmBtAergKysssXtNv9jsK
lf5sgZnWaHojQYg7QOrV/zt69eAQEMSK4a+M+B2au9jmLeUxXmwXlpgfGXSPSv4BA/lA+73Oo4Fz
EN0g6t0fbMpzhTJAkg8FScdbzWhbWPOBQvPxoA4ZNyEF+qzyrIXon/Gtb98qpwm5UTtyGkXxLE7h
wPcFXXqxQLfpfa4pr0JdsBx5IMcz6S2bVuFIIDQtBPPuLyTeh3Bi80iKtih03oQG+U5I+F7hkPm3
RJ8ghFk3nmDeAaXX107nk4eKX9Tt553YUR2dWPJVDy7JahMkjTyCfGUF9+ixBRzqG29IEEYJj1E0
dcII0zyMYyoyLDqGoPY64mHUQGs7AKtK6EYEHjUzVbVWdL6bBA59UlFflgFOqCJ0pNt44cJRiZz6
MzuZmZaZ3NwqZGY5YvhpSJQNZZhrkjWt/iR3maRIvC/A2xY/AAJ09he9h5keHADx4KyvKMpBRSNR
AgcdIuP6bM/jtI1wRZ8uPMG2yAZx4DFLwb2amhpPZ4bBiBWU24ywuBIrFgFxhY3gcNxVdSz3CVQK
6fvWbbOPIGsm6AA6jzQirgWZnuhwZiGnrhc962PZJBQbp/VChBWG11YsbKDttQMZcaZAnjF87b6X
+iumb9qZxoXWjafkp/lGmQyUl2Y6c9V9IrqPAdTAdLZM95tIwm0kjcE7tzVLYUBJX+DxQixW0Dg2
Ffwf2JJ50FQp0HTSfQ8ApF+4/tEV/T8JxjN4iJoAQrruKby0pQhQ9IZ0E5v3V3Kc/9vNgoXo4tob
1FNE+TBVH20JaKS3lZ6GwzbzEo9dKAgBzBVElaN6OTacWSeICU/M44p9gtsA/Rgyo8rYJy5BN2IV
W/qLpKFEWi2qiekiEjSgkUp21FKHc4J24kRPz4l4aVLvXwZUNfcy0ToT4axHJCY4LGaig5Y5zbVP
GBY/Qn41nrQZM68uiDxEgIX0jbO9Lm9tNSzB+CI4vhAYl7pnwGEQ3aCuJ6BnfiSmspmyluriel+p
4p9EYTN5bkUI5Bm1Xn111M3mQn8rhNjR5ZbKwXzmZbApoS6VI3zHvkEUjJtcqAjOZtARpHAxPB9W
M7ln9zuoxAjlKfTN+gi/wHzdTYiA9QFnY1XeqkeoU4UJEkR8t43ziqOv/U18aS0MUSW/ba4as1vc
/k28PIFtDMf67UoHoW4qMw3phUAMma7+qn/vJakgBDWEf0T44YGidDBcjAghVQS+KG/vwNA29Tk5
sTuJiz5aTiH4MaEnUXNq6D07PBWwaeuMUXF+U2x3bU3k02A6lDsZNOlO2WiIo2JRy4Z/uoGn5gAB
Ma50gb2qNkjwmiuNRBXSZ5zVcYohZosyYWUtexXP+NXmR84TWE6b1GDF89F04aFB/6PSmOcYkk3d
HiXDY2lHwLy1/Z4etpMvy34Xpt2mDkXIzAfxcjJLrU3aoyfmLKKQGKWxusnDLpdo3frZuo/aPyKg
9I9QO48xJPs5s6kOaxLMsqEtUBoc1t3dRhpKj+swY4PibFs1403ZmFsEH42xYWI/1VYOUBDBtOC9
zKBcru538r43R3KtuixhidmnVZOcXK72ed2oopxyPpbhmoXx/cjgIwh5OiwESyVvYCnEt5xNdN45
ZEBpiOle11K8yVyfOR7IgUe3496zgdE5cf18aaTlcTBBeP0YueGZxPdccUhgJrnZIPVquMhuCNq2
AxMep8oFZl2fv9meeu36vgqajKAHLvPHxk/ffkGI6T91pX+qvJO8UXIQLz8xIlx76TY/6ZMWn8UK
1Et8v3J7LDR9t5ApLhqCp+lCHfi27cvAZh9tr6I50sL6DyuzImkeRJfk/Kk/AL3l/AQLdsxzJIDs
WwFlngDb2Wk2UgW17zO8UEzcagaSbKFGPjgl1UzWzNAMy7Cw+WLaQt8pLZlDv49OMUS1DB31Btkf
a3IY+gNjEiTt1Tu3gF7O8iMywRGpsZsi6z5m9wqKED7JtaNApuqZ+9ckjxS4gy/SLXYWzUv7qqPV
mjS5fx1LQ439/hY+rc4FZzHtzKrN08cRwNZ2xbVmDGS2fb1vCCFrEZfaJUYoz+Th7jlpO/OEpXU1
wR5xH6aBlIJClwVMjYQb2pyTGRvgF1Z8VXeRWx+7UpWF5lHTv9KopL3Y1Htk2BgvLPQQm+v4hAxK
9or8Gyg1vSVhDNgDApyRYphx0h9CpoR7zNC/K0Vur0FLZvD9Y4wd8iFs2KI4cuSmRyDguYxNoeLE
nVvEr3FCbfb2XsXZ4hQsuSCJcaZkAgJ//j1T9S2F9qY90T83uL8JHdfp2HZDnMmRZkW933NQaXg/
1cU2JcfjIRDbymN4eKDBALlQIQfGtke9KtqSEI6RAubgmFaAiE8g1ElaQCDSr2RCOEhuwqeUOdXm
a7LlCF4u7q0uc8oNtN6/6Cxe3MySUReFTnThaOPgdCTntfDXhg1Ne8znHGu0XW0fk1RyLDL8uUzE
mNaQX5th0Lk3pPfHXrQ3Sp6qvKeQud7aOAGmTeFqeRc8OpVRV8fOZa2dXIK7LAIU2QZU6qlWTGBp
4XV99GGFf3PAYxD6Ifxkvq7Y16Z6oTIgV2WjzvXZEvEXeXquBM09lgPSKDlOQCh/etaKAxlaiBS+
XT7tuVTFD4KkxIvj6QOEj0PUqzUSZXb9Vqxx1Gv6mhMtUyx5iQzEavvTyP0bEY5Qi4Yv4ueIajLq
7oSCATOq8ql+klnG6YX2xpYDYXcz8KPkqqOIhX+55gykZZFTuSAgUOhFa7euMiEu0/b5EE3SVA4C
Els4NsoxsoMKhExAnzKBEn1UdB84ETNPRsXO4MRErqVB0msen2qeH6t0H0C4wSdkwUkBKYYtMMwb
iSB7XWawZbRS17AC2LmC/MBppmkq3T52esvFe6PZFa6qGvcs8KLL7X0R0QHncu3hQPnxwP+ZRClp
ctxj0wAWzrcG7gN7YlNue6fwzrJKLbI1XNKCxIj42kZLUAvZzXbArL5JOiH/4QadVaH6wwTDktjR
1CpRZZgxYMbM6HQBl0IUrrs8inJ2M8g3keML05kG4jTNmTsfry/iwqP3vUBTMcwbSZlpuQ814oHS
+TgqdRhaD2DSJxTagasa1OavZ3kQz98VaUqKm1Gv/1ASq7OqVVMsvaam08wt/vUZmqXeNlrcI2tK
U7j2Mdr1+QjMSysxVPVIxEMPE8Ji4NPXSItAkm+bTAAUeInNjE5u6xZCMTPZJ1swkxw4eCtpceU4
8l3bylbwFEVZPWxsSpvC1l8wAu7ATT30YskXxRNUWP5llD9elZx+SZW4Gsvxs4lA6THt+v98CVKc
o2dUrZbgh7M04mKz9hwCz81GkdhzgpDzX3T/etoZgvd5OZA3XuMCv1n4nTHe8jXdEVwGMKehq8uf
G3dDT+t9Kwm5CA5IQu+eFP2/NVFDI7VLiSQ7+87dWG0r+6gu+PSBIeyPMTZ4ow6Y6/E4inI0BGIE
P/RRZSYrE/oHcxjt8xD5SELgzZusneBiL6E+fE3HZ3aLeBiREQiNoW2USaNKfJ9BZjW6byuzp6fG
77DlbrIUkm/nRGJBoA5vIUCJThCtpCIipE9Vsi/65reZF+YS+/OsLt2QtcJ63Apg9qrG2ZkrJLLq
LBXAegUr6LCgcBHT7t+WgA54kNhXW3pjDPsBFDWmxP1RYd9MmwN1sqCFwHMjNgeTLjUDPNLq+tqI
6WduipXwL83773QJ+NHLB7eHy++lprbD7GdlxQiTuoE8B7lmGNpDZ/DMQHh4s2u4ygf/oD6w8Iab
rDFAkFMInWcEEMLG0YhTc2pF8VIDk8cpdqn0anCA2BbwOe7OfRnKcsxsjUA/m1a5os+PE7L8nJcd
wOUI9tlZXP2y3afvyswRaHDpDeISmGYoWvhxsMIAiNQeNk2LgeJ2+SWl28iyWVRFiQLG/aflTtzH
otInDOwauPhB13mcwrom8VM3SCJ/orzWsexfDha+gPI7lKOqwI+IxEkpF4ko6twib2DI3/RMKJO9
QR3WQFDqia+aiONpJmHvthGr/KJugAZBJ1GQqrglgflkXKto8tmUEXYYCwUp8H8tvOzNqY/lZuFp
uUU86GSPqk9R4t0/PSBCipleNu5Bwj081GOc0MVCcxTBVvC0aRZoregS+lq5T+i/7hPAC4XIZo03
RM8yrLVbAbfztanDTLZRijuQfhIkKqgfk8U9SiP6zhS/WBvPGqadPfbHa3T7gjztaIXBitwN3Ve0
szCFskzJRsPKmlJoHazUp9HDsq37Ye6B3Zsx+a8dDKF5e2+jpJZu+8iz5fOGDSnCONBGe3JrmWOD
TiFin79VIWiGIBwwf1enuZs+RmwEEeHBifzj4KKTfH5hTx+T+d4V2iuqlrNbWSrbVjhGkfGadFES
+kXL0BDH1+J96Bly6SSsykMMXYfDwIAXMxtTZNTZDf7N0Qv2H1Ymu5ZDlNgVpt9zmRobXYK3giyr
qL7TlQP/ijWvPPNrtSe313UJApyxnzTkzeZ+rZfXlY+dnz+uaXALlLHA3d0d7VaFOlbEEPWv36JT
4gXaBasw8nrd5yysu+F5QQb/z1q/0DWvzpWg9DpsWNvJKjDQzM/t/8NPRce3XLjcj4FxXw4Dk8CH
7xPdAM8AgXT6V7ESDRsYs6Y2vbdWl8uq0Z08cCUvZJKheJ5nGD6JdeQPIMB+dS1CJFXdGCFG/sNg
iWs03bo9+eWHP8Brw/S/DymMiSRaMAsjYilG9GJsKHHwavjRFXxs/shmfmc+y2Z0ebDwgfo7YdMR
c6t/KSA9f3i/1vzAf5S5jRpCkt/etYOYoNJarUvblrYYwJUzfubwzBzMRUfCC/L4AV9WYvOU0W/0
dOz3gq6gNruB6/3TfgZV/cfTrKk2NLVU/ojsWClIkr4WKatlj7JnTd+XvLomIarpZ3P0fvVYDVnL
86XMmFpYAgWTnFCVM5u47rEufdAc+WLyAkU8dA+n0LLBOAynRQkyEcdNZxzCqvNRJ7k5ZcbmvLn/
oZm00hEUgNLaN2PcPfU1p8Yv1wM911byrMC3+Bcl2qVjePYU7qnR07JsW/+V4KmXbC+lrXreMdwm
7OWCJ4pZGM7KPcs16xSZoBDGOUmzrar603zk9ZTbhsNaOghr+rtHFDFlyaqleONicuXldBllBQyL
sJFOZY2AZqChq8NI1HxyWQVgCiH2qjySijcQDYsc09ww6hwTwO37ajzfftb9OEMGhfkAInM41puU
N2/13CPseuD76TKSjKHY9lY5Ttb7OnyuDnicVFqb8XZG9B0wpK46V42n3OfyQsS7g/Mn6WHFo8Hc
y1GpZZOpf6ONVvWGnpr9FPyrlGNtY+4TBM8B16CKqdsZ0Bt6PzJwUIMo6ijNvR7BSanBqkxVq3PP
lrgBUX4Y/0M7hgEr21hqMhyJzAcYg8XOK8PUanrC4ZdNTUU0tIqIkkiDGlh94odCcoC1TBtFA09p
/YmHek8n8i45u8uIKj17GnS+ZsdOfQUUplvOcX2SZy5mqBSTDizRYBLrdAMzJXCuOZqUBOpFVGom
UqgzbtPYrjE/F4kEL85Zx/QJUNBaMJwHSqtHlk5zWTGxUa4zuIEC6WP4wszJq7nrupDZjffreUdd
vGAWKRG2MP9QD6RokVftyzNj7tqICqLjPqlTQe2Fvc4DQUke+bMx9xEHx3YbuwZlaIFiBgMLdyT9
pyf87Ml+sz9nwWzqVAQDhKyYOmRjeGn0zKeegtxpd8p6GTuofYh8Uf0FkgJ+Ae9ZWsnaoaZFgdti
+6ymyQm5ugc4YjtX1aV5XKv8Huq+OQ4t2DMbxivTaZFkKl2FTHGL9PwTu08HhJapUHKXF0jVNBLL
mQbV3KQb0aHGhxPapyBT6jwjW4q8V52IayQPxsO7g4ADZ8px3JgZf4huA/pbT2mn5pL8TXLpepG7
xcn6odAeDjB1fwxti1vE5GG1BgUVzq63gHV44EHdYWbhYPEtA6CE7Cfv4n10+dCwRJychKeEcZJz
QQu5rjDvFl5Q/Z8Wk9/D+jQRUaOyCH4oH+sFu5FVwQXebI9euFqs37ueEIlNXK8NqZs0oOeWV4ru
nShqu5p7Do2ljsaTmOi/XbZESvJeyrAQ08slBQ66PLUzwYuSHWisia28TZb4o2rroEtyp1lLg2aD
HmMMNfEAxwfyDJcRxdmCEAzvLQyCuQM0o4bhihqo9Kt2cOuHFxCq5ECwybt4Lv/WVUr3KP0t97NU
qBwVWicKiVzJizEoh5/9CGTcN5dUSYrlWYBcO5UfUZ/tZKwjrlyFPqPWWma80tGfb3oTGqyeAw+3
7PjRCgHFQkPF/VHSqRVhQyHH65chlj3UwG3Y5NGInLOVbA2YhnkTMq0zvQF+fGkwwe5ZpiiSF+ZK
nijvXMJkkv5ALJobMcc/jMXI5dxZoBPyZ5B+3z1CT30w4U4ygew3u3gKFek7s5yeSOd2gje4IxvC
mjIeRISv8w0YRDJoTqOlxeE/lZYyeOUZEADL2fmc24dDayZmywUHuYyPXYlUeQBl8l0kdq0r8YGr
fCJorEmB8yvfJVm893ROEloOoDS2QvuG8f7Fp8R/UmNSgC5LOychi9unWoC0b+xOJ9IMgMyTPXCM
3wbQaMZKYl8YtMyExR7sIpG1TkZdCfKPLF1gWPHQE9TIfJUaQ6yshusdU9NyDlmbArMn3v0xmbnK
vBzgKoEilLo6DwYpV0Ugx4yKdlUGCp2bsQV8DagY/3xcMPHExYH9uULzJMB+YelS5/xiCL2o0NaN
wExGGKiQj4n3XXziXjBIpyTt2oGFKs1gDtsWdCZ9kEPEHfsNSmBUJFrpFWR49oBE0sKzuOVepT5O
Nz+gE419MgGDX5dOCZ7PB61QeecAEiiE5tv+ZoKLawCb/nvsX0l/qZB2WrOs+1YeJSvXBrG8qyPk
9/fBZK5utxgF+SYf/m56d4fdhMcxODwrmn+2xEef0wR6Kkt6YtNO5Pqw8YvFovdYMRGxPWgudbi7
K07VRvpm8OKEofJyGHD8srnJec/81bBLB1nAhWV+Zh8ikY/1pLhC6TAtW1480+nDbW+o2Z0+my0k
Bp8Ke2flL77WHF580auSle839fFtCajId8xyQYygWdbEpAyIiSCyfRq4e8GUbX+wGNbWr//1aS3E
DSVmLefyVrE2B/EmuEqdBPQ2sMBOouoa4t3IE64RXd5iI8SPlTEVdWwiMeeq+HR89kVi8TPDrpY6
hfLXW7+0ZKxTniaKW+DBcP/qLZfbc3hJu575JzUNusTOknVmk74L7P7FGVRT7YRxqbTcuiPC8eaC
K92mh36qlS5LCDWVo0/Tw36e2X5IA81B1WN9MI6dFzztJJfdiSsgrvdupEa2EuU5kA/BNQuLAiyL
hkqFCTsjK0fKcf4AZGX3e3nI2LHHgKupP5fYnaFVtfVehvJ0Uy3DLh3FEWuPHzi/J3A6B/dKPnKg
DV4AQqnIjNFiLCRNfnByt/QF9Fc7IjBCfRVvE38xPi5U10HSt8doWFDemEVF0Vg03GsfQH7sLe6r
IllyPDKwDvfA3NN2n+GOvFBTsr9dvkH78GvKDV+CIUIbriOQg3vQQpH44TmUJFZT7pO/kgwImY5D
TQBHzQkiFOm50IgfcizDlYVUDyq5KW+a9h2uH2t/9GHmD0EBXmVwB9Ps4l8ll6IcYB/b2BvryttO
eGaXdRQvAJeX9hBhpQDRldOTiGU2DHzwx7qKWG0yazpFH4P2Xx41B9e1JK7+j5uBw1QR4eiKaZNX
gLfXmsJwpQk3ETMQD+dFaFDi0c9Gsqaa3v/vqoZ+xbI2Nr1Sf0RdoE865przv0M2hh59r58CMwa7
1M9bnCHVTMPBH3UNJCoO0FhT1MPOlDsyZH6nfdADBds+LWbZ5FmwaC9Pv98ch2LzqzqnaS6R7B3d
5ZfXRu7rYYJJ+wqkL1cPl3P6nJ0qZ1Z/xULPpArGAE2VhAtpp1xWFfJ7UJ+Xa3FAjrKGNyZe6Fnn
z6Mc1MDYWglLNL3kwR/OVHDmCX4OgIKxKVLyrHpDU/asOyQ66gH0qK0X2LAuzgI4Fs3wcvhXCY0L
Xdx33PV5TP+LwLMKXIGHDt75Ur4UcYCh7tTB5eT80L6wnJ7A4OEV6BqiCPWkpHGz7WpzKjOwtjUg
R1j8CsgcJmZ2WR/EesV6KD2SFqIB0O9ZJpUbEffqo45HXo+ABzMi4n/DZ53OIBSQgilgIkj2qM4N
PfG59i0r++B87CGWfPBW/YWO6QMlWZSQpeJiLZkSKeikd84+dNdFtSybxXfglWPTGttDNBWhr9NT
R1Y9Yg456VV3qeHLGXppwp9osbPE87cz/F/cUm9+pouVjql3kMM3U7cnFH/ZZWS9VayHc0lGZwOs
kYe2uW0cfa58UVqMaquZtBbrpAEsYe86xiA3uFEjUHoGcwlhitjc5yRDWUAL0Bn/VAr7oFXGEvvK
CnV7GHB8XTWvF//+ZxNGdnNXuSvVSg545RGzClou5HbE5F1L6LyKDCIqCUQd7zoF6/xizy8hNEtF
ww03im0bxI+FjgI+2XeUTlq9rubV8TxL6UbLJWYm5VclbEgbCMXw2Hhn3ed1TqCDn+pDXneg4ZiZ
sgsjh8f6R/VkQmHrt/wTaZ6wbqU8dqGa4rZOcqG01C9OMT59le4c8TPd2i9KZ1yH2DaaSpUhnr9f
VzMjZN6bbUA9EkRapVEaQnPg4sDVQWfx7nuxEKPkmzDZ5sqNPOrs0JeJILR2q2IFym9jWr05KUkr
Un0ZdGncZq/rE3UArrtHCGya9CkEII0zjFIfh/oIupt/Zpwz2S4/OCffI7vulM2aCQGUPFCQRGRe
zqRQF8dKW4xPFDGoWOq8N/9V/qhREUz/tsIPGoYkRqJ6gajRIw6L1tRZ15JUPJ3n3lF0ZLq5Ct6f
Eg0qjrsCLeVjKrdcEpJCYEN0vGWce2tMrcIjHjByLHMKaXAkP0KffBf318paeFDpfaMLgHeUcEzP
eo42El/3TC9SpqqfhYT32bjgy0O5ZyblzQYOYfGgBeoJjkcQt/wdhXo06dmucEw+Px+dvG4IVAiR
p+tsw/1u698IUM8Jwlep3jHBT0eQpsGYSdVjzBDwJ3Iq9JcnRm7uGgSzZDCoHsWkMXTxxEip42g8
JNqwkIh6wJq/3enmiPpTwx+v9rtSSJLau7gRdF9vauYcoxoe1Ij4Rj8Rny70fL3iYyIWcDCO2s2j
hW0ChbMa9q6lzfoEIlbkTQni/Y98wfIFpzlCxZ4Ge2W3nUO9v3PqWndJw/iZh4zrYlAHIk/rA6LJ
u+zRppNHLAAFibU9+tHHUoUG6gDkbyQZ2PZQGc7PvzOkmmxoJV28gCOiX1k6Bq6/UIrvj6rziPAI
7ch76hgfFDcT0ETVkZzZjpV/5+lAgVTBq3iiFBqPfi8EqnOixopSiUCj+RLvrHfuPbNaigyi6jd1
lhRFGalV2l0laTG+x0V68ABESVBGUmId1opah4LjWCYVDiI/mZGQRde07foFi/cXxpZ9t1oPQvCz
wuzS/h0CTjEkjk+r/xzBJ01nI2kTqVBBGr+vd9DZF90BWlzBzRhNgvBEW9Qd3pyIC4Lv2YHq4tQQ
RkwdHz8lWaekFR8fyhEGxDBXRvSOBD+veSS1CvE+MfPWC/h6GQFqNZ+sEIcelrRCLpHZCdbD5av0
oQ3U/m1391zcW0GdGqNPC39a1ideu13Yp3BsTiNrxcriWHmyQzxDnwzNrdnOV3hk1THxcdkWFOwa
M8K7jqpYCffSQRFWtvYp6/1flXWYzXDenzq/kcjRAmJcmSBd4YkjhEPG/txGYTnKYPoC0jeaGpO0
nbZknDENVvkXadqcCGHl2zNhxlynPRdR3Gq7WwV/NvL6iF49VeWF6qXOTvnjuuosY/2CFSYugyb7
iYoysJiWqznkSH20xaUO3z7f5R71wpJ1qGRGit/MvcocPWgkq/RZqkOC/CcCI612x37Bd53ULrHm
pPhOf9p62DGRe7lYhxSv9r4bT6qZDZLDKaQ883m7Hz1J9ppC9YHSHCi+ahimPqGLD1m7LZTio9vK
89V4NSV5Y2fTtDfL+U17wspcoHk6t+PPzpfr7SphOlYg3t3IRwH2YAlhfWoO9laAv/6aN7K1sSah
P42sqheFHCPYJi+6uhkSi2zd2EcFKp3RkXjV/Q/2g9B0Coi/tvPubvZ4fYc8WYUKl0YsptkEdPkj
GcJNnZgOBQn93tPmCfgfl8Gx9paasE61BMOGEn/yJa0HYk3bzd0luRN5fVnHq/N72RJtp4ZX3wBu
FFdKu6e6psp6lETznwV0ctXu/TZNsSTwa7M1ddXRycDOYAGIqRGsIhfOJYszuQPzmgs76O9Nz4sn
/4tA8VOGp227HH6i3WZKN9BcFxZW++M8eV1g6xaKrzGy7LFN20FFVh0EzQMhTG92xZhx/M4M5BzJ
M9I8hEwLbf4GtxFYfMkaFe15s2l7C97sPaFSR1po6MNWTokT5L58e4PpJxA4TGgk063rWMlCHDnl
k0vfpI1aguhT0haIKq29vsSyADcJ0qOG8ti2V+VAjuV8gMQFc9eheYLwbMN7ByCeW8n6PH+fmZPJ
+oQ3KRzGoapx26WzHjloXB5bTH837GVSWO7akUeeErupwSUCX3888rLFrRU4BwLul0w+FfATZeIn
xtYu9tom7vQP6SFYqx+efeP50QwZE24SpjG5tlsvL3paXyR83Xfg3Xa+gNrrKwQrBiMt4NTO6zwB
uwCGWIjPYWqck0Fb3X6hq+O9yPgE87uPlxFKvkzfb5EPN43hYTjoMVeaeo2zOVFA/diIZKpjrlHK
2BDrDI2ZZVEj2Yw01YvExy6HvxRvN/JX3AhmhkM51TnIugTHELSK/3NHePw8x0FjllwCufQUrREi
zQL3pkwOoCGZcrNHYmAsHueChg/DIx49+l8/5M13OKhPlFsZZYbmibVLYFsbmLjuOOHBx+6Ka+1t
U+pITfr9+pecIDR4/icBKgmu6SlGnqVEgPu0KlAS2D0ZUdsoXl9nGWpBSZSYUEXnj1q9SejbK4LD
1DX7H9acFEY/uKL5/7W/EX9S/MQhly/cosThWgVj7mHv1QQOKELmxeGn4ddsCeVvDaSatUqIbXur
DLmldXZF/nNtYE4QVFjoLpfmdls+iDDftnemyUP4YaeueFZOdNBp38DEM8R2Es/6UOztSXxE5V0T
2ilGjRYjZ3ItNievhx61K3fdGUo4stqHjKuwM1Lk8B3oVxib1RfQyClPos41blDykKXa/kqqcNOb
criwfL5wUvuMZYtNsCJN2mToMqvSsdiZzTwnm/8CXcMislTmZ9cPSGu86EZTldT+uDrNFge8xB0c
dB9SjjlCuiQkjAQpwI9kPvqXpH7ns8L83mADFWPyZfnX7QAq3q482SvRHmmHJCRvTUVmlUKI+Qjq
R2GrWgkv9ioZSa4SWJGHiHycACoBoc3znJ6tCxotniS+8btQjwcXjbPsqVYYw6WYWF+Qv/dqOy1b
Fby9G3N6Hi4qYdlaEOQpTnZf2LoMe7BBYzpSzH5FGcPIVRkCGNy3VWVCwZ9Eo42SdDCdpB8FkQbZ
Updm4XuU+Ly56WLjpGJu948cbnkVej0usLTcUCx77rLblhfXKkhQY3Mb5V4kwE0oIiDaKyIWEVom
G6EujucCXPALsXNXfvWr3lYTa3nM28YN7c+AdZxzPl1t0H4mAJJUXfj8JU6lXzWueP5hsvO48WcW
aZS333SNB3AboEN5wCXJh5TD9TV9xaYCsid22vrCkKvGzOMyv4KvAh0aDWsqykY9qxyqomvv+2pP
1ymZTUxu7DuAvFeQat2+vClBZOYODTV/nbkY+8yx9UDjA6EzJz6T3dBj3RjnmV08lwgQtOtZDpla
P1sGKL35cgsiyxtRvRYgDueZgo4Enf+XT40UDSzCQGziVa8N0olm8VGO9LFtv5WVTUqJcQwR6CXg
2SnJG/t5PsvCzBLhy0Qd1Sgvtbp1/zKw4W+nRioeFK9QTzpDgQGV56r9M2Fi+NEw2uy3USVZVgqy
3wRAkc85Tel9NAEcvhefbFD7oUubdz7e8LPy4z4Z+0XKHo7y28zpGGX79uwLLx4JgZe2OBhnZWTT
qFVq7LaAMezajaYudE3MF7p5tyRDqwufPIU2oMAW1KgaL3XsP28gKBdTwLHa4hIPfcIdm4OWzuy8
NP3RyoPY5L5gagzi7dyMx9Qj+K4CA/bp6H1hzmuIr74bX7idg+9fVcJdof5o9BYB8oxH7QkErmcm
mWALeKOpG1Q1Yemd2T/OimS9xu9X+sfRQpS+2LhnIYBCWVZ43ZMpujerjUvokh+5FSH7fGLnKWU1
ucEiteWcPbPmkLhS5+UDatWKS/yWbGaAns3hjiVTQ1hW88mFgTbo0YjwSPBZ1TKz8dUtrENqffpL
0a8QM+jeGEo6Z0RD+/zBzkxZZCkbMsq4YcXOv2D74wUyMZV+Wy1wkYae3CnMegxB5nEEMCcpY8NY
jatYOQj2232RZhTPBpwVOTNwx318UH0r4dj8QV8skZ3wjCNFO3YCSg9VelKzDaS7yZk66dKkf15a
ldJBLm8TRq4fQ5INfNXLt7u5mz9xAbyEePpRL6SlXYyaAY5iQWGrf9VtI8vNOFebcY1Gnd+Gxmbp
IOA2+fsT4qtr6655vHHyLdh+0N9O50qsqPSNv+0HG5rcnX9YuB77XxctzlWTnaoJvBwSlvXJPRR1
Wv0TfXtq/7ZwH64S5lo4WPI6GDfXmgibhYFcUU7I8zTxZNokoctfPFvwAYtfMd7qYMtCX+onbpKd
3bYl9mwJ3/lLZh4JuGiskm+ykF2px9SNIsvNg5rP6TCE6Ad6YY8SmX1CXjLFrfika8SMWUnWbn87
mB5M3f/LJAamoBOYxS0gJkRYsbkimnxHUOOZt/cQlv2uRKHATHy2GSGfXADQmnEoZ4JC7vCvE4jk
Kl8eXmoLPf6nOGZ+Lfks5mNy+xMHWeL3IqoKllWsBskOxNGQsmqCybawTUeUiN9W41iPHW46Oi8F
ekM2QEqExm66PXXujxzTE5ESQFcvJRisYAHzF0d4VYf5pa7kNxy6sZNkj/9nDZZaK5tyrVZzSir9
OQSo5V4Vsrxyg2RFcn7/sUeiHAMZnQ74Sbatug+54UsuobbDNZo+sml0ikGvQa3dG9E1DCWhGNB6
0rxSwvkwI9OVA8eL/zOG8sSSmP/PiI7PY2nTcwkF+73mG9POY3ZKEkMc0cawKSh+HT7yaAcGPDao
D0IF+qfaKvv5LCX1E+mezCLTG1W8Ov27WT2Atc5+9jVJ1KUmgzrluFdb8bNRLR2ufscCPTjpk7PY
/CEc2/cPRu50sor3n6FRX4KpVVKIZRGFvA3wG7Xir2HrDo97uAfZdWHcufr/ROXx+1iwh1yWVglw
1QXYtcf26aD81Qy1xTUzdYazsnA0wJfOhIiazOCvyZYLds2Me/lNVkzAJhfrxts4EfTCsHkMFtFr
YUyNlr5v8ebta2HzlMeliQUfJ4BhkMAJdT9VnApjCgpNKMCc58Aod4+3ZO/XDzwh0QJqX7T/wAQw
VhnVRoMNxHVKyQpyzrcMKnf3Ttghjr4Mdwu5l56DlVdPytUqpQ1KlGZxyoSmdqyTX159dy9BcSiv
g5oUkz9L2zS0o5gUyMV5Vm3wxS5oEdJC9S0L5189P1edv0OG5krxTx6hZ4xakDSF9e2cNw3oiGCt
f5xIc43GzAB6nW/YtK+2VIUO8kyerqAnRLpwkFyB4J+aIeP8BYVivFYrGdj3ABtWob4SebZt0bD9
XL+FLz19zUb0Xpreh2K2mHsxSPo+bpmmgvFKCtuRpIspLSd8rOEQZhNFCpQ2PmE201JE6cbPmAxV
V6hx6cx7RE+iOWp216OnkoCV4PN90JJs6n/5unGj2bci3QIY9bJshOOsQL0Jlzb4BMJ9HGVzEn6R
xYIT+Z67pHPu0f+4k6K1+yNm6CuYvPoxlStLVvKD1sXue9tRUxARwDY/dZoYGqA/k3rpQQ7JW9Db
2i4zu3Pj810soIhqQW2aU72Q3GC3NO9aNRPN+qnkuuNH7GmC7ahzp/gvF7e1WSa6IuPIDPKAc0mJ
IAKUWXWxbKbKdURS9rJFadNBIDxB9DELqZ7bU9utwwD0i5A+2eUW2fVW7lcID1Fat+LdJA9noeQn
72Wo2twiuLveyZ4mGn4YH/pnBUyeuuXmwtJ/2DgPekDVFIoPdBGByr26IYcCSogYbdbhiZnH+9iF
2ALYDu7f3rtVChO9uqgjJQLL30uFn3m32agdhX4iL5ivZb26aREwbrhlNWSSPsC4no5mBVARnAqF
gnKV+undaRXl+mfi91tbQOAURYrDILRTr07ArUwL5ZiSc2y1Wgb27jTSnXwqMhxsHJjT672zviU3
NTUkKzULCDmPsEHdIzYhyIwAQCo7qWbSYUnV5PKSLCB12EHloGawq4+GxVx8vjWYfgBrzN9VVbzU
i2jUeGHxWp+oY8Pxk/6aQaZzQR2s+DRDISswTiYzfkgsZnnn5HxiE/hTmOOMn67sWCJ5zyQQnzXS
deNlhsccl0Fu/FjRS/JGkIT7bDLI4tk60B/Qj8itK/1/lCalCvPK5qZek+W+pc+Zqk4HJbx6Uh2K
uqEUgc+Rh1P+fh52JsKusOH2fajcKLNPc2YPNe5VDE9S+mKgn2lWC6aM1Uvho9IdMATfEJmO94Tw
jw0FMMWDop6POQmQ5XGWgTCoKwFKrbaOG+WE98LuY4ujyacW6NmzzAXPywg1p0k4pCBvgMElqcib
6+Jqn/ADWMFY6hrQiAbDT6fCVtDZtmDHIoT/oOdNzNMtxr/C0WRdoycJZBH3sDKgzyMOs4S0L8rz
Z/+X5ZIvmpthBHdY72qFWfBAScEq2I2n6YM2pH3m69emnV1zNCgzSsdsgATRNx4XlmOT93IyCLuP
HqIsQ/jWwQgCH6OYbEzu45YDRbe2XwkKyyd0xRLFfiILECs2eK51FyhT3pwWpl+IPKVhpbxDcFin
FUqYSUuMtZZtgniM3Gz8/q2ddTyvzh5x7iryFTUKcLYN6OX3wpxVXNwZXa9e1fHc3HCVk9L7ksFB
9H7jRy50gCTctwLI0zajFk9tDyGoF9Mur5rEmKs7qZrzEYI+bVUxSSOnbgGNpnUtVHXQxV0gP/7t
RQFVcbtswTNtG7dl2v+ORozpmOMgwjntU2/Q7gyEUgvZuYaaUsns0SCf0jnJJJZrH2u9p+5MYXcT
R0qSD6yj+heGBewIODvxx2My5u78mvcg+OFkBsj7M4uFoKGwMfrMBnvkvTseJfTWrT5fgpjs4Twk
0Xeri2CurXUQv77R6D0tHqHP5GJyEUaW0cyYme/uLbTKj54tnesxXKlqFx85Fjd3Q9a1fodeyr+W
QVobl2/P5hU2LDWMewmDBFar/pjEixJy0ZYaXeCQ38DpdnS4GESTtefvt1/BhQETZGPBZOoAmp70
bLJ/A94xFD90Du4u9AJK5b4/nmSwou2a0CxuVrnI2XRaUxVmO2Cvfhtmykw4T0ovTatq5bhYElBU
Qj6Dic1zcCt9q/ulGMGtOySTzUEAvB+mTf6ZHcneXGuFiO9y1gYQ4DIugisZuDwVDiX/DiMca7Ak
qVun6T3B5ZBsLQ/7n5XV6QBdJJ8uQ/Es0B3z6vmOu6a6sEDXKkF+X4P7oqtujXYGWmSFZV8KfDSY
iWUGMmZDYEbWZOEYCJL2xbQda8Q3UHzuO2GyoczKn0hcfglPugvrWfViT2lWV88QkxRLZ3vIzdes
v848YD+N5mIDpbI21pOCEiatnQMrJiSW+BkE0VJl9v2wJa3LDgBcM5JXNgz5HRCCSudK7bsA5VEe
4xhJSmVTO22qTRJJP7gRS09EBfge0e0lvgXqf+2mMtGP3NKtetuiKgpRotRlqr8puEL0rga1qIMd
C6M28/dmMeyMvadF+2xppaom3pCLZIhT3hOugIMY0Cvu0O8DbrK6dGENK/9NWQSMpokaiZ7UX0Ix
IB5KGyoSJ0IeblfhtdQsrMJq3hGQBKbVIVRs+/2LbgKjPJSB/wBSRZoJYlIzY8I+2Fih+08uVtz5
7mW7Oz1ZFIwA4zsWpIWUrXqTkGejo9gp6WzmcPdempN5DLnC4c6nxeSas/ik03vn/BrwXZlq55Jm
xi93Wwy2GESB9clSlVmlxfE6KTzmAFq34DCPEAyy7FWqxuznh9CIePU4aXr3JEZwVoM1rM2f4v3r
4atp51ZlxcBneSDsAplh35v1bLEpx1gH62AFJT+Q5jxyCezllh2PjiwAt3lSKUcHNScU2u+Dk2+o
Vusssws/YGohBihzCOE6cwrVW1PyFN9mag7PgLjovop4pg8o9RMTApNoBjVGeGvFL2y8Gs8Mf8Ex
JKA5wPLUYniAXns5oPUUucWccqQtbT14wuSv4kTQf2xi43ZLJ0ryGeJJ0WFmXS4HXt9dfFjauytf
jdBUuKUTxC51V5H9etPyZrvYuhJyVT+f8+xOJUmnGPjJMN/gZBUbR5cVDQCuppBC17cNhzpg3rmC
vy4e4wGY+yBMAXuBT4xs0HUEQXjJLBGpQRSDeHvJySFobtTZ/zhxcnoz6yzB/9wMbs6NzOyclUuJ
vshP3+eaPXzHeW7D2I5/WyETb5IZXm2hmumxiz58AWZH/blQIvqwEYsJAJLp20u1ki2xZiCti01H
eM5mFNgNChMX2hWY8hn21b0oIg13CMM15fbR4ifwoirk7QzLf7/iwW1fQm37rmuftvDpAw/+lVKD
ijKa04F36vMiq1f/oiARtt8GtbI4cJQlVeQ+CvBspJOX+tn4d9UMK/NE97/Zk3kLYuKQe4QpG7n4
E9EVvinN4ee8b9WFhxSwSq11EY/RPmykVNzj8fHTB3z8ymR5KQ6ib7/GUUBqXxmXRes6vV3SNoo6
Qp87M8M3tdObweRBgfq7zpKrRqe69Mczbv4+uSbMtRfFgRZxNIogCPFrCavw4eDlMXSF1+a1UcM1
bz/pcg+kiuTVXdQdYoJzPb9JkbzO+gkdPkH03v3wXHYyOMYU+GLvSmqgPOxCMjRjCX0aM7jMYx7j
llIT5MavAHe/QgqsjyWCpbaKTohJpdVBYuBZDQHPf5oIaGly5Gx1+L9POIGEQmlYYf6Qlb0Rj6CS
h1mYv4YayGyIDrs5ddBW06Tp+Zw/ynRVAWvgh3Ju9nPEWu6IMUub+baNA5vEkGBxz9liowhfK4oC
qesJilIEu+PyLUXi0+NKbMz/eqHaSYCYb4sUrN0XODpErFNsWb4s4KscLUtkIdAHafqR5HkJysOE
GDM3iV9/wWvS0KoiUcULrzHGIjA7SqTC/pPi7Hy+07WKa8sCLnrq8e/6hJlkk7nOlR/zYxbCZ+Rd
jXtVJeCMlPKs4YmkrVISr4gzHv1iRjzm3ZgyX+We9Lbj6goeLjbE3TDsH/A23QBBJwIVRYcL8or0
QoRJ9Mbpeeg10CXYopBzTIBA5rzdGKy9GtY4D0nAHU37LGEDyHWDK6gJ8ZSMrvtINEPNAle/VjF6
CPAzkvjKG8gQc/GTwKxL6hn71M8/ed0ELJad5z/VCK4fb0UPnNrY5wOt9og9HqSXyoB1vdK88HY1
ZX+d3VKMoEhXl+VUAnw0+0DgCSELr0bBY5wcRjAVPRWMBiIwrKBYx88IA+bAoVfUDbVAY1GDaHX7
bc4ux+6lLHd8AzmAy9gXsWktEUPZPVvXndnpo4Sqsx6S33V3Ta0Lc1JQWufEiFX4oApyhlcFvCrg
TeZi9H39Hm3Fj7UJnS82wbCURsLdRCPfxjXzs0L+9o2jQX9nhw4rvdX/hA/D0bwRwDaHzu2E5raz
WlyzGhuBkPkEWcjJ+DcS/NYvyCwGqF0kmRLgdOaijB4+vIPSS6tAyLiwSyHwXTeDX7SI52Rw5Len
zSbO316ksWITj/drtJnaxEdTye7ErH9Y2YaYSlBXChizXqLTQff5j1GO051F2+Q4fgqfoHzCJPPZ
nfoCMKBRhu4bAKO/jRP1b8snjHniZx8DT+FKfw4dKEJ2CPPYhVPMTJFVLxcnhFgisT8zb7LxYM5N
TVTOaLOjOPU+csbGTpeLc8r0X9bfY9zR09OOd74l6aXIaOxbAu6mcIUov4N2plH4NvRstv9podx2
IcguDTjkZ3WchMjhGS1Kfj6FYbU+lhrm+ZiV3ET0zkZ/MNc9gW1TzuWTDMBrc/F1yDgQGCSMKQ6Y
tuPH2rDDLT9z/qnpxg9FVw9AreES0houxZohUEFjnN8d9kH212EUmaxzt9Jw/0aJaFkU7uen4Owi
t8aPgDKa3Fl4G2FCbsufeUgujaJRbSuD8N3gDqNofO7AQ1GQtIrVIunm/0UWgZbtgNfeNQ6Eqhm+
DbdYpzBiAMI+LgrLzdlcd7Cesqlv/mcA4Y6N1yVZOdsLnF1yx4o4/dUOxjvF/9m3kN0JeGaMvMp9
fqSsvf+uhUCuVzefO1WObONlMvxSCShxBe6G69JpY1b4moVC/S/D49siUkCdqRniiWbpPgRPgW15
IT46oSQoV/W05l0zoYQaPzg8FBYMfvAWANV9N96kaVVyg/KQxjh40CtEx33rRPg9KUfN7YKz4PAI
hZoHqYRo5KOjuEPrrb/aQC2I9kcInun0lU+gIFvn98K5Tp2bnjooOYia488jKqIC2k/tFsQ7Q9av
Um6mDqUo2qyMyw9pkPx815Wvv7UCopl0ve+zQM5B+s8jIIFIP5CvyoiG6PpXyUUo3zQpDA/wpLRu
4ErBkmrGIMqUyUvosHzF5L9wNrb2Co0iBuGPJK587Lfp05qxHOfLPGqoGZgTD/xMQjzJgUQHBPVt
P2PQ7sStYaPH4fnFFh91L3Gam3umRkErZFkFcVWiCllq9v2ADSHiYisZ3ZiSDa1QJZkiIjXq1ZSd
9LqvtL8jU8jTmfV6J/kho36OLxAlWTQze4TdQqkH4T8CC3jryDRklmKuY75NwuaZpOVgbZ6kGQLf
h9MpQKjpAWplTOmBfTsqgVEmV+acYRJ9FsnnJ2Z0g7Nf9+wAwJlHmXe9/a1XvlNojxjVpL8aXbHx
14/Pi0CtRgnf24JRj1TmJ04OekgyjO1fepWGv/DIy1KgYjzpojoIIWt+1CKlDB/d5uJpxbkrk0hx
B3ZX84p828Tl+rK5tZOcZ3XJLr0ZTPvMmxL47dBYdUNh0ZUrfZHtkdBtnetIMkRVcebLVFDg+K7Y
UeQpcH8RqRHNNrdFGB+vkuqQzjtuiUN2vQUUBcAnxgrq/O+f0l4zKok2cpvuYQgOeps0EVR24xCz
8YCUv6DTXPwGpcZDYfzIBS5KEJQIose/eayEPrV2G45cegAGirns1KPlwo8a9RDyUb5kc4xqIl20
p3nNH69u3AVhLmtAEnnVxJ0I32XJJEi+Rl9xf1EvCPx62jtzGAhU6Dx58p7GJsXV1PFNZXRGOtd/
QhZrbpnNTZKILeiqzsjsoN0ryiff6lJXqr/lk7rsknZUaEaMnRi4QcSLjfz7jF2VsjDKVZW5DCK3
LhmLnHWC+3DiErPUeMPg2XMPf0u2xJAhQGCyisfA4OT42qksOKVTuBOe8g2LGUaZbzsCWan9pMDU
blojW13S6ncgw0Pwekuj06u4DKsj+i+U1bix6uXN6Webn1zR3jstoI19EzLwVACGhufnzy6hJuyM
GZQmj1mskXNVo/2GgATxf5c+9+doQrTJsuuZT5sThIB+tqzi7gGnmVPtxo5rL+08ykUPZPAN9rD7
AYLXBNRMbY8Rf1+KTe/9tcUvF9wUzW0cUdy1LVRebKg26E+N2d12YeiKTRk28cgYPYDIAAK18J6x
5zg1K8mvcEddR7FA405OQGnmUhYE7qb4+3RNBR0HgOYXxEbomU8AS1vrLpJdRN8Dui8jSBKmREjj
3v+Zhz1k6yFWpYpAbb3gr82PeioDUfeqHw/19pgYaFHk2qhg5PIvuxxqTk2ws2caVXDTYg+Dpx42
IhKlIqCuMeVx52HRj6ARwWxZKYnGuIZSPYR4tWjV1Qesd9rItqFg3jo9F4rte1l8LBMt5jzMzjg5
eZoLnyTU7XKtC41fbUDOS0iSVAi0gJQcK9Z9T0pJbRgZlxlFi1RELckMwANL2KRYRcbqe4CaGN17
0CMm0GwrLN6u79fkx9IqUmPW/HT5g2Uu7I7/QrhT7tQcYp3UQSz+X5BUNfM6o7yvqBYmPt53Mjbm
fHw+jmffN7WOOftFOPyn3EOR2yRDE9Jh71N6iRWY5z6munkWbw4I2am1ujXqDyrphGTIrHuncN/t
gBjfxYrBRZT/fczSuXSorYf8FdMCT9QtyEhZLBc468DCS55/xpcG4KIPC3J+aqJEP9FrNEOtgShA
RuKCMrN7q45q9TGnfqVpZIbsRq9TLROmqa9c717XjS6CgLJPVa42vQfpToeo4l8GTfRh4jBbJpvK
UrIZLqjoan/9bC4RZkA84DgFeZ4CJhVX0kGJjit9Y4S7/dAkTLHaBbd0G0uDghukIKDyjvR6g5cn
ODOoi+AtHRy9JK69D2Qg2By8kqsb6gcQDOeLT9iaRRawnhD58WSPXiKFY1SOXzlv5i3hRQMCIZel
hJhwezcOvZVHr3s6JIYyUzIR7CnqJ8CUzcTcydr9b8tvH6jL/4Kp5qZBt9GHLOfEVqrounsLymxp
DDokHp1h/IS6nPkcE8rxyi6WYRthFCi3wmJJU0NRvdNpoUzhXFQ07xuQBnMD3c9xvzbgD4Skwli8
KrHNAWd5IUkPIqO3Sp4//WD0GJk7ZZd8LK6IXYc1LHHjCOjD+ycK7vxZmfQatEtifCOzWMJFL29v
vQx7JkrgBse8tL53RlgkTWtJoyjXvt2/C2sIn+/GflfCJyK5erW+aXHDnapbxA3+Y84sKCKjdyJI
dvePBePGu1HuDVrV0yYJjHFrBGyn5tIJuaoe6YtWQuQ/zbm7hXAVnSC3suI7RoGSASdeedwtbDbI
43NgQtCb58Y4TOmtUlZU0QVw0m/5k2biI3DnSHVyp2Y55kVlxH07sqKARlfHZc/f+W9+ClHhW0s/
SXA8wVuJhXkgX2TqluTQ0ywOt6sGTNBf9DHQ0pLyM3EoTxc6Ql4xsBH30V77ezOeAQ5OH+iDHKOm
d9Jplj3ewilFuoX2JyTY4MWGcdyU0QWU9CJGxxm/6w1OEzN841PVSS2TaFUDg4luzCDIGi7bhbVe
h7FHQY9FSYS4GNVVclEpwKz0p/HVv8ACIKmLUU7d/bVa42e1V6aeKiHdON8E0ZnQn49DVgqrTAX6
0hVytLolMfk21ApejFUaCTs/AsSx1/apJWTwCA3BjoZccYC1tejaHFt8XsBqlymDUFJRJ08CEpRR
Hj3um72wwkNsS02HkSM9nWDLUGklmuu9lE4kem//K+BLbxWvoSACI2OjCMgcCY/yhA2n8R20ZwcF
WISHn7SYxREqmzCfuF+cyqkCmlRjNjlyewTrXE0y3IUEgB07EVE8AMC3H/8mrY4P1KcE5ba98/RS
1P/jneZkDMXA9mtqgb06c3pIuZlAhIn70bglH3Gf/GiG14qjxbnIpwkIo9DKXiUY+FzkoNNCDcKr
ynxNiHOPDM0xERLlm0YlvZIcXBtPXVbhW17O96iLiK9g8pxXcFum9M1Y1hhiFjBUukA4W5nyqqgB
O8DhG5HX6sfhOs/AuHATucPDiAqrA5HMKy8N/PKPkrQ737Hu0QDLwyMvZUPdbmt7dDr3uer7d+Wh
6wg+ASfvRQB6Z0VfCDyU2vgguugtKTLW/4FfLxm7+VKjeKI47WkuGP/JcwFCOHfjSdoClo2mNJOy
vznJcczzEeN/En9uac7X1jdyScJBKEHpcqy7FubwTliUmvhJv9VbA+GCpi274HQTOBOzs4UWH+jv
GEvimghQJX0wTe17LOn1rtoeOmAni8Bdft1DM1bqV8nF0Auu7YLldG/XgbqgwR6HDEssSIU9ceU/
CPBQM7t/XsYRF2+h8+KGTB/RIhHktr8pBW1VatsrXFTjlR0/8jC42tzV6HnyLqHcpPjH3MS1lRvW
ODoy9SGV5OnmZL8sYafxHaTI935e07g0EFaX2ldF7dfyqtxEKUQffJKK1JPzM4ETMX3Jba23241O
m9X92iirZGt95MrQRpsm9yQA0E6m3P0rMfatos5llkYb/HPS4mRK4HLVlx5ehF/xjfWYq97Iwcpf
krjL8NszuOmW6YQmNE9w9pAn08QfOiaA1/mcfaqoItqpFr5psUFCT/zlbuHLLn9SVsigGD+PAMaC
qm7IlImfpUnc7yEAly3uZe30oNLTAkh7kGmrfZvDd1/TBZ5f+Xl8cS3gy/nqjM7NQ4SQUjSXqbJT
PogQJO6P5GT/0lqiSomf5uWHulnV/cZhwPXWWeVZ3heFKfw4Evzh1ch3oTttxD2ptan6cZbImlTQ
VA91qDMsZy88IkccMCgM4Q3g1T1YBT0AM7GAaVpOwPSdMjSX8XpxScQsRgVVIeRvnzTBCRR6Fi1t
lUDaIxPcn9SjT5RItM6UMfVO1bFVCjpVWR/I86j7YzcmY+tbG4qIgsX05XoHFVZt+6aBoWG0zLAu
B+Hbr8ghyo4rM8Xf/5wvtKls0CCuEJGpaRCSsW31HWgVBGgV2BhIiuXGi/kxeSWpGUoyMF7dLp+E
XfCesqXW3DGLNLhRMMAJNfzSWkWOcBnyoOMCYfGfGwps2uoRVfmMSlIVhExDnZ/qsTPRM6Lfhpl3
CGEm3zpMD9g5RXBHDKRxFevDbXkfLkKdZMfiylIVdDh1jl84Nw7vdO1H95o3khW12WCLG41Mb5ga
c1WB+o1pzq/I7sgm1DE6SkaGFh25CxJtCgECjRFWetoTLIpWosEhq9nuWtXZVBXrDBUuBLk7gb1P
BNJy8PiNKt3Jd1neohDr0k+y115fGnUTkK+eB4hYJHBT61Jz48o2ARU/nlUbuh7Ld1pCppsnQoCI
BjHOC+LB5rcGCer/o8glANULb6Zbbx8yyEsUXOvbbSy+pv7ePqMhN6hVE1ScrwfeYuexEIdf6Evh
Rihn3+TO11DT0Z2sPMP7cftelHq7vJv0vvU97Wk5plDKrhvXfUnanUY0n1/m1aMXir2hkDIDRBoP
DasQmc6DFtQy1bGnFDmYuoboFFrNjViqR2IfxTAq7KIjSx3NaDd0jIvaL20S2dg+4jlD2o3Y1PYD
iJAUwJ1YddtcFz8mXjVKDG3TzkKiYPfxtid/CZ934OE46kryZVLbiHbUiu3fmOmsz3GQABq47gYH
7vywwWDrFXGk4QyNt/0Jofw6sgFBhbPbc1LmLeHz3TCZj8CBr9p4l3iyzA7F/scjTEOoDaAjtiII
3vwlps23JRA6rcHLikP1QY6KDlLIXTfFpGG0ZTCvBoiZ72Gg0L1MTzTVyGuoHe5jyPoeWq6UPau9
L5KOGAa/B5lVeSoT3+ZHbmzNqA20pQ5gid6drM2lzARRqI84A1lTnIbB0nss4KrB8vTISVSdtIvj
hrJTtsR81KnjDCVS7GXwCeRb3rXYenAW749gSTNBKHWghkkKH0Ffmqmp46StbxegTuF3wO3l1ZTt
OI91f5hp57QkRjFtWwXKdxDyrIo5HYiRzh/T6OaIuLxr33bt/DiRDZ0qdybExmKelrh4IMqOdoql
dkTW6eqPEbDSHILg8j2eBX2GsEOkh4DukNUO17XaYPjLX6p1R3X9uyrO9mk+PI9u/MP1kViHdtes
zLdVpMOVfQS0U/9Bz+ibBjCDR0KVuEsVKuWynTWHwTlCf8OyM5enE6UwqdrWkqET+IDdKwKzOX0R
PWFilFyKabc0ftjzjiMDFMhIaRrranrC5jOjnQ4j5niibwi9W5OZ5LAlf1JLE4d4JXiW//Jj//I9
WrwhKQAhCQ0XQ2COlEuJdIg83FBwpF5y7c28u0zbPjhu8a9M+5sSXoxgPwilHbZMMvd92qICnkGV
rrvQbL2PB0nPi122JOzwdC0UxrhxT1LbcrD54mrI9H4c1KrM4axWv2e7Aw3XaIDeT3ovWvSw/RTJ
AvsXxFT829SKKNfVUm3GcLd4KbDOzzI489aC5pawzTxBBLSxu30R4YO2BW0sU5ggHSJ34Y/Vf1ZS
+5XE+M+n0Hu2fOEMz5NsQV2piKOStifo7Rr+2BLkkntvg0xz1fwghPLaP+m/hOSasluM0IKk/F3V
1zIXRd/6t62YZ1s9dGXyQgGcUwCwzFgb4WlidX2gh4wal0fAq8tl8LaACmL655DYsZGKAcXd03wH
KXwXA7arI0sInNKKh1tbedNB8+67E860D4+BCOd2xIOBQe9kUAkdN+1LrQ9i0AHwwCjBTOAcoVpO
KvnBkE85WhL04lAsPF5uYjWcDddxYGnLpRCNoolxFiLdtWr4ShRYqjvITNrSS3DCsia4790cOhC4
9/tQ+OUO4xJcKw/deeZE4S/fn8DEpQUgwtEKoDCdQjVpP+eCy5nk2QwaJjFJHa+tyOcex0p8aj77
4LsXPomS+HSTC34QTeDW7o3YJn4SDDosv4vlRXOaeEItdfPrDxPV7Du8XVaa5wmnx9y22jShlU81
z5JoNUf0VlvILHn0x3fVvqgX4e2rmJjVp7SQ0mwTyvnPmpSvzzf6GZ/39DLivZeAqe6T3BFtuyVk
93k1fF4+bHQ0lZEgIItZckFLVQ/5BwyR+5D1hKZ1JIFhBPgyMaCa7PLzcIrPs8tdweXufJoB+G6o
nAvi/rYLJt+Q+Vw7jh6abd7UsdvDZCzfgaaZUkZrA+m0vibdgivIz1N8gqh4aMEpIVqZ5DzrFpRc
+3cx2YprP4eVKt87YT4sjjeiZn+NogDM0oVj2f22AJL3SQY0FdqLXYHX41W0yaUG0kccG+hih2GX
58FGD1eC8IESvcb3k2OX8QzSz1PJh9xNDrp7LqvmGQQUt6A8K9H7nVTIj9T/ongesEJFTjCdpjOw
u8uVuupx69e2gwrzNdj0D7XJbO/DRHNIlOxK6HJri40EGMlIxvdaWuGn8//1Cy+tWJxm9BkeFBE6
8K0biTUNXvsnW/Cr8zGEVEy9i/epysA5Zj/FJ60QIKfK9/RVmFgv1NRrQkokndeo+SG1CDfmx8va
K3oEjYReq/NK6L7cy2pyt1IFmGybQk4pOsfcfdhqNGKA1OLqEDCcEP+hG/iOc3Osvqiki5SKYJhJ
dssFP6PX0Mg1jYlTeZ3tkWI3hawcUh2zbK8R4Gc7cx1O090w0zwoigDdTY85/36eO8p8wD2EQBan
jBmTpzlL12fSH+IHVsbD6i5izJGvIUG2HvCxMiiOu4wDItgMhVRY1DiY3ksAIWEkZHgUH7LwXJ6w
f7o+j9DTRGrOOwpFWPL0hEG274dnRQa3W2leuFFYopzJbC3y07Go7vq/muqy8DFkbI5H20IA1YAm
uswM3GMzKn6LMPPFA9CigU5PM9x6XW4Qw1cy53lpo/VG4MDm7dPX+XFnL01+SHBi7QGz51depC7A
aqSmbvOYMV4mvINFNiJJJwfb4XuF/e/gGZ0TxSdGkFIHF/G86EeUoM38VyPoKx/Gjmw7r4VKVQw+
v+cB7YdHWEe1O7jymDcGVebUSmMhV3eH2+qjkXmVwOQps8sUqFFS1rgvkBThcRfnVhPNyh/f9owN
XqrPWUeNsfmpghIVKJX7wKWkZUiTzQ6m9xaSpErgL27rE3QUgqgykYB3Y1KjyHvmxoAGC6dHGy9u
N4M3qd5RmJErtq80c3P42z9Y+IClRUCv8DJoBafgJYNE+L+0lNJkudQqkkb9Sd3Q3y90Xp0qa7J/
xMvdspRBE7/VBbB5JmR+baJrvu32BiO3VeUhvXNbh1AqAOZ99TdiQSpVKiPzFxgT7UIlQsiBN2s8
d1QfzbwrzQTdxEmnEeAj1PYYkxnSAQEFiKvNLOMnOkdWVpPBIRZyJ38Cn+m5y979Duy2kQKjccZc
ipMDGXiLZXsjqiNI0V5FcuJPVHEbKQA0fuLtxgbtLQM8G7IXuxGcf6zYs0ExMyal5x2FWtqGIj/z
zyx4tnf6zgI5zwbz0o14T+VvYJQAjOxA7Md+pJIjaXOMtgbx1FPAIMQiESKkJN4zfEEX73RNIdk2
Jd1VzA4Wz6hljiCEoKm793YYprPq76vYeN/quehzpbE2qymjZ15C2GrmexkHj0BPGIXPSx2mYH5M
A+EKtBqVKXqiJsUu18WjzAmbzM7dfpRW5Ym7BdTqqRQjM5EZ9B0YklVkogTSxK63DqgvDa0jS/Qm
QaPeCg+Q8HbDItbpj5lInJaghjpPJez7patEOEWS2HxLePQSLX5Fb55kJYud06Fm9wTDDbnccb5u
cEEBccCH6/DO3vIWhBOaksFEpbuE9AMSPYkkweJfsSoweQsSv0u4ENQDdz4eEtNKfdomdGaxzsFX
E1+zTanBkmOR+95UR0+pPNGQoBe/8NNBp8hkYlxnvMDaeHvfKJbk3Y+FW2FRC3F0pCmymyUn8qpa
6hN3gFK7YnrjpJ7gAEoeYXqnJ4vfPlWgl9HwlMrJgPWJWokRoKVTAWiMFp8lSoTAxd5hcKRTWw7F
vWhdsaxR3N9Ga+0ejG+J5V1ZAi6IR/DI8jqac2dciZ3VEguVyMIsq5AahbfJOkRGrRvVPXgpnXLA
4OipPW3WC2rmR0ltiNEZqQfTJNNXsxXBaXHXwAp/Xuq2FGWo0zWfD3AZokb59Jln6Sr2fvQkfrxy
YL2KzSBOQxGDgLgR63h6wNTiinXuPw3kJhTFv10L0CBCbnKokuS+PAvLwO66DeDZHPhX/UMXwp1R
VT+Xvh/R2sFu0ZAfKfgU8usWkrnGg8zNTYJrPZA8Sa/A4WxEwPMPme1zjAzATT6Cgpm9elukn+0j
eVcun2shriGgw2xt9gWL7+NK/1atGRXElTH5gdmXoa+50axc9sxDkXZ4TojmZ5WFUzV5/SgBXOIK
kCkyEIaShomL/ibriIslF17CU3S5hrhIl7TsA/uBt1G3Y7jFaytd17534YZnuNSpNVSeC/TdfrEJ
R7aAO/ZFdN2+T3sWBDNktexrEAs+2ANKa2VbgK8lh5fWbAhKQ++SJAVDoNloRKcH3z+znU2vw1Zp
/wkQowWXwfmijkHhYgGLvHhhluf7SyLHrTjnzGPX74ErZu6xbZM+YoKQ1fyLzi1TJHq4ICWJHiXd
/5hFWfnljcfDB7Z6Uu3Q3M6KJNVKpcv4xjdwtFw+IVhVnAfB/xIjaa+EWY2Z/kg7PlozpW7zPVtR
g6ypElOQKw5Lbw1tLwLvogMNQf0sH8rJAal5zkHATyQ6EeFLb6xA9/rYSDZpvUZhoKK5F46NaSyo
8or1ocAE/xeP0y997/vxzt8gbzusSbt/WLZWdXc8tP2q+pOyUj24UGA5O7vb44HJvjYP671hwiTD
DDR9IUKjJL2f3JKNkebl/VvhFEAx7cmqGqgXEggq5ZE6yWAErOWMbiZnuuJofikHaIar6Ow0rdaa
+wW6KH0SJTxYgwYYqcI/SWkAv0zDGG5/kjvX00SpkpAA+fZrjmeoqSelYvmT0TtVY8Fg+Rs47IaD
NZSSqLXXmgWx44QMeBhISbqMog/DIQ3+MdzJyUCQyd4Kra9sitAv5CnBktUEmXn8okb9uWkJrQz/
zlWf6EzoEiuAP9OPTNjf2Ajdx5J/IZwFCpMsB85CjBA6k/ia31Br7SgdVJ7LbHlVcLQTWH/1zpSA
2goUJO6Gr1eqfkovxThQc4ybO6dHlEC1YD08uGGwwUjHlk3+JtOlybJiLxwRaE0viD9WyTiuusH3
kefBmaHr8szDgE9liYDqcKNb5yU/3ZH1mpZ5KSGsxuj5SUoGpQZpq6yOAGxFclggw3f5QRQYOgCk
Xm5dhcgM5qxCFgPckkEjMmoRZq7fuPuqttg5PLgdI5zGv2cEK5a9dgWlEah4Q8KhjxMKKWQH5ebi
MZCT8LjSShJ0incsFiCqettxoXGXWH5w0E0JaQka37TwMxpO18u2pER5H73cPWMOXycCIUwKE4BT
+ZqHDJrlf44oaoNOuYH5++hZtgIW8+tPK9bCWc4PlWp+OHIWiB3F9S/cHO1/Bqw9c2L3B2HPQ0wg
AuyhBfIjgT15LxJgijidwIJrT2502vMjxMkUXhayxAj+vWZiLkrRxvUiLloFbG8QMTDCvidGcxvz
zFdHeCYmwrsnrYlIJK61ZG//t8ZHiao6/OtBrDrXsmrrx2rBF6OxKUoqZWetOWax4aD9xXApBVcP
AhYhaJbrRdT/8VO08psrMAYM1wsWsYzUQMLu9jhf36X0KgGzIEeUY++703Zh48aA9sgykb3hS4bG
0sHJSsyJsovkQCKAyCq41rC5oPb5ffHt6pET/dax7CHwDBSSXjzpxD81c38ehV4CFJ9Si3LL5e7a
C/kOEXvOW1/l0AMppCRJzmM2ZMYsBPUG2XDSLmz+BhK1oBmOEgOEepMyeE9mfWaywlgMb7WBed90
n20G8b5wC+4K2oZMTyqVu8u8hPOv40PPJHi5tREm4tHZdxpxE68ehngTkVEQRICzmqznFcCLHomW
vIb+ciqLjOpFB+V3JlX8jsvVI7PfadNIeDoEwzP3C7ToVNmstBaFclc0NdwdSlkxhlT/8H92pKo3
gylm9t7Fcog2Z9HuxeF5fem4a0Txlri6kScu72khINiEVKIcNrXg0tlL1dtUB48NsK9TBzzIX4eV
GPJwHJdxXirbzQ83a74LyIznYPhmiy4p77FbhCVDt/nUwh+jDvPPHxzwz3Eds0p0U4w/h9N/ekba
CKSqvx21h8l1AZ2UtOM5Cd7SFFZkFQwRjLukN74iSTRjAC6mHe16ocYU77J+Y0ZuFFU+r4OgkW9/
axn+Rs0notkrT0psWBvpKUeCmY4BWsZgte1p/A4D9emnTMDGOpnwHf3msFjVlxhH76aHpbzqqtae
tgx0vgfK/HWl28C0ATD3ZqTmUUugiV7eibND4O2L20oNcmJ9/asi/5E1IPB7Vb7NVzcAmS37ydLY
RTwukN9tDxuwulpETVZPjcGCYxf41eP5RqR6a45D2i/xs4o/LYkHbTLTpU8rxcIUv9iZ76eOYBTY
YtOEfUGmONJcwmXa79W28qCpsaWSahms9WXi7UMxgIE63TSBGTmaahpX7VJ3F5aochLsDgoowaM5
//rQJ/fWLsqmXjfHqW9IhmY05hcqNwtulQP3vjdnUblYrka3jHNaH5Q+1QecqyJpv3apLgB5UGtE
M2aVJ5IPBiP4kHlKymF2I2aj1Arpa5JWLpgTfUWucUBLVFwlRBIkqWdQvEI8Iks6e3N+QyuUlqmS
w8VoLliy0/6pwQ9NWy3Ba765VEs6TnB3dTA/+4Dkb2rEaukIi25h1ef9rSmV2lAYII1KD474StCq
5nFALzddmGMKfp2ZcpT4Qu6lg1D4dv+NM48ta1zVr4cU9Hbn0uR8JYbOh0uN6wGHiM5gHeK6HpZz
71DXj9lyAFcxvFz2Ltj9NVLCk39nJPklZYlJnyBlAq+sDqr/MY3ziYfruA5QCsozF8OLqRBuYxx4
eDmc8U2a24wvrnHKimcuRnZwe2gigoGK4BqceuQ2fwteZuLZLWyJTcXFW7i2DJM0Y65+03YCL3Cn
cGpXdO1bu36Nbxx/1gTHhRdoqowNK3HAERyYUQ0uougisB7zn0fAjZhn85zI9tZZ01F+nuC9dFLm
OgLmyUlkogQR1PPsx6gRz3HVrSmbkChvGzB6/G5nfiqMcud8RQxZOkB/Ml5+svpswS9JePH5FWOL
Cg1B9gqcKutzy/oh/Ll5jzgEoFWJ0WfA6Hz9n4vqQIHRZ2swvqgc7JwfZF/FnozT4mpLOvFr/4AF
us0L1EEH+lnz0fZafdjJJjmh9QDkXdfqobp+l1FwiwSfZT4Ki7vYWdR2Qkv07Z1Evr6nTzSrmQtR
Xo5GrINfA7mwsQlCjAqMfFgUJWuDjcC+JRFx7qwrUepnHy26chAmaL7XRF1YOCSqQmYZl3gI4oES
1WSvigb5SrdeJyldOV8MF8Wklie+hhhdc2Ahv8czQerKMZWrps3etYeieRetvb4oeD3xconCns3s
YxVgGHoc6peBopDKOOXHYi8WI/oYXjl9bshem1A6YjxPt/F4yHQSmwuoGpHpiI6MRO1SYXd6bibE
7Vk1NKWpK7RLuL6s0gRreHtIZhtAsvAavRr0QKaqAsauqSjEEfSXPxAme/3pLc39WyJedRxnWXtG
EJGGqUT45IHPwVQ515S9Vr8NcuuxYFoGjcYkL6/06/AXbFAk7FCF1CFzJ6p3OmSim4/pxozS+3B3
cKKMF6/8XuRhnSXq7GtTv6RgnmhqcRCvwYOMnyTmYIBapqqGkKjrLpGcfOqJjG8C/CFarZ8plreH
dxwTwQCJOORT9nDCxryUSgUw2OV8wKOe7ai9UzbRXi6AuDQY/wOD2v1s+6JD7Nkg7Pys3xQ9pqHp
XuC1Lg1KmhS+fQc4PmULnTl+S9Vhw3kXw/g8GLbCmLYPORGXRpZwVzIqgPuXOzli2XbwtqMf+nm0
XnTfyeXWEvMH/xUDqmuMvsL5RnDgql19M9c2dmrDRb7EN6TGWqMnyfzap9jXZu5Ww1mrFLZ/SXYO
WeqShocgm/hnjBKEnsURFwJOprFgn73RlUVu9erA0PZf8BuENcLHs6gmYwTHr9HgD/wqzOksrAry
Il+NCwIDjnSMLJ5TOlW5mJmMvjh27dXO8acP2sR3y6SecdZDaMJS2JzJ2eJHfmmyMvz7JBgNDg1l
rsCthlMx0gRmpYnfVbCrkFn4JnJYDefOyfvV+yPHhc4R2OInGkDcfF6ffQZjISeVJP1xEeUy9TsL
z6QAM9+iEjDnau8/P1rjyKxqaOb452v6Gv/YSsSJADYUyx5DPA/H7XWZWCljY9zaTmT+RoYwfFlq
UAi0I5ADKb8KWEGuH9Hp/XoGDN+5WL/LHiPth0JEvs/ybANltvFALtqVmoy1g0EP5/82AIMqLxLi
ioQnIVkpjDJw5/U0oA4BUDNsVtZDUudvFCy5OtJeL/+zMdYsJoZyOJyeVJGlQ/sKGSr0fbc60rVG
LTD56/gGzJO6UUxoiVmtkroBWdWsC7mkuYxaL8EgSMo4wBmcI8YdW5CyXFab0xkBIp9MpSqPrBMQ
ibPjaiI1HSyz+eb+SCK9iWB6vGHSGxMWy4D3JFYs3UqR8IU6kLL/9ERsPXPWc29lcFVrZUMChCOq
9DZOJM2FtlEfp7nIyxqjAbzaOPN2pT598Qd004L83ImbGQHcpGpnDvOn6Byv6VmgRt/i5djfZY7P
APzCmBieLBkSYVSYXsfp1BQu8xiqzzRav7oeVDBnk5NM0SJyhPZbgDUpU3VcHBYb7gPV1Oot2MSG
zYMSbWei5kjouAYf8BvvdAp7TGxkmp9NWJMmNeap6Xz8cd4riPSKW/tZX58C9nH8UkeDocNa8dhv
2osb76QzXnbryAo7HspYtD67pVh2E01OyvJ6gjvcvs2VZO2NeBk6ez+0iOfoWUKTEykjGBGZWeS8
tADM+CfHDRXYGHo6X/JZdjJ+/Ycy6CmZ7QXb3W0LBftCy9YJRdbuw0dyHdCvPQbXqaM79gi0xSer
miTmTUM6+4E16emSANCXA+PDxNnPYje5QCi4m8SbZ1KHnyRud3dSOhq220I7Ng0RARrIEQJfPhpV
9nuI9+wL+iMsd3lHoGi87nWH+yHjqMpREvc/9nrum64vMFAuMUE4ERTssSIXJZvWzuPZKP7rV5mk
MX6wmUb/C9kgpa2jlG9r6ZtY/EOnT72g4upy0iGd3GCNMBR4KiianU+p3+ZvRM+z3Yuw/vn0L2KH
hIC1Rp9+kMEUGEEeIE6ngcl0hgCRLq98dvqjid9zEuMlVEJBnQ/r0Qalb6lhU5qmpgVQ3zTyIzvy
TqAQis+ioR7jm0g9ScjNah7eSH5LNmDmAB7QlEGp1yqtha99QULo696VX9MbV/iq9Jol5TQn+rQj
tKOMZ9iqpi/nj+jVbfXMJTrW99Zc6EW5SD+EouzvYKeiB29biWdyTBswyvSGWhaAXPzOvBUtP1RX
jIMsq19g+mXy78xNN+sWepNXM+18YoevVqK2WOOtO2Q3FZLCSqX/HfGwwvgsOhwVxQIJcVnkIatH
hGx+PRs4q/Lg5+PJmMZFyBPk1DQuonRrkptOQjgiqr9j//G+3KYL2JN4NquGv+EhuaXJYDZC+dWV
7d5u7GrPjpaxlFxM9P8iwVVUGzLLMiK6HPIUBb5S5X5JTosWspyx7MZpZXt0DX4BqkPBOoN2KSwD
p41ZW7uT2sR/canz4S4bu+JheQpa+dx+JhlKxBqcFOP4sZzmktm8yA/W/e0LLUxZX4z6pINZfi7H
XNO9Y97AC6erW2MH9rKaIgxG60KR6EUOwaRmF2zfUb1hYhPSG8/zccoE2SoE0zwvMXm4Dd8QDslG
3sVZ/gNCy+27kK/Yx9RYw9hsbH9AmvJrLinYaeyPukpNdDkccr+hn8cUfa5RTT778tzJVUD00yqs
LzZd6u87sufSh/i0mEka29/QNPj9dhu6LUgTKc2y1DY0Peof2/VfO63yHhYxey4Rs3EnKvPLHzPB
iNBY89gMx2T8iTvAgj6OmK3MZQaRjl31zWsF3w+S7/5Uv6lzF4pfvC6VqKVstYw1GgEFej0K3uqA
klI1YSXdiCeassRoWXHChCP4j2NgeM6zRIWJcW88kXZGbwo1UHEKmjzWU23ArjuUtFPNvugqlcE3
bCr8uAuzI8gYMacL0P/lYbgNuu7hrgTRnupQSLh38XCpMm1YI4EDHQR2VYiOrkdlxlGu6DyQPKN0
4ny3Mh3fuYZBJXfgQXAs0ts4kutw2pbwjW89nN3hbB5eOQSV3xM31/ktMJtIIFiBjG/O73a1DzRz
/0hjmAlHMt4M+cZkn10u8EXkEwOnCYh0Ax1RUSdn+U+2813KtM2Dihh/Xu7y1Y8Gd5dkM/EPVlMz
JtL8sCKONBRylOBtvA8MxK73huYrxaZqZ4BkxxrEHP+qRku8IvyI8gT/b7cL4d3/Ov58mql1qzB5
seK4kpYf7XiMuW5yBTlWPZkedTJWbNgwEnlCrh59d8KrAviouS+PwfMI5PqfKSSHe0i3ECyeWidX
OfYpvFPuU+DuBFV0tTzqtlh9ywTETx2dcMnUp8Wi7EDg1013DJFDu2X4slC8JvxbzdvkTRYJHvDy
kzul9qwtJN+sSbX5LYxasYOK2LQxN+2fhg6q1gGw4ouYKpzPIl3pq9EOUb+ajb3mr3gJ3yvyHc8e
DKfDeyvkWYQOrDakHtcgLU8oT7A5ZkhwdvNthhx1T4GlyX73oRvshLKYvDyA+406blVnlE/h4P+C
k9RPgd/MOy3wMVt4e+1S/dYBgKOA8gqOXYaXU2Sl6HPmQLFvHLbEqlRSlzslr6v7rrjfVHlKsIxJ
G6fpP6kj94NND0Xf7Lm+Zaqsk+ScZ/jnanwJpuljqIm0bLQ9TpUl7JMyGCisY7FT74X4eL+HDUfd
BR0wNGFcHOhUfVwcljRUIZNp0/olIlPUgzPF2mefIBzjCsNyrLdvw18KH+hq+UxiZJ3SAXazINXF
Q/f2eWfwFP+rYu5Y39aCl84mvNzEii/df5VDYX+hNtM2bl6SaxftsClZKskqm3iakzGJMyMOyfB6
asjFA3a2GKET1ACCMnOu2h4pNmJTICXGtp89L6YZcM8egem9kTb4Xi2G/G2abSXcnL8TcPTW8gu2
oPVGk1r7PR+4GdD72hKpKCm07Yk2Ke8rfn9ZWrl37+PwFsPD1Mpx9+5PDqeNG1UMUMZnnHm0Mbz0
gkdUaXwUKwmaJyDtNOlgOh4znGKG8sKuXvUIkqaV8PQYFWpI5oPdpVv68fzSJkYkEgcdKpmUDlJT
NGsb3GkqiCIOIkyCpPJTFkpP+OTMjPbO77QIDFRUPN0lVCdnPhbI0jgaY32T7cAnVvtPKdg/51k+
EotMsQjspduAjgzC4RTtXUGkY5WoiJYeIj4fHkw1EjJgYZKOa4xV2v7D8WII9i6hR/fIG/57dzPZ
SYW+/ZpNW035yDYMA7sq/2qgkGY157tZSOLu7kid8UXCHHkvaoJDdWhl+KCZPhD2/kPHVaPMZxA2
g+y+/qCf3wgnucnYi8ESXFRcImHwxDySgSZn2zHmSwT3xGblPMLHTUmLIqAVqIqBK5dOKh9NbyG0
ce8o5E6A0PgOMXbTWAhkw/lTzltDkjQQsp7zciVxJr8LEy5+1+vftiFJJl0HfuqAq89tQDLS7nXU
JrETPb27OMAATficJQJdXUyNC0IpYg3HjEks4loYRpf6XiwOjAVDUb8aa/8uit5Vw/CHkF2+CJqq
sITEyECyEMAOZBEL65IIXZFcha7LQ1q8+1A45j5qfbcpi/PgDK5RmATpkYwCgpPOVNBGFz4V7KpF
7JaDfQs7/xnkNDb/+UKs32PB/ETHGVPcnxW6qx4gq2a2B83KFeLX9a+Yhgi62bd4w2xBOXhy4v9F
9oxbQSLbv5ETh0WZ61NqsSlLM+5T4eY+HeaGxAAx+d9PSA1EewS4bnE4hVHA9mT2KWPH6PsM28tJ
bIGks18xXWY6bX4QoMTJdWKzNNHWza7x0u6K3ectcswh4SDU+YJftCg+a5jbrmnY0tYIvfq8Lg/H
+0i+wRQMfJQNXOiVUQyNCs35nnVyMfUVyWqqVSgAETE5UtHDi7sa/s/vDunM1dlv1QkwjZjVznfI
ByGoKRHxFYYA+81muOkND8CCW1eEzXIRWoawE0NexvTKyROOyY4fNgrOvHiDEqkqXipocaB1nJJu
g0Qj41aNCC+nUXwO3Jzd1ENQlfGdETJq7QOKTz9NZ49ctzOsenyXqrvz6qCfHFBSiPqYanTBJc85
YcNTFVTikjGv9G19uw83jiJ3UmjuIzYH/0RaTu4nFjwFcPpFUBj08XDmoTNRWcbytxX5eh8ciwaq
t9qMRQ4ujxqbgwVOtmhgsSslVjIkZD4nGHfWQhhzK6uEVijm8HZbfckZN4iskkboV+LLDRJl/IM2
dTqaKmmKHNFAzI3GmCxafgurdp8K5NwQEx4FnU5rVlw/BlU7diFs5zAbIp+k6q9Wd5ZOkXOG/Vjy
8BGdo2tFApr3DiyaNyVX7mRq4QQct2aRFBR7rnZGUh9fJPgXAFJqnnfjqMKElvw+/H1epMumEFBN
kuRSXuXg7QXOqoPA2wU3llWHQXVCKFCxx2iEUcVkH/qWfEkx90f/60bq94AJX44eQcGhwzGBTh/u
bqLwUFPLUOdmwTd4vA/UXwIOESAHxd20qIcvJNFCG1YVxkjofhyYfgxqlxN6lj8NQ6+TR5OFd7Ce
/nMvRwDJs6YBj1lb+yOhvRxgxBkebqauz9exwQVo5xCL6QZRXDMZbeqjExnyIg48HWHY7+fBM/DQ
9ljFlBQxWmSjqG0A/LUdMX96zIBZWwzO2Myj9N7s38E8wYB/XINyU4xk9mTd9H4rcg31OCOxzLo1
KxY6EBpw8P4z2Npq1qoCswyPIOw/6FywsRq0/D2NeWAors+Y63Wdw+HNgDYWFizKekMwcPXT0EFb
IhlPIfz3i6YuN6q5fPfPsywMxUS5zzMM7+8rB+8R/5JXe+2RE7X2SkTUhl/ECJdIQ9BDpx+XA4OR
+BvYv+Gg1uVkk6cdGMzCPti88SpDRtaGWYnS9vBEf9goeINcsEPGz9avKlpHdA6FNUC5sbLFTMVk
5yCT3WFdaIdaCSf0Qdo3lwJc7DQGUfhFkKGkTglhFha9nwC7wEIjO2IlgV2og37Qrs74+Y7eRowh
LFXAPUPN1ov6e7+whCp0B/tswCoe0V5BZpvOWym2NEVa0ccAF0ZIcbPJA4UEVwpDcDmihhHV8ff6
SY2xAFE+s1wT7tzhOudic2k6dOB5MtObv+D4eQOkFE1yZu3rVANfKXSdWmAvGg8PJMYSGH08emMy
aMu0wvm3yIr84ZHsdsAQvCulVEF8ZgKhC8lvKASpv1KMtcor4dnsqptHtV4k+oUdYedcwIQ92Bj4
+Smkll/XQvNn3ATYwZR+sD7gvvXfSaed/YW2Era4cCJs7145ZYXRw3h2jpu5wJbaOsqx640xyWWC
c182mApNH4WCZXzLrojFhNCJU+M62e7aWhl/Sy0krTfg+EGwDVSoklyTVj7YAS0AQxiT0R+Rjn4h
KmqnoP9UkosK8qZaAMVGZfbN9oNxvQP8phIRrSwdSi86mSlYVM3kqkk5BdyzVPMculYTwtmpWbWz
RQgNRGSccvftQdOMjpAEwWhdUQprmQkHckyYGOTcpiE6YCi2LOjQQci3hRqntDJjjoT8CuBV6LW7
DUhkhjw+DqdOYo3dE50WEUNmJw/RonNwIuvLnX/S2mpJL06nv7b0TFVodrWw78DrJezLWclcV0wo
wWUtR+uqI5gRVG6CmVbn3HF3X09jVA7Kjyqj2/xMu3x3bWkKG3Fd7nDjmb/21JvgrUuEWGMlBn75
RWuJ6WaJFj2XtPHEeVw39OcRZSf6wV6O3FMGsZGro2d6+sotIlV0Fp4UBBBvgRhToM0/V4M47Gpg
8jWWYoM9gG79G7YkMKBP5zXLLCbpbspNDj6pVo9hDRAhGP/LNlj6p/HuuxW/BTvpOtSCSnI/ZJWi
nUaYDC3rNUDzZ3yVokJi/k0bcVsE6eNUnk7Fncpt3JZc3tN6Niy4NoDbl5hQWYJRWqY/iqUwK8GH
Yq40tcmAwKHEsWsueMVZBNVFlg2ReaX/oi3kOKwkBtRFJ8XUPntbP7O9ssfoSohTZPcZcbXs82dT
0qHl931qGNWyJczyq8YumTmVzMWS0mbKRoGGuFp8fzaIHA4rdJ6Y22HTPs/wmjXLh6zmQG1hFbMM
P7wA7NTCTwRKMN/XSo0eH2UGLz5k7bYtUXfBL+EvaV2+6WLfbRsPS3GKWfJtxo/bUu684qOsOEeu
E7U4NkeIA4/XgMDsxA9NevM4WDAcJHGtWpWZy1KGUKbUv4J19aqrE/kyatBwhcI/2IN1P3NCwJJb
0KEPToN3mRcg7VQy/Xjf2MXy4Nh5zxx6zp0tTEh4dOGAmh838n2oDF8sA05a/tq0whgP1cTfk94W
mdbhe1SCdm239WBO09wvsuQhmrW5133KPApwntqNNdffR4Nnwtwh2Bdj1rDcHkHTfqExWiZ/2CW9
bHc5Zl+uJgUKFiiBgsve+00pv3C7cqK1l6dMmLJGkIpAmIh7usOu6C0STuIZBN3TLrAdlmOv+/sj
pU6Ue6YkaXKmBxMtN2gDqy/ONcnM6OL/JI/KG55KOqxqxQxjrFMlNGdF63uxz07eNYzclKtlS1PR
cjlAMBa6sqA3M4CKctf6TS/Y8uvH/E4vTPQli6gyFYf3VKIVrATEHS3CyQeKxjTpIbj7v0YWIe3q
tcReLEyQv5jBoL4TTJkxQTZPmpnE8TGQzpJav2sK2aAh22ihq433Cf0+cTRdPBxvBJu6c8V/jDyy
TPkbpmJF/N/9X9IdRSjkyG8jw9ohqCwqBLwgdTwdWTUCHShFpBxr8MsfQ6LKa3swfVgWBEqxxf3u
S79rQHfQy8BzpjGuoiTYKtCY9XzOBzXHhdr/Y4OlmRohD+nhZvisTs5InX+ErKRf1BEuuM0A5Jqk
gX7gqQrSg456xV5MyKDQ9dYDQ595ZfnjbkIq0p0t9ON1H7xHZ9QTCAaDxa1iJEecpe+VjacY/vq/
P7WHQONQRcA6+gr44mXHSGmJBgzYOhss5n3i6nYB4IhIQYy8FmLsEez4jWQUqH30g7hVfyxVNGd+
uZ7TWjoXFb4x4uYEkn/FZhFl8TfPtGokshB3WAb9nY88bMf9tZ4EBbbIbsF6Jz3kN88N7q+Dd932
U2dywwQHJ+NinQGSp8XR3rpgN1llpp6D2zJgqZUONZNOcTyLDcm6ChZnrmA761UgoAI5RjHH6Fp0
P7gV9Z+FuEndxzQ5kLbTA2J8ft00KSFEbUlJxTt+REj3InvlF9S/sbifrfAzuTc473RThkzf4sjh
s6k+GPNukoOQlCOtJULtOgRtENGNgsZDLI+5MeA3TYT0dATThetYik6VfqyzdFiAqXwfeGf1PYn6
JrH841AVZb4ZXdRvfa+bQ3/z391UV1iWdQQfJcMjBRq0I8bIjgGr4XHO9CwL2ykxKsYD4YAmzx/m
4soeSmngVCKPC/nX3aSXXsauw6RiFq7bSTOYcUxlA9tSQQDUGBVEji8pw4QAsoD8atnRZDad5oyp
hula8sdJWSJK1vS77iLK9GemudyzvPBKpQeI9wyWVkNFuvGLYFODixj+TNVEurh/hfooxHKFOkYj
A4jylrmDC2FBRx2fCjZ6vrNGo5ll55iv27tJPcR5FXeymgW3ZGvAUN3f6EXDDug1H9zJBfqAnm06
Axp5GUtoqNtswk4LaTQ8YXFYeHiyVp4W4e5G3yvs4QNuJfM3rHVxM8Zle06Zd+6xRu7GoK/s5qUQ
rNfCEyiGjo8VoXd5bFFmDvoIq6uj1yxz4AeBr9o6XEy2c0PzIV+ow8f0fmLl/Y7bIpt6Qiv4pcOm
UwMiF1qpPem3Y6WUbeUZX4rzs6jr1cPa2EcjySb+DuQd+3KS6OJtpLaxaxxzHUo0edXh9dcM/GtO
S08TKj7Bow0DWmn5NMKJILq5S31os5vhCBkZACxTR+/l9Ny+4Y6CdvlOadx8NFfCrDU6E3C7U2Ci
NJFClw8QvJEUOGtFlzpgkv6QxI5gBKtdpBE48WKc7YVO/EBmMxG0FUbTBdpR88JNW6Nz8/IzwYNg
MefhbmZyOT6vt0K8ycTcQ08+zDx5xjWhkY9OvHnz3RZBCP5pwn7/ASs+bE7ZNCQdKE17LgOw7eBr
SWuwGt1HEDqWqpAQag0O1cPMhDuZN2jHH2+TQicXgc/jYnrPg13gu1W8F3cdaZTnzFuudut749vk
YQ1qA4/7zdd/gCHFX36po1L/iTChl3QbMmGpFSA7WffMB0iLJXnnu4X+vbz97GdMODO+n0RI0EBa
19mYhi8/1cITGZRG+oVHi0ZCzJKLt/MdE3iN55gypA1CNYi2bN5Bid86CAfIQawzr3pasHUSSUEF
IgerKfcySrr8BiCdrOCzWoYDfm4PEuSuZQzdE/Sxr+DWBCouSvD+AWeGQaP+xBefZE/OiHUKcHH2
4qzPDzuBHrnxLO4glXCyY6J55Wd+YW3ts4F2kX3KRyuue2dj0XNerdz1sYuqKUfjt+U0C+zjDWHM
Y8sdW6GYz5M5oqXnXvbnx2kiCa8fFYWmzx9wvJANJaDEj1iZGGZZr0YUdDl/Yu0YneaaDej/dM55
ejrcMB+1hksv/rVsDd/BSp3ULDnu8rTuqk4zSDf35n7sv2nNU9ScfWZ+aJ+ZLQnkRYs74VP9rfVC
rjPuLTcT8bAG+SspQ7C1edcfjW7sB9bRT5CTilWvdU6Rz2ByGzVnj93s6dR6obgmSiZajmZMoN+X
MiNATaZvxsLd+ZWUEQHOQxmqA8JizmB3nxJcuJuTm1vRpe/mwmDo08mahC1V6KQxOK5O6LVssjIC
QYiZSIWNs8EypSqDyZFVk3liaOj8Tu17ywa8T79ka44lLod12Bv2vR7VThFGwlOInIiMXTKX85qO
LKqh1ftKnsOu/kEQiRCpW03iBTOHeqQuELzmEhnKIpwB+ZOmEK0tGB21s7lZDJgAWUsSZ90Tvts9
X/hfmjp8CkYJwEazOcBQV8LpXMi50y9O0Qlrgj7D79jtxbQKgVHiCDM7Mx08OauAtDjdqTjqyQlc
uJDLIHCR9COe9Cimio/uzapliG1+qfyo1U16iN42zp1PL0538JdiyGm3rqi5YUgvPQ8mwQdF1sI5
CeDrxcELmZ8np33w7nziBqL27OdR2enDZV+fJEcTsLyFJ20Sxxpj26YwOElyF0SpralOJG5Sgy4N
TUs7hwB2SF8S4sazLzBm4yPIlG6UjR/K7XsUZKqqDUAXU4iXJATQh/DkbCI2FEgceFbe7Yqtgk4l
rC+Lq7TyOjBnIZ39g+EIxxpMXAF9iYyoSDnqh64/C05X5UxFzJLjiCnUwyH+zG2RgK/vgpaPVJfR
VCrAGuC5gw5VVrtoFGEnPZGE2uldB2C6ux9EsGM45xZRgvfjnHz9bAMtLBMnm0bEh0bYr/lhhCNu
3muEmI5cUm9IZJTS3YZxuQrBoZmM7XgJC58XvIQ9e/hse5BptjXHM9XlESnsOPkZXIGnXxl2RvLs
uquTdezBwoYPMW91BlIwmxHXSy247rxEWjSqZmbg2CHBXF6csHPNP3uZoMB6KuLmARdg7kat686a
gigcxtyB5knzU+0bkTz4qzN4dGuk95BLjbpVb3nwuuPJUYJacMs4xqkXARhtSR39weNBvHclUY8t
YfwuDVGUEeKWoyBBzT2ApLCkjZ/93vTdONn837RTpuk74CeaJK4X4lN0p9VSwNkbm/1BOkbBFpLI
2c0iveqiLTMcEYJbfElLkSBv/9sfiS30ejwQFx+CzjHktqiTv2FTxF4LN9CepKs6zA5HC/YHjhzH
XXf+krFLkyb1N87IJwoAr8XyM1jFulxFibF+tHax6ftrZnQmtvJhgSjW3XoVKMYo6eP5VVJbD1kI
q/BAKvluEy2EtWgM3+EicFhtH0jHlEYSqvdzqJUBIVRvEr/H7ix4M97UOw4CjX65ZUWGwITJDAqI
+Nr2tNAh6lyToLN8wP81jF/v7LQcRUJRwD2bVEGjEcLRTQS2tqKGH0aRCguiB8ZZqmsut6tP+dPc
A5+A2oYZcAtdd7Y5wUflI+qnkQbyQ3bC6SzwGqFUxkvE5CP0XWVvhmFH9EMbEzooylWZeFQh/plK
hL+8c/b4S0AERwahbR2l6Ouscd2LpUeMK0P/hkal06rZvhWTeLNqIArtPIculD0V3HH3cOklJUhW
0XLCXspO59G46grVCpPGFljtZcARBtmgoh03aXUzm7479qQsXsKdIn4d43ZXlVLWSKJ5PekJOFI5
gYFV/Z4LIH8Me4znqZwjttrDgxToPNPEHntIqWLPy+NbbRT5TKGUIAssvbMHTvxfOevBeOFqGNLP
48tg7wfPBppsW17rokvgsVyGTOoVh6bnnDkmXWgi+hCC7X7A0FGAA+BLOUjbLrs4ymMQ/RRkqgXU
mopmh39V5V7SF6iTCvKt0Es9Xoct9brlNXj8YlcodeNSRH9uUlt12k7o1Hg7Fp9qgmE3sOofL4j2
AmPAuPRkyV7atQJvQ1pYnWvGzOAfLAL0KUWWmpCFOahpBUlE88kvS8sJnYc97ixMAVS1puAvZXo1
IDTacUtBnQOxCOR9FOq6fEWqbbEXkveXiQYfs00uJPUV5Tzubdcou27YVVsKLwKFPpoaOuAMYZrU
wLmb78SPSKONCQOzbfymfXR68d+NaxQpdlMpHnfaJ8l7Hp4upYF4mieeDiyO4lf3BEnFWcrxYkn0
72vOyzwkVTRbJwLXIr7b9mk1y+dkEQEn11chwx6DRHtvk5qD7Tt53Upzkj06Mnn9eg6K1FBHCMTd
mFpsx82Zo7ZB0wrTBEmynjLOpfNRWMIydpDczE0wkddDNdQos8QQ50HMRZfPsdCNSXwHk6pZEifs
jJCqo+c/CqSkkkOUQVQ43YZ0uSGq83t8AV8DPSTprJ3cvWrGKG9aFrY7QmEkaVztRGhW5xPZsLPo
VlxSK4XbYhDHNq0nBRXs8p7HZSimv9dlBldLZlWpEorZOQQFXMTCmdsG5E+gl550HSIjM7hxdbUE
EDCIqSdHwUO50q8PjPhagwAyaiYSZC/UHU2bUd67FoPHuzjxrxiGDXVcvL0uYiBBFrzJt/qFpEIN
AW9XNTx6DhC8cxEM9o60R6rkHU8n7sohs2KLx0dZCTGwV4mXZpiJfJGvatGhpBjJcDzxZjnE0fgO
ZY5u14HEYCBWeCQeiCLKY19H5GRNwRh6QNRP7lSZfU+oF4WJo7ZsCIcRd+h65pEE649lEAUbNQtO
IZFRER6SND9E3weawk8J6c5AvwdcqTL/wczC52KF0iXUyqWA9zJdvCXsesrAkjVRCmgN5Gv/maq+
Fhn6pTnOeCVkucOxOX/BAXwDYMjK/zyFHfEqPbrK4/FxMQ9LwDseSeDLTEA4V7GMM2txWvmdFJcJ
cPwZO5F/MwDmzLSuIM3p/z0vReWdo+1sqASGAbdp24LC+fEf+lcX+W7bDDU2i7H/hypfUB5F7Qmb
0CdEF73+ZdagDcUYRlbbv15xtJOU1QPQvh1SXQ0QnAyNJ33Io2Rn0Xkb2d+rkk/10aehS3W0PD0I
jRFb8DJrONp1lcPCFkoW6Dj+X2fHhtDITMdKmkltawoqorQfSuogUyCcr37WGmeo0kNGGBhHaCUq
QJUZpqKEcXBpDmHdMubfJXL07SsMeTvkNkVHvt4NQjpJZTb8x4txQ/nQLwb7p9uFvHqsqUZ67pwj
xG9jghOO1VJOutAK8FAqWUGeo3TdpfpRZufPiUIYNySwLF5BHOyQGySvKqwEW9aPjO5Od6e5S4Yr
Tshd/utvVV0gJsQdq8PfziPXopOZAU3yAewHc+1SQobFXibq/ZYcFDS0WAHAoyEHujZn1AefxrXh
N6kxSQMiOENvLy19lZ1WS1f4mToI07Ge3i3XI8YfoglMY1+RQzCn1yr6NjS0TdV1D/F+Tx6hKs/F
8RpyzMXUYBtda9nH7Mq7PVUakMm5wcJlGgi27aU2U0yxbkL7fnr0J6ZTPR7Gz2mCDQKuIkKJdmI1
BYK/1K8HhlUBvXbJsaVEnic9cBbtPOF3ngphr/gJKm1EpxQ0lx1dU4m4lJpJCYn+mpKvLOgU1sMx
iqjm0+wyEwR0HEGY7k7+FyLJDMkujCfUad+QobNS+5cft0HL287loPSkvLgcZCPWDzhx0/yKHZdl
WdSfnd2mzMnUnOorVet47UQr1cDhhCdgcRRgh06uowTY3wwb8lgyBPBwy64oxh8XmUbTW+UJ3iic
q17/And0a5HTcM10NQNuhTqjnTm63wJSttMuJnZ0SuM8ChM7imGbz8uPdRoSlr/nW0Wp9a3/8TW6
gQqcemZqtCh+wrE8u33olgDq5tALfpOW4XpHwNPvo22dld/7WS2nrEWH60NJzVF09un98+mEMCit
XtSW2zn0q0ADIC9I6b8MFa+DxyfkJl7N0z86jIaPj8XlPA6KB4rcv+h7zGgK3kvudITLman5sPY3
XyUGJ1OsGwfKp+4fBv9jL7sQjQWOCjLKtFeAUCbl3vCX30+2ts+sz7kSQ8OI/IAwpOhZVo+/1pos
xNllWW6K+Lk2ZPRlasJELpvFfzCasWrMe65UYHYdMz+86d4oqhxS+HygPd4J3h5L3qUvPvwkdj02
98BJevZ4wMEqMASj0HtFttwo4yXM8ZzPT4YPsAA8UD9eViSiyzMt/QvVglrkRCWNnM96pmq+bOXG
XIX0WHdBugmM4xAIWR2PtjO3m310BpmNUWUcC/Ivw6vS4bTk8maTrvREzBnxF7y2sMLI1NHAFfsZ
n/683lXd4dCgD7hZ7eQgwuTom+CsTJrEpYA7hJmC2qpdCHCksxMyNW/XH3ryhxSVMSMMJkdqnnDu
ztKGdZ7nWzbz8T8YXZKtXKKUQvLvzA/rso7U2JYU2OluWxgavMrgDwwTVQN4n7sX2XMu5UPwm2B+
EsZQEj8ZQQJaM6MbVhymekiWju4ivECfydeEKVPQDyoHd1JEhZjGEn3Stwkmzgu/T9+kcU5B0PTs
yg/EMrYb2gPQ+mE7qgYZtCRW/bfad6V+yYrJ86E8sHjFTD4fhwonbivZ0kXzv9YrldDJbgntp2SM
oXqXYHINgEefzN7yP82lpP0EubJdBuq2iDTBOe/rDQ82TdodGHeke4itoToaIsWohQ4V8K3aJHSn
cM4gbOwxPRJ8JR/5aXmKMQHBCv9G5DcMQegSi70HHiX7Rn/Yf0alf3sRIr6SaDMwOUdH9w15QCuz
0SmF5WrQn3bwZXQmPP6O/Ja2RgpYd4ixBu3vbhy/spBfXeSH5iOdaH8FGKOE1B5yhmTbosez0F3L
3YMl5VmUNFH3AGMzjLpZ3iEUnZPBbyKdGYuQlHMaW8I7zNtdXjhjOxM4KnLTVNjDFsqzawibm0Xn
tdblxSMGoXwJ3gAAFNTtwuslaiAKPnXhRM/3Wj6TwtWCg0V0UcPqhaTh+VvnuRnk4rdKskj2Zs0T
KO1K/H19urxCGxB3L9D6LWtz5BfEOSzPngLxf1pinQu4ozJRn1jG4gOEcdE8OUjH2M9oibPpLKhE
Dy2HKwPENidwmrT1HGwUklc6IO7JhZoNp3KkUiyoXtHGy/RT8amugxHMah/ipsFvoq6ERVB50I3Y
1vr+IzoU2O4IQXH5HLNvSOw6qDA5aT2cJkh0vBbJgY9pisnNUyxAp2kXxah3R+Uw2C4KCGj95rm6
+5xCg+DwmCLO2A6haXqc42PRWiRo8fPh9OdBmkiTF1MX/EvGC/rKDoJkcJD7gSBaAbsvMmU4Rr0s
ceYAT/XKfxhSZMZMOs8PwEDVxllrmpF+iSKW9+XsZfZEiEDijs02ulhiQvT0B71o9TFEujnyT0UW
SA/y0Vhq/zQ9ByQD/UcHtOI63OUxJOl1vcw+q9uwzMrMlZAySPH2N2OcxUSwZU7YjLg65oDmw1pI
1Y7mwhMDybQEvR/PizHhIB21mzddcCu17m5apBlWhrL9R9MFcJRrpWbIdhoRAVfakwCFZy/ptZS4
akL/Z+TH4KdDrc/KQs+41SBi8Dj8laMb75uuTyi0qpaW1eCOWucNn9Zt5q0sfP1IRKhHT/tGONwH
O/vYDXvT8Jxk8oaWim3Tzbs9lVSdhOMR/8aDajDQDx9OWUYOH0Tp9LG6WRdu+lY8bMJ/lxNE5qgG
8otwAFe356KnPjaKiIbSNw/6TIZJPFRd2KiG0p1hTCeOyZExb0+qJ6Ixg2gzx/gbc2KD+iM1vHPG
5SaXpF3xK6PaBgEyN6TDVlRftYj+TGqkDjjdIWqn2AHAOVJZiJA0gk1z3Sv49gZDVcarxK0sKBjs
OCOyLPp7Lt5WIT1cWNFs419A121L1YDn+lnPExqsf9KTue4NT3Y6TAIEnMwmiTy1h8/acViRW04W
h5+uE2A3VYTtIqebGvRE4W6CW0qGors2ftZcztqBNOyg0VU33m3OmKGHbUVFzZ2VUhHyqvPEUwGt
37SyWmx1NU75xyts2iul6oWdsp7qKdrbygoSdNsW2aTLDLBwxjEOysvzHzr2E5Bn42uUsrFpBxZZ
D/Fzle3kRcNJ0Iz2XZAdRxTNZPbZIbhAfD2+xqpu0AtVVFFmimLzeW8GRlgUGUOk7szqZonR80pa
Vr2+1aHpZ9u9HSnjIfk9Q4nSguYw4OgCkzUE1AS9WO8y4KcE4mFNxShLn23V3Qkeyemmm7xKVsRe
1uJjgcGEr/J/Rj7UlmnJGy6IizUsH0tDbK6NKVO04vCExpehxCSXV9/6PtPE/8nvvB3WowmjQB9M
XBy7MdFn/slcKEn+EQuAeR2199aHNHlydHUVPxmO8piOfQIZnZr5rMl7jiE4vzu3O5sFhLUL8OrJ
u6h3/BfOPsYYgwpAeDc+Wb/HgfLZKBS22zA+1QIGiT6HfIt0Q9Oy5CBDjvdFVGPICe26bb4LxwVx
kj1UQf7k3lYIVynRr0rQTCQmBUlOqTPB1g0WMMnPjJKjjH4EdnNOZKNoZ3Ssb/+XDre/dDxgeoT0
W22AoBXUmVE5t+jsCq16i0PIUPdDBJEz0O79wHuGc40I6/mt95oHoaLI0wNW+7xQNRSVBGvc8lN6
1x2fK09QoJ8XX0Am11qfkwgQDiBOOtYyswrOSRykD/mSXZ30erNDz52y7WkPVjjSXveXxjt+eiHW
CnyYXGwiRONcv5YNSnYX//Xgy+BGkI0uJR5MEBDr1prC8JDUM7/X2NldjJbjf8YH8S1jJY13BQS2
M1Xxki/8I3Yxl7yemyqTe2R1THCsYT0ey6e3kPHgawnPFuxD0EnvBqCQ4WlivqbEePvOwA8aBGyr
PR0QkHyitC2uojbql7+ckq1DiCSMIUFTUJ8DMgZoN/QnwTngnauay4+5dEYUFBWZchBa5qsaXDC7
0bCV0mJTX6Oio66CGkjIUMSWYdoNhEDSUm06rheieKglOhrGmdoq4jwhxrzKDH1XrD6ajWvRcNBy
wqLw9D/8KKW1zMyWQiJZ1l9loHK1rkoC04y7e7znReBjbo4Aw3IagbiJy5xKMkP2Wr1iRBQURkGr
RS7m1xc49xZOd1TEkY1WANI9O386uQIpjbUJss4l39J1TRnWpLUrCZgwypMBjzxoYPR+IlSnc9Hm
X+dce72IyDxXm4SeB2ataB/gj+K9BpPTRGgnSoF7oywIi+++Ywm0+x0/tfv8DQMxbK9y+bTB9uVD
L6qhm+igZauLY64dI9kRB3NYM0QPBy4GNpKRMm4V19UeDc8BWdTzEDJHs3CutecTSFrqrnPknj0N
R6gojnzks9Ms6dVs81/kYJWhMrvJVjCiijW6Ms2YPaCHV8EYXVRPMqn/74f4VOEMnWUv8VGsMjvJ
GTRMaF8EBtu9GhGQUC0jAGIBrHbD8YcZ7L2pu0nAsYoQuSPyh3Nm3jeY0GQbF3mAbYdJ71DkRkqP
O8CfpeQZxEoNI7f7U64U0+qN4w8Rilwj7XSwCh3jkb4zurud5Eyv3JovBLpGUXE0ja4GxtMMUel3
Q38qOpVtijSy0OeK5bQ5wC+/bNFIkG/ZA+tFqKH3dk8MI5fHwO6QVEvq0WqyT3xXo72tZ7AbLdui
OU8GqxSU2lrhht76z5ZUEvoEnv9AyFJ002cdcYpT7CFNxeUsBzy25tuM+XGKiw7/k0M6b2JhHJ/D
/9+xGfwX3z2wQ3hWzKW0ogVB8TbATjH1HgoggKaShZflXSB1dV5uwh1kIrK+GaKkditK6WPmmO2h
G/JhQNEwAtBiVzvLcZnXv2w5plfYNAsINx6Xk1AW4oj8KlBewKIrWqJPJ14gJ3NFcKdu55kmdpVt
uF1FsOID1PziFng2rUUqlQgRLbpOecIgjPRhSp0dqbyeflUC3J/s7Ul2G2el2XzT/Qi0WIauqUOL
OZatLnZHtd5Ws0DtFpEtk6+26ovs8eT0THg3T5+0Vxm6z7AiSBKOQJUSmqM9V2DOIlgh0h5Ol8yl
ncNjxZUDSKvGW/PNfWMS8F8HBGWzRcCKO0ODNhZaZDprQLaZp1qcSVMICIWbU8hkuLuyahDgUfHs
p0+wWMMv8R3v6rwaFLKkGr8t/PBmyUNz+EX40JwcLOHqoaJbLY6BVcONpQ5NB7rrdYXwv8lhACr3
EgDeIY082yXZ9gUfvPfkHom+uUt9V9rhtvQpFmVRP+0HmdBDpIdn9HVqHiVCGfRjRX8zTErAB5yC
h3vfnY1RKjhA1B0trUj1LN02W6OzWNDwdWA2uTax4Tg5ubiZAeB30nYEP1K+kGXSmLxokYkICUHT
knwkt0UvXRq1hZw6T50qU3awcbrEodU8/6lH+1OmMv2wYk7Ppfl4Jk0WuuSO4uNl7aP2vq+MKBYG
vWl0seCowlJmfo7zUFbW2U7GeSutzc29VfDlffdlTwkSObBZ+ubbZ/vn10piJy1fhauESck/jD8r
UNAUZz+8uMLS1VVHtS6eKgA+tIFRrb6xVj3w99cmwNKMh68eMkTRDpVaLszMUZbPDC2J0S1uApuE
DcP6iD9s24H5JcToo9U4kuqMnttrw1T7FqsX7FpKlmGH9oJ7GCZB+VGbTksb0MPUnVhW2DvdtLv1
Cs4ByUeKD6dKd0Fx+oTmRKC9OQS7rvS8fw+KIX+/UTcrLLFVscCPCm08C1PKrV9IRj8Qf00llbP9
UhC9O8jVTKbmf6VfjttBC7HGssRPkGZ0nTxOKqSa2+c7cabYtunSB9e5ck/JD8r+l0scPl3jkLVK
cz3bAzmYOLZlguAj5zd5/Y+GIlBdT9Atrpu9sLC767J4cGDW/dnvZgqx/e4E4E1trjSEZGTx8AF8
mAMnXDqSguNuU4dNOa2Qp3DXp4OqlvC+RHnaJn6oH801ftDiSopw5+V6cF83I1vPknqwO6OlXGkc
VTkK22pTyF+qAeHTYc24PSdvK2LtRnqAEsYZ2y/nH6wWj7NVp9kFfLcF4WqhL9Nnp80/JUWaEwWe
yxr682IwbSUbuyza6x2mgV0uwaF+IZF35foAVVkBKkOHgX+B6LyKiQt3oCcQN8z35P+CbZPGzSBZ
5lx/KOfe50CqrYrgVkp+kCVsh7jSKSI1VEmgol4834tnpjcOVsl/+L8AMJOidNmlIi0ZJ6+vEDpE
ba9UGwiIa6+S4NTlPJ2G+g7PvkrnC4c2y6rq+nH8506IVwaeeJm01Dl8F5NSIBynxhtZeL+HZnIZ
bwKtQT070RpyVZqCs3T6wZBrx5Qlc4qUo3aHup+ICrXsliwGIGnn7BfBrQ9YYXYIFgr228xZnn5b
4g0X6rx9cE6slqgL/rgY+WRWpRpcAIJmQGJotq9S04HPn9siSzAnJ1hxBfVtNdf381le4ewOjIuQ
ptG3g6Ey6RZ4/buMBf3+u19TOm+Q9Q1lAGYrQbvUu76NESwVhOwX9o03qVz9FRNhGNgTgpYGJ+E3
7r6GG6DEJOeDWGkRm67yS1jAWUfyZfTzIK0IDtEnri4tf+h7u7iKWCtBceXj8OqziwTQGPR+GIse
xgziVeX4/7xOpKjjE5a14ac+qJbNM6p+CuyuuVth3UL5TJFn7wVL6ExW8HrYVHgyj65cdgN3LJlS
2M2LPzH+naMBoJdvJlkzivvytWEm2ju9A4/wR7e/HP+l4+nL9M4hEPdHlozi68TQ8QJZd2gonet2
FBscZiDeNy8MtMjOobydWdJjfyRUcpcAZU6Bve843wBCzsP5te4+mUYNu+JhTb0DXKvasEwmGFHD
hkkSR+My9INGElAcCTnOnJca0pDWRapdLWBA+6iHf4o9CBkRv0+4fQccCEEHLtI0gWndkMyxwHho
wnPbl4QjdkaDVD3qmaEm2JT6tjUpuonXeotQNB8fPDCCWTdCRkTp70AlL6Mx628BjnIw9OIVt38J
Vnf7qvzrQJpv4+ARVnbyzW8hUuz1nV1Zyqo5Dx0Vi+b0URBPil/egQH94/SnuRJBuTfQ7v2b0UPa
MP96LjdSxrlp/7dqwBuRaptn3MmGadn7YhLNDp1+EswpUUoGuOSvZd05T/N5T4ZOa3rK7G+xdDjw
oQ7NfLTlvrWnKXyA+ta9eWTm8ReqO1XtpsEE7Oz0Jm9BL1/AaTBKXZrqBxpF8HhLY5HF5y1rJbx5
UheFkk1a8p105T3ZHp3vgjea6+ZaqfDbL86NvVIL46K3yvlJNa1UCQRigoqOjBoWH5xHBiuQ7YSs
2kY7xz0He/W+s/kJ92cCigoIHFX/fSZ3AFNZ+fc3eM6m6HXo/R0pqUz5D16wSJjSYfikWn/So23G
xdxqpd3A+8crwxpHfmr6adplYifE1LAyj0Yx38kDOto1jru51ptCrlKCMm/ooyDoUo/nHUOF+Qkl
x1szC6KAJ7hmZa+kkhkB+RP0U70/bi1cQiuNcxxg5WHRt2YyOi5clZQaXTkeg6HsZUUZ25fOLlNK
4mAWSOAEMAYRAGb5EFA0zfI7ou6QN650H4w4bf8lPB2RNimw3qx2T6P3ndwD8CBa9qftKUrMf97w
Rz219dwD5bnPAPvabhpr3pCnvMGzqTOS9IY6ytrJ1tx9yx9JOzwUIkqMpIn4zIRMFBQqRyGcbwnR
1+65ioO2dXKtol04h83oTCI7mvMm+N0K7E8umYYMqhnKb+EiYkDY0A9wcDnIs4+Z2hX+viIlPlRe
LzdpB88OBaoOQ4JiY0TOPty7ShoZ9fjEAQ+TXsZ8jwI69HLqkd4YO3vKNYEeRJ6NaqrKwDHIUP8G
IjB7umtVDQ+bJWFvp5GK1v2fZFa6mV2KO9VnX4eUR5hnM6y6eKgQWYAqpO2ErzW9xlgCs+onDF0Q
8WKjSu592bo64riRt+Y27OxW593+QKQ3F1fCVNNdC6Oioes3bxgH9sQqX0XGQka+R+o6z5umeG/c
anodG5GxwC8Dlr2QIaPzACjzfkRir/zLmAG3qmZUDJ93vXu6kuXgOYZ4+/mHMmJjh+AVTC6mxd5c
TK0CVyZnJ83GNTHlseoqSJ3ngYGFSLqFokqd9yGcJORylGD5KAqatcXVYw+F+lbNEmg1y0P+M+3n
sGpxLxec7FuyNI7GzcBB2esDwUD8ek8wj+3VC2m35L8eM8yX9o5FFhQsgaRFdfbK/5xlNT9QLz1X
nhUqs75jhZwySqZ6oVbrHzTFpNDlzlKFlBV3gs39BsGuZmPynw6FCSumT9Qdtsd7WzjUcrKvDJLP
OF/RWnj9I7YG489MbF5uYxlj24Gib6xtdcTVOKfS5TcZkEXwD2Xy6RG8IaWQKO7uvhCcWY/QbRV9
xDbekVKhfu5xBIx9//eawbpmyyg9mw/9FgoimVnljtcF59lMREklMW+B2qAz5kUO+7k0PcVHj3Rr
M4yMHcfv/CeGmTswCFZ65rhfIjumSUXSDKzAIOcGEweg5zntgHRUqTMGwXrCBIACOv4zHpwGUi92
3LH7381ZeL0lzHT6DF3wIYfpNKnEK9jnoza+/OGhsRq+JWVH8/8EdgAsibqrRCK67Kp61HlxN8Lm
v8bm5GsHZXcv3uVrc1UNTuMcHWIgbp952kpzdvlbNRhRsTFTN+pYupXYsJ95JXaMOHfrA3qsRAZp
pXh4Zh0jEAjMTPsCpQSfXHI9QjxPo53QQMdxcfL9ZjE6iHS7DzX58AZdK2ldZUm6/j8UNVIYxbNu
a8BCsX0iQLgOrVJtQ/uWJMqvgFYOAvFUbnXI60kbx+U49TEmRXNlAdDzLusiybor/kB4H/TJdU3G
pVOP9suvKYhdZntJ0J0ZgK5dvmDHLKK/E6l0bIpNZgsmhGydmmg9WtSN+OmRhiAu7HO6qnVno39M
HXFimu8QSQp3/7TjToqtks68TuL7j0HbAmoaUFjelSXDJzZ1rh5cS5Rdc3EYyQfrN7mOdTlvZPzM
OhsDHz5+4Pt0Razxk2EdODsjUEkmKvPIrCJZ0eTjndh7mXtvdBE5oqU98U/4YFhrCknZ0gCCPEpN
ZUcMQH39AnkUj4Rvmgxrnl8j3honR143yZ/iuYAtEewcZvlbyo0b920V+O0wO7yVb9f8hjAfrdqj
tp0/gcyJcvY25Zo7Qs/fQu3QyXq6LF0CmlAF3/9RuHy9WGpjUkDAb/xjLY2Z5UPRDXhP9Hj+aFUl
kQMd/5oNhPBzIAOuFVE4RzvZ4WSewlp9+xjLnX6PZ4iybOS9bnANaZpaJ3PqIs8NRtghU4rpFmt1
e5ycej0yvpISHx+u4SPxhNdWCNZAQvsngSgI+tpMsldRwFNYNbdWttG6m1Epm2WNjM/CK/7+lwFb
I8jR/56OA1eN9FrKsrJlfO/ywf0ZVLl732byGwld9v4XkODgxbMNFQu42oT9ooyctieS6vpiPdhm
hpL9OyTOEIQ/G/gL+JC7BiYB3XlhpUff7FEUBq9b5YkQxWTmla0bctv/4lNQsQY6otgRO0G6Urh2
S415QpArt2nD5A6bKPa1WAntSvQI9HqVRmaZY4NIuRtP4v3KiSbQ5xsVXKWQslGPQrMhBEskWAjb
XIIlKP/Cnc2fMm9EAIBdJ5qZ1hhYxn9JvxfBznsnfvIAcb/EzupcErn7Ueq6PNEHDDPMgB20Q5bH
51N4NdMeMTXSkvH0IwRzRfLq3hnB+WZq5ubYFQuDmU1QCz+A47+PwMIzNJLNTS4Dj6WNc6Q4TjKT
f0t2USiop5zVxCTLj7psGu1VusbATG8Ug4sR7K9UnxzdcBIjYliEBBZrQWoBoWbasHJzR/VuNgtT
MUK3k/koQZr1FYiHaVYF8piM7h50wC3aAgjtvIhVY9Cg4vsZhVgzvyqG7s+V5NtJ0Suqx8scTsc2
eze//bEYWVYi457/zoGhOFVa7JUg+TiKjfDxTsb+tPAjvQa/Ud/PPKEKHOrR4YSZ450qHudJ75di
exYYdBLDuEojpIirEp0Zo0P61mg4gqwy3Qw/6RIrFnmuGmgag7NYPp9xDRxlkrqewcBTiPzAYU+K
zP8kPuVu1xTEKZ183BSyoh5s3lVfqo6M/+z5u4Mjr+xxjLEwczPC/nJ5UTXlIM4Ea8a8pMJ5HvZ0
yneQCzJm0bCEomxxmsfmQZ9f6E5JIwQy0jQAmdUCTJiW3iF6s8+TP5nDEU1OTuHmYF1yOq4oBUI4
35HBZU3c0YrMMaRZRF3J+YuWrGGMI0FjB6dDva/nxVQCegnFLI26kdShAT+pwbgO6xoZ4IAEXJVv
Ou8Qo4NSyZUKGPCqY7hLdZpYp3L21sa2cbKoHdeRVU8E6CNsIr3p3xSzrFIPxIVt0QGW7IYI+Raf
cS1ZHj0WzGKTqjJzi+o5XMyWgEPJvlgJAQyh4sGpE6+IqbMav6ZkRFgtXPDsa21YjUD45aLXGvq7
eU6GyiM2jyVism8EUo7/SMw1uxBT02GWETPCktmqrN1xgDUF/9gHlVfQNekQCiG0JDmvf1zA+s6u
QLlxRQkn9XG5yvtDWoXRShSzBZEuT5VG8e8Af3ORcQv1D6dYm8jxPcKwsoKRZIEAtKCN9J2Uo+99
Um7pDJszdkgmMAN2MWFdsrB/guGYexBnS90V3AX4bCswyAi3EQ3VZOYjVSIvxAQ2eybcLDRcihgU
1UIzTPj6Rb2ueLAYoYeLq3PAbnycq6ClUaoI5VsRFRc4kgdsQheDbIwlOsP52I3Kf+vohNaiNYy7
Ww262dd2JuOQD9lX+kcPlG2OfBybsx5T8mktLDrWZYB4UF0DoE0F5CNIJQEqSff68X9G+nEOvXuu
Q7JPAes5y3HLtyoIke/JRcxknPMkmNQCRhxh/dUz7ZQsuoAtqBrqeH+p3WYvepQRcwmfxx498hM0
MCedbUWAEkbuu4xXTEc8l9UQGkPK9XGpxGZ6h2YyQd0J8W8FkcVECrXD+h8wdZRPHBniIHMH+PCW
3z7Et9IAdR4bAqU33Qe5hzfpHEhEXNOM+2e4+Nl2+knfjeR9hdG7/Jiae+iKr4L/J09s5U32UuVW
DEPrD+J+uPQdJaTDng3chfpivCQXVrdM574rY3v5LG0JHs4rz4LjYV+Kb7QFl/1pKcSjfLuxf3Tc
0NxXfmI1HmBg3Up2DC/NSfgL4IjLp7uaaAdMpqxCoCPdgFbEgcE2yS4EAR1sDXP4KEtS3pOQ1Pqa
jd1t9y7R8AZVATvF0+jeKm9G9mO/Fy9exYh8lMyq0iraTSDyW0n9TOHDgtvEqo6I3MWUStiMadVB
ekKIGX4J64Ge7wIgy6Stg2vZ3vTRX7odC5FrleAMHiJjHZjI+/a+jY3paQPx//ghTiAVwAoy9OsM
mQjyPgJep+YY6UuvHDdl4DCmkwc76bGyTvyCnHTMhujBZnqvfoas4WrTLk15XLRw4KHyA3w5A8eC
W9Ud8u0ohJ9ohiand5f5MxlqyTGbiJ4IZiGq4cZcpXvbkCcWDmYyCk1pBQ5B+5KEsaaFmBF3G94A
zf5QRLApEHZxcJ8/KXRck1R6WQHmyqg09VKVOVllRHO5Eb2UmvB8ow1HZQL79/HEnMRkteeT1cvO
bJRFdq5lcRKaVy/YMoGe3rg/2M0hidzLg8MtkSri2KhosDMtdJRIRigF3gE7rHR7XjnXRXhEigEd
zvi1QmYSOUriAKQsUDj1XZBfhbJmp8lAmnd5lYpi1Q+r9UhXwquRnwK5UEUXCpiPdQEaXETyuRg5
kL/UZChqgoXbFxFa7Pkuxd8Yo++yzlDa15g/HA0Lll71wUUTrSDiTbfr+c2wj3bDxx3NaKgzfxK0
2iNcsggEb6bPVrlMizfcVauzU6qh+VFtFE9lGq3SNpJelDy9vVWqohVNd3xFOQovYc9vfNjUlMvC
ogoEPWKxXJprQpHUnpe4P20YxNoqFpM/0N46im8AOg4Jtqvb2bJaXFtu6MG78elBhqL6vA3JoPFx
na1DX3u42ByBV/Xa8EioVdxPxHNpkJcqLemi6VB75odo1ho5sBdVCke4Ye2H4TMb1LOP6vUtvZR1
f3GXfV2liLh8cHDV8kRgZla6DrWLy66iDmKIaVQRXdqw58APb2c1rchVvayShhmoz+D6viswJrUv
VS5qKRhQRyjkED79RRvJchw+O5FVyFewWYD6SLjLCSbeFqXvcUIxoqryIv/sjIlZFjcpAxq0UeEF
5wBu6agHyfXkDpW4sg0Cc/9kA7XBo5cb8ewoPr32lyLvxeYJThY/29HILXnup+AuC07aA26yMDUI
Dcsj+rz0Qsa/K9Ysh0FmuEAi2GvqzeR494hSFKqImfTj+eodbyARBUkiTNzZm0wxO+vNxzRoRhnU
2ehgoH0h2r4WAuW3SsE038O0wAnEv3z1jsObgKzrH9Z6fUjE920PRZ6xkVd6yPNjR+eIbTIYWeKa
1qHl865Ha8D8H2ZqgpiMWHCZuz2W5crp2/rTw2Nu0Z5AATVnDCW9X8z1JMEJMNuyjo/+IexxXYkT
Aw2kP7w7j8wo/UqKVGsqWBmbwgDYp8Lqvjuc0B/aQGqxNHD2XBz1WeyiJdl0MFAq0t4yt87SYKpj
x3+CqbvVCPTIREUBX/WnlcgJzknA/mWEu96pb6/mfVLEEybQBYdb/IuG/vLY5KzRHJ7QP6ZAQfvV
rGtliihMjh7wGQBgFjh9vrO1pFzxAMvwfp2QwEqfQRSsbuC1e2EMkBftWWHzUZlNYx9AhdxxlwJV
g375bPfa2CvQ0S1gXXlmBRPobo8RrWQyKE6HB4S9qzaUbfZkDO/Bp1rJH19eeGOKyZyy26UCOmY/
QJgaWhWk1jeUyeSnAcSTayTGrF1cuix8HfRQL1agD8Loa0jeCtYe61FUqXchF/Bt84MFIN1jxBLR
PNuAmrB1wcMbumRuzRT9cOj13Zp7vrm7PMRPtZk6/qK9y0vNVn7wjIbYVusQ0mhQuR8+VQWTgv/5
CMnJ2LuKJJ1shSCsZXiV+YmYe4/urUnMEB5hrqWlQ5smtoXsYvW9vWJXv+gSlS9ZC7jae3uljSgS
6GxJcVld7L+49kUQH4FlcQIm8JGiXyZ1EQDIZe11v1wSg2bZQE6CH2aBGNLwfnuzbLy1TvcjY8Mt
lxMgSn9X2AXdvI08R+l6E0eDfhzadtQfTE67FQhPV3k7dEoUQbFRqNlWvJlegTZyzII8kd+UIe1J
154jwV0RbSMNJrG0GdBf2d/GPSmFJpNyPpdAz1KAayjWlujdnIUOafFXMe3m8jVFj2h8lEs//eAH
e3lf47yiysBZGbSghwzd+QcID7OLKyViLCuGjCd7UCCofH/TxIjZbBHr1xjbEOAAgGbiknWEMOiC
/XEJQCeoNZ9RmFtyJlQCuBbBBuS2O0vc1h7GrM39i/lZeeins9Gd3czs6JG1+L49dpmOc2m8D3Bl
TnLoAthpOHJh77cwWq1mrc+8u2zemahp+W3sgqyF9WrqSCCzhrpX4MKrWKIqlzxvYUaw8ISEZZvP
PPFWM8hpaAafFq/RgtfbO5IHDl6XMw4hOAi/R3GoQ1YoMxyT56cOsGgEcudvt2KV/qD5CUlS302t
DEivAoe2412fi6l9KH1C7MJmBhNqQF0t78hMZWGmRqgu++bvducjmX8NR2tfbYPQvzW/RNJyUR45
oPUmWC2MSC83xQg7zR0UCBlNdSS5ulky5pwG40++nCwGsI1Z/ogaOpJkjg/C5bjqB7bejrbpCB9o
0eeOL8MUx8qGsPavikihTPaNBlwdbKVHGmVFkTMUIjBnDSASfdGBlfwj1KDq3vP5v4uHd8Yg+P3u
iBzBFa5C/vq2vqSrO5jwwyFh5Hxgr7p2UPR7D9DeNgKGJRKQc0XHaOkJP+GJo+KSACCGYaYFgFV8
dlIkitamSFhSZBRbgrJFKntOQ3Rig1bluHLuy3S26j0Tsaiykno+ABM5Zp3Qiek7dWqoDatKbQR/
xDCI7yIr19pXRpM7EXxO5o5P9rGtct2P4vM53WMtBuVkQ4nHrRkl3Cg8z+S1YRrkL9ikYHczvou4
EF3BqVAL2Yu2kYA1zHcZhS5RxcggvzM9HHryYRKTpKaisOxWf0dvG3WnMrguyoIEOEzuAp+iXoGb
hfXccACeVEpQxtrweTYBU0/BaqOrX+h5RFn80EPHkN/kpROGkHa2cc2iHKyqoMVeSKXa8twbopeU
ut794kKRIyNKhuG9TenHXXijBduU9t6dkx7XRnvhchC+vgVVxXu1EyBVpY1kcVxPc/g7ur5u2Dp4
3nkXCRKKyxUv5Sw0kI8l9v0iuMH6hv8esIEAWy9e9PUs3eR2qGU9N/GbU9mo//2bZfyjpxIte3us
fA/RK8LXddK5Lb1Q7XUMPJSiIZbFr8kT9zP1skKQjGw22Qm88E+nDsBZBTqW/PXhDIRhN/1GURpH
/kaf0vAyWhKtTouOAEo4bmoKlWxhuh6pq+CCsSuFAmRoAGURCA1rljekGDEq6byOyBlQr4Fp9qij
TFbtDoeFOc5aVypIau8Dia1481Y6/zYuWEKo45qvSNjF/cabbnasGcjtbJK5/Ha+930UUbfs4JbZ
vEDEwE/cQkoY960xvHltYMCEkcJNzUXIfjDv2ERVpYxpl+Jm23YnkJ/IvaPYsmY1AdrOLr2SX2Wb
CiSHQvbBWYqgQ9KchlQxu32JGvLL5jekgWcOeP3Jlm0097nxuPkO6XhkuJNALIbQK7fxyIk7cR4B
f9xLgUu4PUTzupEle6QbOBLn5bklViUvfF6auH9Xo693zl2UfTXBuGzptsucz//4brTCOQy2tbBr
unhxOpleJpCh9ciEoSN+Sk62mnpuwdMWEIDpQgZtIAl8lCEjEJW3/8/FGy+55NHDzm/D6Y+sohe1
pL0Bf59mFW4q3H5aggfLDinNKGneVNuCRnyZAntB6KijGDCQwnFdV0xE6gyoDg1xMD+d/anIWAJx
XhaPnBSiHjfWWRfvBW7SuUdrLT6Mu9DTgYJCWxrlB6hLKbgWFoG+emcmeeUPeLjpgu8X342XKlpd
8Y6evKRrXuSDoZI1RyKPR21sCKRgCqjo1qshvevDgA/vVCa0qZEJxw+TXFHZoUM2fpNYRn+SP/bh
YnFVvf3ykxmEEuxKws1r+awMiZ6dpirS/XXSPfX5JqNADXc+hupZNOa+UJJm0V4/kZ1i5j4fIA6j
VLawyI4uMIiCLKj9vOU+9lN7RQ+JoKHIIp9YTCqx9DpMV5cvvnPVcShhiYL4cKRBJraQ3ofmj+jg
5PvWKYY2fO1yY4zhQlSbZJPrQ2/+WaatBprVz438s5+6yOV5+AjygUORQdxtD1WorXksapoYcgZE
majZ5ZrRV4E220Pa3h0dpJM5tpNhmkUyh2xV0/e67jbePdayzKDDFrbyiGa5zSQNUdbg4oKH9RB3
uA17TfRQNnSnDHONAc884TpvRZ7A04n7qOsgZxg4qjW/kfrhqNUHCd/fIQ1ZnbsgoliGwCskoQ2p
GhIRK+QAqYfLcuBdxl8yGhLOE+hQ8LPZJClMznceG4VTo7VvdaYr2KSeOW5+DWuA9L1YKlaIyg40
E7yUGRTEHOjZD/Xbi6fJCKX6j9Sihh1oTnK+RZDDM2inKcOCifZkH6YtlWAWdYKJjL0QMPbxs42Y
ZrVy1xvtikybtpGxvl6cNPW/X0/DrsFcwM+BxXEelVTsQHTqmsQbXIqUiU9e7CMIoqxQVmGls66p
0LKNKVELLEOahpDhal3dubjCbvINbg8j412Czx9LMrIaOoWimR85rWjso3CE/j6jcGj6II7SsJtJ
PL5hEOVZ9fzFPJnLs5TBAtNq3r/4DKjqID0MtnG6HYlaktyLgpZcOTwJJw3B1UF+n90AKtdJp34v
W/cq9f1hhpAY5Dr1GYp0MtKlVGmV16gfQ8YD1EUFHXRSdwZqXku/Ig/SryOSmjHU0xhcG6+Rm6Xd
K3xfskptWvZ530tdl8Dl2a3/3VJj2ZDjJmptCXoW5bUA+qKLIhvjOWmYHfaNXAlMIw5bk+c+GOfg
q25gZ8mTXHV7yvRnX+HTTeIdyXlvpbjr9eS6rtnOyn+Kw/sNzm4EnaznvczZGqRxoOlfPq5Qaqkj
YA63U04abTvOPfDHqT9bFkpF5VaFNp30ErtjDxYNnl4PBm2VmuzYe1CBTgwbp3bbpKvVNa76YaRX
ruBADnKrRsaZD9CQi7Hr7PhY/brj1Sl/Wo/AkkMyjcP3uNBdHSXtsdcWzv9gSPtZ3LcCZQLh4r/a
x4V2nX1T6Hh1+YYfZYaswpoPAPzkhd/up97F7ed5DxfvzngGdYD4NTi6XQqd7LeqnsFsgggkMQGF
CDPlMvRrZH5T3EJu0jOGJ2z43lJkxzGTFIAhjF4b6/T90ZmZWz2eDfO+EhxcAzFj5QbqND4m0M0S
gTI9j45jhHgR4IL1Cip90DIV5c0w2SrTy8413Ha+hsnHDbk6/6/SRQQ80TCE0ROj6tt2gHjCzEZV
rHpDpQg5ed33BL+8SmqkCJ11ALIqmEDH3qFm6/iBH0dHG3TJ8peHwAT00CCFlbTyBks96yoNznYZ
VajiGjva6k8dlLONOTDPemvW5YlAANIZasWfF+66m8gWYokb3EnU2ARDFDxzZ/wYHKIUxhJSGwfW
GVQpHLJjwlOCi75FxgGYHgngrLI2FmbjjUMuzB6dgDOu9RvD7uE9a9mk3Jm/46xjaCwY4lIG6hAy
TgqB6VhDUsvOHEC8XqYnqcOpMUnd0NztIKjZn1QoKruekvur18FP5rRVy+27A4O4l0Vou1LtZ5rC
ocDBJ+SrSBA+j+DH/+iHwPvJKrL+KLlbFPBtd2sAGJ+KFHfa6CyjztuHJYfrCN/vZdaSQFvxtmBL
h1O8U/Xs2SIy4WhYFWxYlBTzS5O/9eukgHhTkzmgeG6hfjn8ZGGxuqSU3kKUWIGf9U3mm9U03Iun
qaAT3pVQv33FdRslIy8tSlZqQ/OLg1Q7r9oRJmOg/n5Di5np1p6MPgqEUAupC5JvZBweMHrqP48P
CHj0HyNoIsMYCmdnR9pLwUmsqu/xt/BkQwNY5P+suGAjgPCzM4DQYbkME0NSIoVhX6BmVL+lrcJ4
E0e0sXXS76Pjwiy3bpt0vwZhlGqMNF0LmoEukCaNYV9C2wMnRbekABnGv4uCQGWS5rhwJ/LBJJF4
DSKDYIoi4nRD6DTyoqPBM2bHTzHXOXv3qV7VGKgYi+n118o5RnBflH/aahScG2WLa+sVasahLT7r
sUAREDUOdL9x5neduwwqznZEREzhu6khzmg7HE12ZJet9OiHst+Tem+ro8VSOd6y0UffTGFGy2bJ
6VwSZwRRnl4QquC0Qrp39gNPws5SDzrOm4Cjh82NUWRde7wN58984dD/UlVnKgaYK2XeT7Bl1l/O
9Kuv637m5osEuV9o6ssIoMW1XZkA5CoREMgqJZAq1JReIH5lzB1Nt3ZQUXmkx3o9MKZqfPJn++sx
YLrHqjy0lq0OPuWmNep4dqkkqQA0kN9gw0007EDOmCrlAdgscfC05iUuWn0Mjf5k5VCuzlt4gEFx
9j73rCPIYmQpu0127fJrf+UKNZZf3Hc6WaxTFWKWE/04aZAclzCrPJGLzIli0LmVtT8qxhs6L8vK
RbYoQnB8A4/ZfJ8mcArSJI8RTn5SieIHg4xbUOjv+OdFDtMcrTRWx61rL7ISzYbv4pvguzb3Ygjr
0tw7ZisWeafK7n8oR2ciVXaaNDcOWwyZpju+sKglB+431S61Spe3JLZRgHeIZqpiZ20KGPBzn849
ywRy5pXZxij1jiGLTCyJJbC+nqxf52O/FJHDTgRfe4iN/U9yQXBT8RVeCloD6KMihok9ecp4gy+8
7E//NqzF8WiIChyKTtv/xjhmDYMmOcqanSreSJqPBqF6zEUkOGHjHnLYLVx8340WQ24IcJULySrV
FYkD2BoYSmfKS6BEJf8PkIMpWhuv2CAmD2PKaXdCZ8K5pfw5QshMhRA+FOORIDwhL6N3gkgn5ns5
cynpnBUbtNgSouemscCr3SQgkQOmEP8FNwAWXhdjTD5zK69Ea33jgJ/mOdjIyPUjO72vM7g5XJu/
o02gzzQXTH3zuTdX9zYKuhRxJ8ZotN7vazgs1TgshXK80n00hqPHBzW3rtj7g9AWfSYPdxH6xoik
7wUOsjguLmgygsRd2O6uTA8ZFVCoYKlISa/pHHc0cO4Qdi5P1L/ACg1GmsPM4F0Uv9ezjMwWJJsY
uPoE4POuK9dnSINSjJIq916F4cmr07QNHlC5EF4NPqozU8w8WmHAg2G+5ws6F+eNNnoBjSU7Vd48
8lQ3NHAE1J8HOZUNkMiJMX73zNEbEoRAGP9lHg4jQPjABbprhkv0IjWSAzR40a6OA1v6O8uKkfa/
tHfTQqKhF30O5tHVm6/c33yD8CDkDsZUlUL7D18GS+zwBbrZ/pObFD5tw3b9/ORSNM5YLrpuq5jJ
Pg18Fywr1nsFLBnc8X8p3wW8VTC+hvf7HhIRMy9+KjI9WvTW2eAfFrVtzlqLGr/OKXZ2rlqWZe/U
o/jZlfhm0sj5ESqbwmogcKUALx6Apsc3d7ivVvQK3hCfFzE0OhlbBgtmzI/WB4EB/22c4JaDzuo3
pMquWb5RYaJl6Ru25snPjkRWS/uw84cmuhvVbBzskbqNgfMSxS0bJkJJuvBuqg+geD2+5NK+bu7H
By/O+bEHCi47sEz4oeMeD+QvtckPPUbwqBwq60kt8F56VBtQl4oBKfuCx8m175BKn1DrqLQG/A4E
87XsFTwdpAw6ae3kK3iP0eMHf0fauTne5n5pOVPaujLvkQAJpo6M1ndWNJT8KXN2WxqM/ZYFlL9B
orYOrTqKAnou6sVFjH50x1AfDJQxcu48X5sj+trne+Tj/vFGZ8pFvNSOKUKWqS3XYZFQ7yiRor0q
M5nW94E60ksq/kvbZ52HLGJuViAl4R8WhKphE6JChB4FdrhfW5JkWKhUTdP7NobmuWOEJCvW8E4f
a2aS1X8fjNwj8UR/qEp/D8S6dh1/O3sjJn/90GhpsicKYWU3oL0SyR+BtprTCXuNHgbV8b8YR6BU
ExakbN6gm5FhDaCVKuKiaKyvTVQOEu/7l6htcq7BjcX8EvRmPlJ6PKduzDdyQfxwUGBQgpAPbEp1
B391yQNvKPt6oE+QN+DPtAphg9qOhob0wPYAzxq88IOubR4O0XbeKsISQ0zR4x3Pom0GqJA1h0jb
j15Q+DHFybvLZ/3qzNM6wzHw6FrbMSw1HNJJDUBpTTQCgj5rBkS9wRhGnOKxChG9cs/3lBDE47kA
ipRMH8lS5b6ZHGBuYQe5yG5laqtt5V79XPIhVpGFHJIEgWb7IRRdPwHK+34HkKnDsmBWEqG+Wfh3
igQAMEHYmR7U5KLZDmTzUP8QA9CfoEeBXy4PmWqoZfoFDhlpkYAqnJZtY2gF0bk0sQhaogQn/ZJT
ClI+6GfybB2MtVPwikFBkxywzhzfI/9cXEqKcH+AQLaAfRfQ0K9Cc0fhvTKlDbcDPJ1IHih0QDrW
sm80MA5ySvh4NmxvzWsXAq+lEJSHuvaJWUkIg2W7rZITrZZ5D7s0bXg1Uc1nR36X4AaWH2Ctkhj8
UBC4BnJdPO96YAbNKFQ9kllbeAfnaVTRLf3xbGjNtazPJ0vOKv4Be3QeSdumifmRvfC81N/UIf91
U47jzPstRyYwaCZqPZTP8w2gHIoKeqdOwx1/uYm6pM40BlnzcYft2iPu7Wf8MARQ758E32iGpeJs
qNbqmDNqNKmn2c4WzmWngUr/9jZGuX06xqyH8IC04DSsdb/ziUPVTjgIcly8+xkgMr3QG0JSrZ9Y
VTj1aZaU0DVsaHng993kAidKjo5sDk4FDMmREguiyuRGJcqQvtJfufwSB5enwq3VdIfAPvg3/lZn
aUlhvTe61rZRJ8gXcXqEu5t/JRr4eaYOvqoAFnvPLwnf+bGf51XPEMCYQee4CpGw3u57pvO5ADx1
pzBoZGGM2NJW0bLCAGj/lZQsy4A3DxBIsKn18mMb8SLIrqLBpN6NO0ViNrUW1Qwz5u0fVeLJfnum
CXYQgHtyPh4C4cAAFoh24OjXiAuomLyKQHmXfU65HIx25vKgQq7xj2A5Llbdu7ILaUYzt/ULGSXA
+2DIEBR4jhR2L1gbVHjNncoj9Nt11yB7byRoGWgIAFm69BGR6Ck4fZgjfbe5HBywMrZzznsllIRj
t/sq328kJFpQoGA1Pnr5B284A3E/jigBfcxm/3EvojDTfn3Bl0/i0cctcZ0fjRUDMTnjYnZklBZu
OySpPR3J516rW21lTn9R6yV+/uULPcyqI7afwfrfTM620JSstrS4YaGw0m46vf/IwTXXwqx6alRN
k6k7bz+FhVGI7yTLdqE3h4TbtgjF7aht4lb1M5E+OtBIgYJjdv6JUd8uAomq2+0wlX2lYkruA5HM
OeVmknmNpAoVhyD7irEqTlTF+bD2w9mYM/qc7BFn8aqeDu9mMYpxJgcVEHiqVL2NfAaExarbJlBN
kjs9hpMrqKleImyqxcSkoXf4Hw59i59HzBoqrVPqbSIX/Fzqp1u0htmVhZTNm4sm3itTFFWUO/mk
OLjuvF8fPVj/C+Wa9DbbA6G5uRiqDRDzbTiu240g+1qrrYLma4M4qahCXhThBQVBd/v/M2C1FeVQ
n6c5yFxixyTeZ5buUj5CXZzVfJ3F3EmDg2Amcg0YuWshm8mwt2lctUjI3dOkybIoApgxrfyNfUa1
R7UJCRtVXkd3TNyATEmW5+92Vy6/lQdwPTiaRI5nM6b41QeAGLXsPO8/ETuSNkE23IAGPPf0fPeS
94jRCRGF+7reT+YCw4m+ycQeB1WH7wycf/O4Bj0fRy2xiUKqTnmx6bufv8vgz3VzTQ7BVb+/zMII
OYl8TUKCPiKdPu9g6knQu/QlEKO5qyBi4uEnZywB+TlNuENQzC+ijM+yLtfnCX3q5GyHvNWsM6HT
R5m9eMulpkUNIlEK29RY/oZ8SLnOniIeMvQzMSuPZEhlq8ZppXm1XRBOZAv0j+9lUfRPt5B9s9xD
9BTU8A81kLA33XJajatdMaF4XAXVL3gaTtlTL/uA7Ls6XhOOG3Uyp378fN+1A7N32FuJXT2pBde2
tGFEULFV0s05mCBEWgZgy/3gfcfkOp6pK67DAnOFkNVrd7iX1DvBGHBrx2mVU1ZtA8mra8hmsagM
eTAMAJMPQZoIW4HXu4i+BXQjU6bFyfYFfB6bR48Pz7/T71asxPlIRJbmVJ413/7mBFaifXJJHSIM
Vt5ip1hB4SDlnpzBkh3OODYNdOUbQXQ2mve68GZwdDoV+zWEF+jVAI+ucu6Y6y2vmYOuqRSTaJNs
XCnPIYHbwojCJzrH3+htnSAxQCRuYMgZEORJ9shAz1RBC01ZOfPCNG1taP1/pphhxqtNvmysF/7I
37I1YAnei2g5cEEzuWvlVgBs9rnDSWe6GGR4eQFlbt4b1l6HtnC64tyeecirfOKkodXp11AFSV7E
aP4Z7KCz3TAG5n/SHGCkWxTwF55Zlg9fZCd+TKX9xPyTQ+z37aBfo2HwykJGgCaOCRSZqQ8WuiQ5
gXJbe9pTkbznU8BzcU7rDchST8yiZjZNR8PeJPnz4EfQSNKKhgCDeyjsGK9m4a+AqJn3dDotM6kl
L8dP8BLahH0DFUm46/wy1DGokqLkHbRKDadHk/u07fnbkb/rx1s/8cjD7erYSL3jvhYoAmlZEBpT
Z3gyRXKfgR0yp+SapO3vNnPoLJ3Lmff32XCVBFnTeoHFOZZenF5fISpIcu7n/940ahUpGFlZwMXU
dJEHQF0W0Hgk3Qy9hm956ptJkB4t7l+vtbUDPHvBUXhaWjnaeTjKroBIE8Whz7u8VrjagROVxKz6
V1Wr6ZbbZLvKZWB1x+kGh8HLrWhFC6eNst0zqydtsGYB7AhhhjSC6Pq2djAkr8qKzQswSJpWHAMz
yiYCy3QJwo86cyHiBR0q0RA9I2g3i4uZFnLbS8f2QkS9oF72Llx6YSL8E0/xpAHMAWtPrB+EeInn
EhuiwCTDsL/eV1mp0wZxijs8FzputMK3NtVRA7+lzmREstNVYGN7jWm+evc/HPj7dEZLIbIn2jNX
oSZlz1jxiazlULtJ+BbaB2e1/hinVmm9cN5QfqOSryyqhvs33Rs4ubfkcu9IRwilEdVD1SGjyBZ3
+JkFm+dD4EPFFCX7MZ6z6dk9PqfUicDSOOpDb2kmf2TCkPeL/QyMeLXNEw+zmiX7ybv77LFZoB3c
e4040pxYkb0bH3OlZ6FIQqgQ88Me8eGDLwEuhEy9po3mQVrBChPcGh6iGkOqj2xYdQuV847NxGP8
b0NC2lYhNuI2EEVgXSNjU3ydjIO4CPTp5wU3NC9WmLllkq6q+0RcltCO0i5adnPwLLrBa2BD1TlN
41wLjndxWbpZqGZQKLhJoTENLc3RZLkEAl5HJhKFc9M97M1u9osz6NFbemPdKU63Xm64P5opIvFD
8FPzTj/u68t9cDrCISzYpTSy/ZP52oW3VYz4LY8cMxZRm5pW97GS4ZBMWVOFOLO2wbju3mrnHjp/
4sOIQYqPl9hKxPu+zvImBY3O4zq/LiA5/VxcWlNSoo5IaglLQfgad4e2VebewPm6yrje+ccpZ4C+
CK+iQ+PeFvN3OCxDsb4oI0VQ21CWgEJYv82Flx44yT4rT7gcl1SEeUASJPbNpLwhqjRYUOmBf1CQ
k9nDFUsEVHj7o9Vwb2z/CavvCXS6oRs9Kd2WtGkEF2pRwdUFv4k2zyo5dPhUoBoqjUfEF5BV8fb4
6soYh5LWHDrMTq9JOkjTVgz21lntoIwkwB5PpvPSqwFIzEt+X98TZuKkbMcEV5qScL15m6bRlfjm
IR65RQR2TdYvFVo3gmqk5EHNM1G2gA2YXvkeaSezwY8UqvpHeqCk2aLIWn1kcOD8Yyyd/hOkDru/
90zv4Uf8xeh/ZzukwYAbOVmm3OhFCO3Hl5/bUxwkMEkFwkRp0GiBLdGMoAYPOjgjxq4QRFSqFUIn
gfKd7GXyyN/AtBF/4JgrEDHlYZsukDZZeZNf4FtnYYhiPClsmm25Bf8Vq7F7rlmUGpJruVIaCEkl
XwrEqtiMw1JTfnfBRFUiizcYWLWxnNnAfCz66G374RF1HOZgWdJUb7ehDs+zpUfEZBiXfAG7MMC2
Uw6LlyIUycUz7GxJzU9UoOXAdFOjqlG8ZUGAzuJT+ONC/RQIME+x4aevgLYTYmMm191QotrkIur4
h55+CBMHwX1gJYQYf0Nanx83ysQevTGxLX8BvzD9btkGNBIVR2gBsn1JFl8sB1bWHl/2xjcmSqII
oWqwimS1Abqbuw8CaMY5sSzhSgpa2i09HHo7QPYlexricuTr3vYc5smxbPpin5dFV9c7VcQIEOuL
DIu9BEigkPJ9aacy/JgDTD37Op0kGLyWiJOE0tPIeDhXL/ONueZms6odt3Yg4EypzzHMfHerafJD
bZvUf6+GtqPdOiI9wJbh5qYQ1WgEKQrXBHqQkg8zgNUpKcwd3BAFJXxmLt7QJuiI/s5tIs2YvVlP
KeERNqbl925Iw5qXJxfL32VklujpaDnU1xXwGe0mMWEwPgJTwit9KJnySqaio9bRHkkwaErOIFAu
XppAv0qTMZVaOHrwb1nMsehGNlMzFGoDkMW0ttp06Zj72rFo5FNU2Sa1Rkqnxl34cD1cNHxUuBAT
CQvbA+HzN6G9LdelGuYLktrEduoNbwcC9uw7AqCjHP9/EQ8Zjz/WCjUjnMdpey4HuhuBBKwmZbrM
KtJVJ7Prsi6oqHVAd3incTrcqDOJBE4BkpkjiaD53EbBVSLmXRg2IPb0TkU/KLPAzfJedrOB9UM5
2Wz1XGSAHHFRor3yYxYTyuScqobc3rXuFsqiTqTDb4gshQKhwQjID5pKAzCkiYiAZlk3eR8sqfEX
W74cYRHQhToZMTRA0WmHbPqzDDlCClH1IfX9qG/SV5fxRz8HVlIbz+7z+/p90KZy8tob8n67YTut
PP6LNYCMEWlS8d8eqKV2RYgmxi5RH0ANJ3BJnwkIqeDwUvnckihBBlUQLS//Kw8D1DxeJzmm9yLv
m5+Bkse2kBLpzilxWdYcZP0gCtnvr+7/hyZipkZKL3g3pXQTHaSvrbzsSd8bu7v9Lr3cGGKilNdI
FFlL3HpdYQ2UUsI+8t7IkG9s4uDJrpbcaIjYhhNlmfMj9/Ms6w23TemHhEtggajLVv1s1MhUysZP
UcppXeCKv9XuoSJhDi+17a0hSgBuwBDIVZ1zk2/8LBibzRnhscpFYrM7H17FYtIDkkuchnA/E2em
7O0JFG5cZq5xCd+MyvYckRGdAkoPcANqjXhwxWi8jTcK8QlpNywGLR1oo8wHDGE+tgRByI47Aj34
/zt6DlimYT5n7fa6WJh4Ef27fxDz0LUJR0ZvTsQTDgkfov0Kqur43kZhM73wx01poszfPCzKNE97
K0tQgo4QCKFxAUHs0cIBNxwIypFM7zWbvNnqHOC/No+21N1NBdy7j1MFNn5KDJ30nn8yUYVQtSrJ
Xg72MVYFzVTDHMByH/CQdBKaieHASzMuqEqjcX640azJ194H1GlTXdKYoLGctwqUDa/K39ZONU+Q
DE+GcMmpOG0UmVqOfNsLKO/tkFox2M7iow3k8cfsFlHbar0A8hgKsfgFhpO71Q3yYQ4jO9S9/T/K
bsT5kowbpjuEugn2/mIPjcVkTm58DwfkqlS5+meLB48aTZ7lJsjAA4qjgZE1bgbEdZ+Ib2LLg1ge
mY72glE4/oHVUCMTLdG4NWXnyMBPlNGMVdn5byw24ZCc+WUKCIp5olq85B92moJWGPh5kjaN8Mf9
45F9T83Rt6WRpKbbDe9xZxOpMb6P724EVBIxmRMZIdxOSXBScU6z77UP2Cr23kWSuMma9nRVRekV
hM3IzMVtSl7kl4QpfUEmaH3P9m3NQUe2XkLYHpH/kaagZDT0y5/vDyGvwG7SaSccB9TFDko+bTYL
054KLG+PgSqDLJMSIWW7kzK9ZHtOAvHDo2LjVXCO/zqlo2i7WMNisUtzdDhB6rrwFveDIGr9QEAp
/g54ezHj7JB7loKQNR9odNXm5ZGT1aOT0VaX/oxuUAwgZnlO2clOP2B9Q5hwgxMzfPmbXl3wP6QB
o1SYV5K2C8CvQQ8AYN2Xj721ByEhkTEMRuuWFyRcbNQlfe0SnYGzYXy58ByjOKp+6M3Q2UyQIj5r
DJ+aaECDpWhppi5uGW451McOw/HW0b48p5kcVzndBDy673ZWvScI+LdNCLCxhZIijNSSb5KZ+NiB
K2fA2uVn8Dri6E7m62c+UXFYTZ95vQxoc0/tY/xIRYQFb3yOhNNcAH+o9cKDQ41BToKws3rgbJLm
v1+H5IOj15kQKoEXsBEXoXTS5VfqzDBi7Eh8SbD6WGwLaLyQLJKwbeo2TXyL95LE7JJruY000ox3
3DnGjA1MN+nK/O8gqQnHoCYzQsoz0M6ZX7evqKrPi0/Ohiz1YF/ko+wKztlHZEOddWGReha7qH6M
fb9EQAD8+OjsTWEbEllM34qmYO0VgMZpgbCb7kmSF69zYlo2vc87m7M433AceHPdtaY06Y6zFVlG
pW0e/dJQxorLgp/0iEl+fKxoZ7SvdiZc1PXO3PqcwA3QO08xDNkTFCC4LYNE4yfy0p0ahYtitpta
3abBEzycjaBU/sdvHJg+U+fc0pS1FCVNTU3OYT1C/Kl62u+ir58BgBdBpCLfn/Fz936le24/oPMC
M8mTHKO35sr7dYjj07QxebAUlGkeK0h1G9BpIc+582MllLH0XDua6MJuSrBDrh4Ht0tg81ca9XSk
IOOgG6xbzvivJTZlXOmy7Je1S+ZLy1XgfiKXVLIUO9O1wrYn2lJVjG/AbP/MOH5k/eXCCxsKXeXE
Uqv/xwuZKPMxSFJHDrGVJyxwIDUd9ntLFxLVr8ZiBP6HoAVWtpft+zM5fVCDXIObhviUMOh0C3US
3WGV1RbpGzdh/xqCSttR0PKLcEosbC5S4vD+nuICJ5kSMoqZwu70DjbrVOS6+JjUSDd/DTEZYf7d
bsIo9FNh21LSkNkMkiLK4WaX6siMd3+HH4fL2i7TIPGRot+E3W2JcFYn2TrLlxqT3Uh7hChNFNaH
2EJGDkP0NzvslQbhpJZeNqYGApgmvrIhFhoYyy0Aj3af5QUSj2wzO8H0pBzAZhbQ3ANa2QYxX4en
TUDhZR2zHfK04grhr5ZO64ssgUy82fj4suP+lkHrd96jRQ6Ny7BHm2APB0m5FvR79fDWsgc+Ibmk
k4+nEB0XH5NHS8Pp2iCFHysSiDOy4x7EmvpEolfqczlojZnx+m3+rmcDAxpAPTF1JSzJn4kJNf5s
07RmNSqNmF95Evi905cbKGJxI156NGv/rjX1X2Te6uUhFKGv1dgge7FP69Las7dUI9Bam+0lJc/y
JH+OM5lK+hQJx9d8fTOpUxFwNX88F0+mK5P7hS/PqLEfUCiYiH6syJNlM+/wjGPOFsofyeElbh7Q
LyQWPoMvIRuFrW46sdj1oFVFCugkvJ5sIrvQGqBEbMBU0sN4B5UVskBeahgFAoooTSV5Jh8y3Ctp
E+PKhIzESgARk5ris8xJ0Hamin02PFT6tF+n6KnP9PrxVf2Jdv0Aj3DRewrtg8QvnZc38zG0mTbA
HSQjNR0zrt0bQmHVzO2J4NOw7D27yXb8p5S+nOmyxylWtZOBnVolmcMFTOz6b5CXAa8MgpyMkffU
i5aUq7On61ZKZcRIILOOmkhQfjTtVp/SoXCLGCEC17jxF5xIXm0f729X5kK/pDQ8jIaqJFwHDa2g
ZSl9+TdJ33duv33YO+Mr9ii0xGOHYUKKZHVCPhtsdTr+NkSXCAo2WNVBqMbFFup1jD1BzpwYBado
DpUtWvE819I4PA9w2F9g/WM3w7/CEEkoeLbLxODlKvAZnOFl4ZYLHLn1J4JXMzQNhnmhercZSiVT
tz6mHLvHgpU1EhtYreUAWOki0ZW6g+xmoqcATC2c4/VCeLa4Oy7Mmil+FDDWRiZOkA0tyUDBVPXR
fzZypD3iThhP1cYzljAGN0cqEqF53MQ86Vaah0jByKqrocyN9Vb9EMy6wwz+DD8RO7JywSunddVU
B3G6E+LLxmAW5uDDz+MgCF3K0T2j87T6peDCdo+raLAmokic7lquCTOdHAHJPXUblfLE45XgldQs
SJ/CIOrOQ1AchR/D3DvqAPI8qnn+RbwnNNv493k8yJtUavjqQuf2Ey3q+KF2bkiEU+YlcCEI2kfu
ncBJyktdLJmfOBOxrpgR3VJL+sreE4MdlnOSN3FO+nm82V/wZ4jI9PX1j98Z9CMZEArHlzdKpFu1
i1IjBkXViaRzEColaqpmngleRJE+PI4S/uNcXxg128znWeF4iQUGfAH6X9yzQ9GFpv97PTC6LIlZ
sYKurgvqxpTbBPRPqf4iqkaxFg7y07031SxvkDyTQBpX+baMYnNHyhS/MuI1t9QoeU2o22QrOP1y
qHylHWwqomvWrIE3lRnmNv13FRax/y+4aMySnR2yy6hk/s9ilUnxgJKcByinwNPUITutHqUJ8mHp
IGWoICOUiOOClhnEN0/a9miLeEvTBgp/NRj5QxMO38HFk763K7b9bPKxuRzIuJc1Egs3UGhotV5Y
HY2X5lKSiperWlJ5L7vX0jowlkvmUgTW5kKIxsOiqv3CO2ep15lBD5fUsn+JGjFuXX7qNlc2bRTR
pbkAl5E1+O8sWOP6bN6c0Bttmb3jrhR0ucs2wJJaI9curyJ0CaShnSsiX3O2Dy1huzcLoKCA8q2E
0FSRtmXotxqnS1EhR1o0Sfez/bAOtCfOdczaAeCMF8EGxkhaHdAkS2ncbP1HuT6hmCq0n4HILGrn
xPlY7YRZVXQpGhVJqqXHPL8z+z5jkRDtODVD8MgtE+5BjIaWrC91R/4kUH1JrQF+MxvbiIS8kCI0
aRACJ1k2XP6LFEl8ho7tzY7c6MkornhS6MqaL2yhOc5VGOHeS0PbY++2VVMTyeiXfbzLZObpbb93
JWlazTREHXVLndAYqTBhm23n6NAGzcPGl/pG2DOKO1BV/0ZQ2OFNIGl+7MgUxU0QGMF9sgB5SqHW
rdr3eudY9s9RTnLP1DhTXcQwxLyJj8B/edkEUenzaNuACay6gHUERnkWMnG+0atBaKYlRwPkXR/p
Z1fz+IQR7mAYe/dSWW9Dhp8AheHeZKBZcMR1QvnB1WzQ38l8HXkswLt6TsHzHWK12rbJlk0NUWn4
LEgmuudwFSFlLRc2AVipb3fXOsv2zo5RPMG7GPqQ0tkTtXCAl+j3Ul2Kw01OTVgxLgc4DhGei8gk
K3rEmTVjnnNw6pFLUs4NGOcMnpTcgJVZoUKjvQncqwatmM8eKBf3/fzQdn28dzWZNK8NdGJM9qaW
EUAW81WgxEWRe2faZUcWuYC2j54IyeYGWuvYyP3H3juTmXT3dyiUJ8R+GESrKMRG0LzYyNvbOI5o
os/oj02WWjEJgu6cypNj4x6KuCZt4TkC2DrYGdJ65jxfXqSNwURlI2dShrSRI1uECSuH3ioqlGvZ
m26PW+bOC1Hn35ijcTUnRMaVOqw0lbWqTuDMHvb764Xy2SUlEAXZi3zJMT5jHFwN846FWK93cuKM
ztApM1KG+6ndd8zkKbH0im3h7/3K2UlYiBN58mQPGia49qOW8+PMIXDVzGUD9lBtuxtoHIL18rjs
S4yIWM7CtzxmD2kBk1p8J1wTE3SBq5hwOnF5R0+SDv974Se4cMVmn1fcQne/tct8974gvsJN7lSG
Is3zHLrBPwebXUqmbERblmsR5MWcjZg2C6i3N7oeumJXKvISvDKTNuL0vxZjRrBJdfjdxUXZLt6r
87HNR7C0Ueyu/2pOMHy71l/fSuojubnvJvBZZGmVjBN6mfMzPy/CtX4CGHMd3+YsnHPuDSE+UMic
wXMGh9LbxjGQJnGy8VmFsqsKy9LuNAl1auOhKX273UrdqQ6Yj4JMn+xJpXcuBsBSg/qypQjlvv4v
PPbbIWAByCmixbYVkpi8WVEcxGjdqV/4tVswlJBMGMnt50JSIiJWJIEDXRGTQPn8lBDkAzKHzGp9
HoXhy04QM5mpnAY5a+5NGJeRNcDWHBlVuPqNf6UaZAj39dODPXbs62s89GqZTQd9RBX1+xxcEJX2
qUQgsqXTfkWhw3nfsIXS/sHL/8vYRILjy2EhD/wsf5ovo77eV9cS6Faaz0mhhbBrIdrOCMtlhyoM
nMPfHEK3CeRNZWFwDMehJWn+SxyjCAyRg3FnCwdBslQK/RXNYXM3EiJMb6b8xn2nQXhTOT42Q+sw
FdAaeQAhcngxNzi1dKzghDRN1y3p4AnL/WMr9vGXONLFAHMh9zjiEqw3ZTtvKzDllevtC4J/B+lM
SHc4ZUoa+RnYJgDKC2VIy7HAHrbZ+/wHGPKkuYtFad3ZNV5Uw17Ub1dCSMIwCgkjUFJNEeNKtix1
V9ji5R0aHOZ9ZujnBxq3sQNZbB9fjIKhEh39LrjiBt1ZucIbpJb9gdySsf/p8hUm+LEmhQAXvWnN
c6KQfeLNNUexYHwQPmyuv38Hw23nlsbyitYDOqUF8zZUIKJzCn4qRoSZvlM7hn/AOUFq0Z6sB2LI
OyGTYvCaeSkWDJHuci2L2ESY/sBxURh5YN3zJOHIXRgZ/yNREMtM6aK5s8AHMCEngC/YTptIgZ1F
sWtWG83yc6WlGaewz5pzeGCwsJAWgeDOBp6ibIqaMhRo2Xdy38SFHE21Kb3FNO/8MUy6emics1B3
4GddfDnD92b/HTtW/TyW/dvWo2sCK4navFD0NIntjaDM/koUshKBsQTWazmeMeEqItwVJsGFYgob
7RWo1VQOzSJuv5r48+kgt2aSj6/8PGTQR70vGt6LFw5YAEJ/c92M/7lTPkL68wyQyxLe1HL5KfJ4
rxqCnxfjc8ojV8z7ehIwrt/UKHAegDXcm+ZvwohuQOqvGOi3wMQ9DuqWBPjO9u1ORMHXS/EelU1U
AyG1KzXdU16uTQiRWhXLsThPW7tzde0LBeB/5e+hviRjWG3VnF0rgIx91nhqBDmLEoasNAsL/0tJ
j5g0EsacateF9XgvrZkD96Fs04JyVZA3csFGw7xVvk6BZYxdPyAEP6dT62ftpBdc+i/eh+kelN4K
uiYmSI5odpzrcoBbsrgfgzVXIAYG8uoBT1QfOfOIx/0EugaKe2Gjrc1Y8/0krqgEBIszpXNtC8DT
okjoA0F/+2p40/dgS1G2heG1OofYxGnaZ2PZZa7BVDF8PBnUtn21LdXKpi4XekmrSY5vj8ouOsHP
OQOSUsGKFdWOum1CgmvsAwCX/hnmJfKab/fshPuYpwbyCliMHZtqrOxnS8CAXSgCs4eJICbzAjFc
ot5SPROBHFnm7xDi9nTrsVKvMkBhsUtSyDQtrISEun/CDpfQ7ay7dhoWNqOtKL7kA3cyppJfTd1v
aq7PgtfcOgEejX/bib2vC/DvWHeQ2OCIrAi9gnLq8QOwjzXBSP2eGRIvfzWaehNjZK6dAisAYzYF
97cZ2S891nW3B3po9yende9a6Sp+NGB+0MN5Wc6xCJGJYQgZbgw//NJPN9fOC/iwyIMY9qP+maf5
0XZgFY2E+P/W0NfvpDdALZEMMWqUWqIRBWYG7SHFmUPipjNk0cys1VUHiWNutURVIocDMDbcNmzT
h5T1ss3tRT2wmRgwzAiYuYjcMyG5Y5kV1hn+frkEOwaszdHPaZGVKue1jHtB6Fp+KAVtSE55O2QL
+YtoFZ6NRoc41r06G4ZhS5mJ/rjxzx8dEr/3riqPvxe0BMmX06UBsIhOXpFwcvqNjnqjrIjKVqwx
Gs6JpYWYZcHUOFObsAoCK2UAYCSNueEWNnPAupNupzQDJTv9ESjV31CaLggQVoc4VbacCOjU3mBA
EszfjLFq+ZtilKuG/uFi1x59dU5nZi7cPCEEoYBqH4rORKvUVdommXL+qaJFujv4saocLR2Ciey+
eb97wYIpH9pNAO8IwEyQbsdJV1bueW/oh48S3nYIv+0kYYB8HABs4vGd1tPBieM1Um9uPuojx8/3
KvwplwoGxlMgw5TQtvq0G3+kPtGXMpqVLV/0iEmcoUVVQCUc4pz8RlAv8NRTwOHjyLtH+MOuOxMX
U14wtM5wgJuTSUJdnQZ2l1/DXM9zZet1d8Tlc3y9em/+oWSBxy3SOT0s70MbWyd+45ciDix+J1XQ
U5Pf8RK+ICR3kMl33B8YWtVexpkWHvjnPBQpB9x6oWycI8djM3tLQwTtPW0EA4rzGj+JFffFsxVU
Con+/qQdbMIL/s2FKzR69/ayx7GPdl/UuxYALZV+gddeYDeu18wzI7DuW1fqGUtmM+PO66XsKe8N
xPWM4rFmJ2ZtJHbJR9EOHnNz1xLHglZKb0UBROIDXw6Hxv9Z5aoKTA9ObRydaQ5dvCY9PJQBzOrF
21ZxYahS/VzOv0s8W/P8E7T3pdBGL85Rb9pRYzJBix77c0vpUsp7su9JRC3jvBaemk4/ageXnGFi
euamO8HXbEdKCVXL+XPeF/5pBQ4UtmYvtIIDZseOIvleayiJXQHTiX/4ttD03QgPijY1LnlyBE6j
waAo6ZM82v9ZxwNgt+BHi8Y6UPYiVxDI/NwUKsAVaNom5xmk1gVn8awgrXVu0F0gHB/JRs04FFh/
AjcBgdNG0T4Xb3ZhxBc7bF2PppkpPLn5UYK4anqht0OYU5iR03Xf5s3P4qEMwgheEwCa/9Rtu7gr
MYCwKyKXE86II6J2SWOCbx70oBazEQ2gaDnFLHVCWckc8TNmlqGaLcSMtXR9M4PBRjASsYXNy/l8
iRrQ5L9RxyU4lSOvslSnhezOh8YQlWQ7zDFoaFeHK12ouIXs1ivfkO/ypX0hf++Ex8NbW0w1zAC7
cKtAy7j3tmD0rMXf8QB005+POjwXhf+TFJ2D1QKaUSvTSywHu6sXa08qtXGEu0SdyzozDhNu7zIV
9ToJRgsgqA03kIDmHKgNO7DMrF1ni+JpEyIwO78HFAD+UxSfF+Agpg5XSr/UXXMCdyzaRgSr/tZU
V9zLxbEU3BMPBK2WeXt9ijqyvi4r9b2IwxY5Y1hFsRE25Ol0NwAylxHlxFICtmyzQ35lN+IdEB1c
3WsxVyQ+h+6zQg6pxaUYnVYZRmczHv7fnHKWL1uOXEsmcOJLANo0BkhyYsu3BSHRTTBSX7pTGRQN
4Rw+iUASD/N3K7ZVIpNEtiOna3WL4Syxyztlqqb31jev49NT5197MaRTsYuZ+GmJi9bG5rRKh1Se
SLodk+00rUkoJPaMAIW35fkcGJMyR/CEQj48YHlhUiTPrqg+ye1PLZZkYX+6yzNclUHeSJt4/JZX
Cm2e0xeFOH3Z4lpC3tBRz5K8+9AlvA/MME/7ZdRfj+KmHsxuY5BbicogIwnR3bDo5qHSpeBA1aqF
JLzT52pehzsZBQ1ACF3IaP2ELo3HtYlXHb5Glb7YAls1txTQIVaGLlXGxepf6e8LpIQgd2JN1/7w
L9JmW33h2Iihx2hM8yskeRmRuJK8XeBqVb3d0vSj+074qJD6mV2+ImKejI+W7owv7FQ0Ckwf0si0
uAqTiSbOz6TUkv6wWe4JgXD7mE/kdOpiAz1+UntEVT1hwao/vF8KTvzhzyUo+mChkUIt7jZkaMTM
EmTj36bownWGNiM0XByD1FrCIvGBKQSmH0ycGaSebOHvJPU1p/FaAuUvLjVbUPeJtl1k5rBo3JJZ
hahrYsiuF+Kpvo8C2l9dyLzYB6yYj+ZP0ZRJ6i6C0MxRHKSd2a+Mh7bO/44cfox+tXQNOkzLs9/9
b2qspc6sIfm3MmNO/HUN+xXqd2jgvbqM5lgx1FlLzy8GA+X0FSr/QLmrb7cgpfL8E6E590pCg8HD
ZD5uqZm+jwOUOP/H2YehAwLznX12vesT8OnpXXgT4Cyabq+if03CnOLCoE2TERa/GHSOLaxWUBze
qskXi2wSDYJRlgv31TtsZ27mnQuPecbGXpRddMSjMFiCHpSbhLixrJkIfc/JmTAehb4/ABp356e/
ITRrDXXChoDoMlv1X6TL4nQPLGY8IEg9x7PLuRjVJoAz4E1VuT+/KE1SYfgfXn/osuUxlXMN5Joq
Bd6/WiVLCgNBbVSaHkOncZO8Hp1g4iTW4kWNDBxwgc/W8W9vloLbrmOLkVw1mMEPYR00wilXDtZ9
+xHlQi1lc3rqo7aApNUscE+iTX7C0JLqmSIkySDBawd7z3zyubaMlPaLTeCGmfabrkoLgW1wsDo1
ab0cyggFrsSgKPe2DRNAqcRoaFtAKK2SC5N9DehaWI4p1N4CcMMu9GVdo2ocWdvXMYc5LAR9KLp/
6LW4VeMrgk+9aJeJjixiuMQsY007jEaH8h1VPFwPpC8HGDDGWjaJd0jRkH7fytLur1b+Nz/mTvXf
97yv92Ed+cirlya4SUm8VKgw7bYspvl8ZMBr0cHwSpRFPJ7NF8WKccLo/GcvrHCpWj9Jym9vU19E
8hcBZkjetoCOr/acNLshlcNLlUALvOxeEKUIcaPuPJRLdpxuU4jhSI7RarKNXenEgSZa3ZrUMHqC
JDcdnW0bnPIHe3L9tyT4PbucQ2pB847YWW8kDusfEhaJxmvLouVDc8qnm5vma3CR2k8s4a/Y8+6P
ogaklMnh+cMTwmRXRzVUb3ZfyedvgBJ587v07NEwXBXbLqAVOz5x0ccpbtjCaCbdyyKGZZe4vC0+
mZvtJM8ATyrxcq21XVxcFVuzU2Fl1nX28xbwbEocGzKrlehYgbYOD6tv5ZDggECVU2g4TnG8wsQD
2bJve/tCyJP32kiHDSxK0HA8FRgSFRsVKaylADiMtOgUeFdR7UKJq9WY5e6w8+1i5dC0vU0l2m1x
w/lrDQdgKzC1AOpxU1PyKvIsyyFR2veYJPik690LfZr+y0NuY9F1QN4bdh/99vQFZ2Vqn3hwWvAI
7jhaQypKNiZFoZIwtE/JE8RQQ1O90EQEB1bwbLSJu+6tnWU5LF6Z2TIo0/jonQl4/SP8aCL3C5ws
Dzg53nsYGgFVX/yzUV6y4AFD7DeNtv267MsilvraScQFwzMLG7UXlaC6baNVEIjxn9N1DXmmK9+V
d6C4z4PDtrYfspMbnEP26DNo0nEjxzLfH+agHznsSnQrIXUk90yDguusT2/C7b8gJe0474b51cUw
oLmw6RfHsdutvekTgwyQ92pqMcOTRxvbIHQF3myQDD/KthokNL3+l7kLXZ9YtXdCRjIiY6Uzupy6
6IH3U7Or+/rY8rm6rHXuU3v/4i4kg52bwaebJWYjFZeMq8W3P1rCFLHIrTMN3bV5qXYfpYv9lGep
MSmArcKp/aKeSScV8QudEVAXwKJUUuisdYVfrREEUyOKy5hoMIDYZ8Ks23klit6JibvSMM0zE3Qp
2uxI0A/f8y8vSFDmCCZTxlPXLm5/GChpp2iwiuFDaIdTaESA5WhihEJ76n7tzALjKTm/e9HDhhWG
sNtz4AT9iIWllNtECrRAiT/eJMAosJzArNXDrOglW3GasiSm6pTe80tSYI1/APibkkZHKst039sJ
ZM8nUeqorW3KQdQQGetv8otTq7sKCgksLeMX8bUV36ZXE7VJROcnGbDhvkYfjRqV2L0lNvNQVQec
UgFXPNtp0cA7gEsF6H49eEDeSQR35jVAukZww9lL3vkYC8tuUKRPIz8UI3z1dD35fQ2l0Rx8pS8M
d7CswwdpUAZHD+prjqn2XCcPr3OZivv7T4hagqj208svWVsM/mWBr3hEMqpqBKBs59pdSZDHGPU9
XaIyqPPKpZu9iPOJZGTBoX6oGQjRojw3GJZLNK+6YUiUZu8IAqk7BkREcPV8wKT/8r5AEhgYZcd9
Lu9AI8KBgGOTjtv8F6MP4BytRInY9MlWjt8pz60WiXXf/DMt+15UE1fFvKjHPVRB6kpWBijVO4+J
i5I1izEXtVMMyVaoi3KMFOAo+OnQvADxU80vt18dTZTJ1FVN52DutOmCNJuH8xX4V8v9gfkZ/CxW
4R0sMQGkCvxccYRHLteQrvfI1PeAqtCr7nOjmJXFZC17/3PcoCY9G0ffg3xn2nUVFiGR7jp1EAah
m8oS35P22Bxt7Y+qeShZVvA/s5X40y3zYortbSNUY3SehmC8qUH1Fvmu4RVOUqe7k+9cBnFr9vcC
nq5EXlK5+0nHG7gdzhVWBZTMNQRpoZOz6YaNyguAHpQUpDIHsGDDCRmRJxqx5NQA7l+OsH6e926j
v0U0Cx8vqt/RdC2HY+NWakdjxpTMs3RUHCK4i/s65fhdEJRqDFycAFKp5VtXaLzlFinsCZiliR+f
3lXPECb5iJ6yr44Z7gaAC1eygYlUuyjjfpmFkrCK7T8o+gA3m9llxtNR4UaKjmPJOKLd3FoKnUZ9
fFXbVkhxElqyNCJlNk0Benk4ltQv2P2nbFynrPJ7DtHELyCIyrdDRyVfWNR/VSTHZf+eluuzz9hv
ar3cYDZouoZ5G4HEsx+U2+vrT2Ud9KrxgwSYZrcWnBBzgv15KdXd3bILrO2Is5SIMZaLswSc7bzf
6DgasFLFIr8DP274qxNHTc/2ixQqz6ySBBDZgcnmT/PKrihm4cEB++idbC6o0EKvjPdkgSA4UGn4
4fL6jvjqRmRgYRX/Xs2Q3GpvVqCz083l89bmuRXvNmZACSo6dVHWAX44UwZK/3xAtxQsXKc+Xo/f
e8YGKbTlBdlmwa8FewtSBaImhw9iuttomwi27arW3J8ehxWNmqQyF8y74IV3yYRi3kIvt/eOSmGN
Ygn8M3zDB1pNvODZLSF9VNA1Pn3h4gUKkBYhAQOPza0rjl0oDaci4UPVyOltHUyM+jzUKtXJvQ7G
kXY2LUWSRGCFjMFV70AK5IT253IN0SiIu0ldvrkNHa07+vLaoY8OTpf3/keAttbsUXylE3ZhA0vA
LW5BhCiGYD2g2+6QfG8DDsk3fb4NLhxj1IqTyQeZfnWkDjD5n2bTjQ3ePfTRSPLyT7fzU6gJPlsT
lRMWSUOFSL2gum0xm8tNVDsTFqHqWFruc7Bv8roeDrKaM7IkTlSXLg7KFYSH0S8a+7xsq3hV+pjy
NMaMKHLc7ICMiyLzzwH8joa1+y0c8fnC7oiwZXGGJR70jL0O/uv+ndlKu9GwOnOiJH081Ch/vUBM
3Wp3jwF79mXbheZCQKSwp+pEAQWSiDzn53gV94QyAuIBSm1bW9Lt3OJBOtaKjGBeiJSvxbIh1Woe
4kDqR2yIM+8PxYpXApzkLpvdBymQ2GB9YYYbiavBoSpSboEZuEeRb1y4wdfB7IM35uPB4wABIo6w
41FL79WQIHKz32qd1+JL1dhY58aHnUad1uxNrZW0nQcPgkMDG3SbppvbHDDlcHHN6maoUUmlt3/c
y4eYE7Rk2VrHAA3NbamVIh75yAatQD5e7eX9vfk7SAeyFr4Ff+QGox3JsJ2vk6G5VRtU+XLuArbi
jwpPg6FyZkMfv6dZQSESRL2i/ujTkluYB31YCFEtv83b160Ht4lQHb9vfBWh6Qrz46ZtiVFRYYb8
cFkf9Xk2jONholCY+R6OgYwPwDZDnKchwZnz+RuWPO/YySP0UwaccHLI4BHkqkobB/T7jRlM2Pwt
aGqYl3pZNggDtLu8EOsG8KgB6fm5dhwNU91Yji5rx7aPnk7MpSrK1nCvnT2xGq1OVxCIyQ35UCHb
qXRrsVLCX633KmeF01EACjjmaZQFpUpNPIpeWv4L+XiZP55qoxR/i9LD9qUg+EXWWaaomCMbHyxV
2uoCZUQ9hAuQlQaza9fH2vDMM0cqIfJQWlheuxIg+SueAhbX0jy/fHjxw51Aqt/l223uNMdBoFYM
9xadr41GNEz4r97GzOSZfJMHt3ocaaistgm53xSiwrwd0Vtcr1+UZfHQipNiRuKNUmYG+4AcOkAh
x6OrnQ4Jmau5hu1R5Bu5sSxuSvzT6pxBGflo1qZ8VOIxWmew6ejB/fwrlUIEfwxXv0AOW9mYtnoP
yzgC2vKWltEOQqymtVSz/K9kv5Q5Po2j67Y2Fa+yT/wWgQTGzjEoH2Guqy3t0T6JXlUXStyGYl15
Wl7HUj01Mvkv2GGQM0GRpO50HBE/kyWi0yy+yAbypRUUrXOVe9/90PT9UTWDjHcRxBIWHMrRLJK+
CZrOYuGwZAv5mgRmG5xUxf25cWWNiRTiF9TphxqYNyR3OHYX1nrw7LlVJ51njMKDZK9D7mT8spj/
TytX9HMczgFjrqw8b4XHazvhNbrVGld33Z3oqPvb5Y2PeB7muFgvDL/y5lqSUBzI7XZdFiulBoPO
Z0Nnq5ft6MToNPQ/RE5of6IzrPv96/LNhSf6TYeNnuo1LEf2delZeGLiiUgLYP1S1wAN0guNvjzW
EdNl3O13/JI+PnPmiwV7yOayISwu/jutak8QkM5tGhq0sZAV8+jusoubP4N8SutWJKQTA/oa82Ly
k1I/r/6zYw3kxZeQyoCTpVBpGxtjJteYzjyXbvDnmQ0Yl/sqYydAJnoLIJvZHuV10B+8TF6e1xEh
Q1YQiBjLjJRpFPSp/u9KzN3fCnf0hM+1+ZtiPCtOGCBdqsTAMyGDJGtLJjCIBjOk+9fKDrZjqmGd
VNEkr4fHfEmSgjse24nmaUkB/CNHHOnrPUKl5SLhwfGdoH+OdIXpv4g5pucvzc7EceM7jH+7qL6g
fof53xywwpH7SSl5qbTxZCSubxWecLmySbwNGHfZW4uYUx5FWuyMnD63OdwT4dc4drnc3lm/bEUp
zefuXPgdwh+Va1mzbsGPF79CuNgahBf/UNmDCko4L44GBCIbFz0sbKWUsmRXu0Mckube3qqKyHo6
KwHWtjoL24KhWs4GM2SougJAgLKcFqZRqUnQ4Eqf6wnb9NZbqJUV32WNz06fzlv/YVOOgit0X2RG
vORLArQFRS6ZsFeiyUQa3L8uLemEdEis9gKd+g2t5pnZkg7VeNMsbJdhlTVoJbjROHp073A3K3om
8JBulSbd8VPmx0KRnWUDoeZcm94io7ulDN6uPa1cbkgJ5wnWS7AlLgomABSmQIhC7zc4/b9gsRQf
rR6VQXuookUIsVkCADF87oElXkF809wOw8y3Zsqcbmp4mUVh1I4jWy73rqc+tCfJMBJodiqFXcH3
RS0nx/hL2qgKEGi/fsuT+hfy4q9Oq9e3KZLpukfo5eNjGI+gvTLQHpYBU8Io00NN2g1VNYbhl1YK
7+t1ilhpQuXvR8ukp/Ie4ptsh4a58HebYQ4FG5+aJ6Er4cmdbCiaYUOXQOeuLPfjBT8B7O8REKNt
s+1do3pq/qM+5pIBvriRxZEA2wMywDKA/+5JVtyae3htFYeckGh2lYJTUvnaJ/lHMmxe2H+nONYt
eCrvoLa/7BumgHeVs7Rf86ISea12O/xxjeb4vKALT8eFCdZQGtiUbxw3OXO3GMvgJHfeswPUefJY
t11iF1H3xhasi4I/WXUorkVGEsyu/l+5sIoXXC5QVOSf3VNBcpyQtKWJRVYXgVIR0afnHwSvWVV9
F6qUQvCAX21aArR0wJCAs/ZaA013XKpxMUIM5zwhvxf4ETVz2wRbRf84LBFFJRqrxBwOaeiNxX6n
6zxSXRTV+eL6K1XUfz1xAxFyWE8YkRd9viKGaarB6vW92qDSm4lkCmsJKT07D2PCHXBHew48ODh9
Ov7Nh75VzQg8bk/2iFuzD3Od2p5aQIJNjkFBQLEo7HvGvUn3Rm78GC6YEkUzD73tkunld9bdQkUF
w13ipAePyUVovD+gQysweJPztC7Dr/jlysMHAqw0uVFvRySCfeuujhk+VbX7K2T5UgjFFns9EOMe
IwcoawKd156gLEgT+ikOENa9aUkRD6AJ4gn0lHMTpCRQqAsdiUxGGdfQdQarLqWmusl+cKEAhCYn
l1DA3OWF92b4om6ZIHO2bXKlYsCRaPKEepORN3t849ssrkDLD/iyjC8rbroSeNozzlwkhJsf/m5G
FmyPcFOv7wKnHz9D10lOR4aFkDurCTH0KeOwC88U59YlF/NxNj3d85rQkW/O8AWdj1IdXJQluXWS
iPy86SVsfzdQwzC+zjMLRS1VbimnFaQfRwEIt05O8icWIT6EFcGs2rsOHFZe0hs4skIyjwYdvv3G
s2vgYbfipdQ1LgMQOlBVZBAF3osZTPkVIBy+b022fniKBWxNUWdBjts5k/c478gynyoFefZXKaBR
1ejHyY4I+46mOsGz1x4ltVYwo6PFtFxNN3+6qx2uKjr+/RqmUPs0S4hkBgIXvS3IcqrYu7W3F+4K
AZiKOH52hAjHtvK0rlzYtsPBEL6ILwyWm0yJcQV/ZujsWqaz5WZ0S2K2l/u9GC7dZuoe+9t1h7Xf
R73oGFhWRkpLZPwJVPY0LwQ4rrAvziHRL1pWtPxyfz8Q9pzghdjH0xQt7oe8dQ/xFc2HrV+WiKZy
H13p+ZH0V1JrfSGHFTasS4JX7+3Lqi4dl2LzA7G7QeWW2rqCqBWtWRFGY+73cVs1XvS9BaGnpJUf
zlB+Q8KSGDV4klHhMFDawTlK/5YkdlW5Gcmh6M3y/tY4gPCGmWTCzD1X63kVaGalZFAWug4NLeeG
GbjMR75jiB/6wEaJJc7BoHhSQrM3Y8N/34Tyt1IeKTRm78Kn9bcvOaye+1aYQ/oBjGgWGJip5co8
g28JaXLPUbu3Ys2hCK0Y1tS4e84wzk33DRIQXENk7wb80mJcoqqh+zBJYdkxRzAh/mcCFEZUYHc9
3MhNeXovMElirgv4dhZeFwTfT3Pc5/F57Y4SHw+xu7/iTiCimy8d3h9JjPDUyAqXzeoG3a/mSvBM
m1Qopxq3vfeSfypCbRpKQI09vd1Y9oyVeaB3xg8Dc/755cCZjNvKcPg4HRJj+Nim+9Ct+G25FQ9t
rTx3mDN8IF+XFP07nOEcvY5Kp3Yygfuth/uSEzdC4OrhhmseGpV3c4wRSg6CqzalDeZ8lV8A9usF
GXPU20oeDBs3UOLuPXE+k9dE2n4nQv2fLP0cOL9N57/r69Hyj2QlyASxLAKjbiobqNmDdY5e2VFX
3gz+nWhT7NPuDQ0ZX9VUaoctCf/zrGP5odk0HJvG9Yoe7jW92hvw/ihI5E2INnN0h8ikolc+UTVI
iWQjOUu1wDknJ+UHkqFWCyOojzmJY6UY4MKQnZuAxf1cREBbEmIAUkON+z59UM6Dof3nYYiHIjD5
wKYT3oxUUy/f1eCVowKz/9A6OVtCqR1+kECUTJ3ES3CEEwU7CYg1g3gnKZUN0JGBSf+9whFomeDV
KTgUurOt0qwgUA30hTo5b0AIFXFAvGfZQS0z5WvB090ykR8vdecTPYTJmilG7nPtCSBDQ8RQ2g4b
PYfL1xGobu5nj6yvGBamA7m8th7Jh1MeCAEzS+YCyHPFw1SVQZqsNrvgG59bZ4WHsjujCfFYBkxA
PrlmnnukmEht7B3aZBQ4UxO1rvGtA9V8rWpQpniEn9721swSoHfomPQjaXqtkbB4mI4wjCspe9kr
Bxn42NdmuAkGp2Ms/sjSoPNww9nes/X7vEwO7dmFchl4hD6yeKwgAP7HRDY+hKbLU0gcA7ulw0et
S+KtncmrVa+UyykVES0rzEZJtGZBR9ZHCxgVlofaQcSkGt0UNI9k/yzAFGe/YRWNpb0gtl/gtdc3
PE7N3i6NYOoSPwf3B434saF1S2CFy294qQ1LzyEzck44IearXKrlu4Tvb9KnG3GH54DEjNZBZyj/
V6Kpa2wOHzrkIdwpHsgk60K4a6lR01rJUUbrSBpAipjVoGjMEm5D4PweWC+g41I0HplgSQIAfakr
lS9e5XcLGrevXIaNbPj/aaxTOz+Yxd1j6vxJ85tnar5LBDU9BkSE39yUPyxawiyjUCao754y9ObU
lzu+XTEC9uQHDgPj5c22r0+49hQExbvsIO87KYQBxrBTmaJmEZtRghLWqL0opmxWrlb6N2twpeKH
aQ+UZnKWKoDBoF2ki13ZFkdZlA79uX9UJ0ybjSpKlt1plwpfqPtWijQ02fS392awaLhwPcyNzqdl
p4NhI7EbrCMAj5wBZD1gZL3PsscgtRiguUYnvsf5h1nHVOMywN9XGkFET2TwRJ3/m40XsXf2HTRQ
vULdJt7/k1D/bGnL62f5kuJtmtcqIWn1uBNHKp+kKFo5MTz/p5q0QB2QL5/GxKvibj5eEselDgZS
Tdif8Zcm2hATrz41uII0rnJkJmJ4isrB+yZAOCGtrEPEy/rMS2d3GYa0ppCIk9Km+V1MYGQt9eVe
H82hDlR3bBD36STA/gCpNFX5D05bIseKYOxUVXnlbHjNVye5/BFOw/NQCO3WtBtDMsSrNxUR3J3g
pHXrI51Beh6Km35CUyqGJIDyZhIDMycXBPLrh1w8QOBVg3keqK9bsKJEsRTI1AyQkdFoHmhxOuCQ
9GDYDhT9RVLuiZ8/zsCwS19hXAxoWO+v23EszBa/5OFUpDZjKsLmHh18rJnVYBYBSuWgBdDRl/iu
NDgbjNrMI8XyMvKK8/YriiSIVSFQHkiYTqqC1t3SWGOoPBnfFcluVHni9CgPEhJNhg2gtXnb82+d
I8rbb2BaIj44/bINJNUJIIg4grbQY/ziYJFveekmat0uRk3IbeyWwS+4+nx4bJLDfXj/XzuzVmdS
dJrM5FRsrow8K3gPOoYmp/AGxxOwcZbr29NawVj1HH4tgCYE8PmZ2V8O0tK5QSkjCPSPyfTK3tAy
QbLhU9VPE2dhece5oCzkDD2B43QrNXqtogscLWyCzDDEUODM1liyYcJUxAVWn2t28FWstSrWjRaB
DqrEW7WNrbLf35Np80qGgni3icpxvLD8ktlf+Tyrx4OIFNehzYXBjfNbCS/tnJzAo1ZD1aIcxc5r
bDOoGnEakPGWAppSpUfnnJkBgg4j3hVzhN4weRQwaKW48M0oJAWlykTKm+3lFa3x2HnQET1UpRYH
l07iOv3Q6F9JFaLfOFnkgJOgW6vJ9LR97v0FwcRWU51nccN5ToxL+lnxObTMgqALWBZBIWhC/fNQ
+N5LWjjCwsmirGZ1nG5lS+x8XZ/y+fPhTtpGg+9YWucf0taX30ZhSrwLN4abAFRE4Ju80UXts4fp
tRsUXHzTC5/07N5PcXpIqCqRQ91rFr6/8FgEP65Jb5asJ+TqPemOAbDx5IZYmRUZMqAlkis+En5W
STpyVlIaNAzYqzoVo5HSCjBfzgoSJ2KVuAPptHxjgukJMF3OOMEHsRD3atvfdKoVvrrC/PSpzPmp
sQubIk/d2+pZc7/pDHZSUev9U09XWUS2PY2r+AtQQ7UxORiLvuRebgTTJjwShNIJlfymfQfcQSpX
vpHjui9vqkiCG+anwvJ7aa+ZTouJnH+kYAxIdIvEh5qc8WwixWy+A55sBST0xuZ3oM9xXVpNa7kD
nuEBzTbFTJNOvnLXtQnduCVh/qR/18vJ2s0Y9efPsf0AVbH3mmudUmW9fJI7/M7eJzpLk+RqTE42
JyfbJVqtwM8CLmRiHz5F7wkIU7YX4OEfhO+mFbUjIHM3pR0rT6Fe8L26DSZkW5p8qKXq+3vkGHpZ
wY0UvAGeX0dzotAlTsm9/wyqqDtJbrEtGyURRB9Qs5ADM4onMGkNnKpsuf5INvzaihYbcxv7t9K7
TzCiIjo0tq+sIaI+JEEcpE7jowwD30/slPNxUkkQ4PZVdT30vDN0qH6HLlcjkVNvDMauG8eAfLed
GWD76j09v7rSXHg6u/VjKNO85wR9zOxQMQ9guZ/jE6LhCsb5vEQ4N59+FP2TP2gALO2zxBlPkftR
/Im9W25wRttHVTV8MenLUcGu3QgXJRu4Cgy9axAzk+7mnVW7YI8S/+VjbUUU3jjhXP8vGwEHXKUa
wE8LLzzdxz3XCMWR+ow4/U24sUBOXgkIwNDcYlITs96AR/OJVnfHsoQvdZC8DSxPs4WPH3WV7lnA
wzo4d/s9jnPsxeyZKEBOU3eWzqP8KwJq4oSpPwCuiz0CfFyMywEEUkRg2y+4VnseBNoH89WyV90W
+RyCyUS8LNbU/HMl9bs/iQZ0z7Ln9FAraSur5+2MstriB3dUQ+biwp0DTzZ1Om7Zt8SM87kM7iS+
gSB3dySgazxBEp++1PVQsRbVg1AaF73hNRNbO2HAFcYlPt1k/R0ZDi/H5YZC92FUSo5SOT99F+M2
UPsh546KhFaGht7d3gcQliIhQ0U1paiT8IZP/AhR9HWfwYKNR4fRli8hV1xs7dep7MiJNsS3S9Iw
nElKWbVXkKvLItIMmwcdkMYHn7azmBxNQA2zsuNuVc9RgB/pTNC9jjHmk8WXt0ZfjAMbvwZHHTFx
CBvg/1c6UzBpUFpQ2dAgwYFduJjBaoUhV/r4TotXpvQ5p1WRPT8amq+5JnnNXvquAbgb7SAicg8h
NBPbHxDLfxrAHoc4oJ/Aq2vucWM9aSf4jWANVGCKineKevXughcACpjcD4iTPr3Watdzql/H30ee
oryqABNNdSPkSLF2O6A5ugd18ydxQABrjgvwhPy5082whd65u+3zUf1jV0uCOBRqD5csM5ip+Yz0
BCNIM6KxOd88KeywG7L3C8WNLTDbvMXonp5hH6KJudmhyVzyr8e2hZvrCHS7sp4LqCCx+Mg4+qa/
9g6RPNw0/9jbwgWswX+ajV0AmMxiKtrzQIajKQBwrHRSm2720glvNoUJBlqY9OrJQA6RwW5Ru72G
Ao3L7xZTj2w9nVPHNRitNLWBvwdvbJEoGAGhkl+AlRAkWP+O+4Pej9xxxYtnIf44j97A5c2CpX2s
aC97b9+oPlWm8/NEsVQJik5I3TGEOBcrdX2k765MMk4Jt0ZXXQlYluAlVF4PXacv76i24qlPzcil
9cAO9JwfA4tLcKjYdCDH0dobDjZ2nSoOgq4YlEF6zOmbeYAiBw4wHOaT38NGcP3Q9jVRKEhm26Xs
bt+kxgMpgs2VYU2O+3p4njTF26DHr/DREfEYCF143pr4Cg0X8znzYCLCsoOKVToCCCSzzf4tstpz
8XvWck8aazvcH/WdwtiL4B1LwuMDTcw5vsP2bqWer3Ql/GFkh0QdrWEAu7pdCpjnhj9GD2C/F/Qm
nxj9wnaiHMPB5jgYu0n/rFoT9cyP6Ruwp77EkfVUVsFxxMi61eiW+zwbag1ZU75V5l81sH89Qgbc
pojPU6VLHHEDKj0wyUSWL775S29/VqbipLWiMVpOx3Xo7OYgoQG6+5LdBwPr02BFJhnplaD+1aj1
VDgUVuFuZVYwGE89yqdUgVSXddTrj9e1Hihz6qmiq80bNgJ09y4/W5vVQH5rCM0kjzw9obGYHqQL
akjoTR1f3YbDhOkdT28gfI/pqQyMiQmUlJnZh7eg+wpN1L7PmAIi2TBZDG/eSq02ZPjeGBY40fnB
tF8pDI/hKRAJKLJX9VTLyvUyLKyKBmY5UZluEWwVBYiMDBGM+F8f//BsgnZXhtFvvWW0H0VX4Geb
6SVVSOGlaZ341HqHmCmWRBVwaBTWN3fjwuyn2t1BET2Hr3/OTSMloLL6Gw6rA91UeWhyUAkE1lW9
cChFpBipSTEmux8LTiW4L+LsDr0lxt2V6MrEsT4y9kxNBLAwxhBolN1UBRUREdsNaJkzb8L5hSl4
B5azBNV5sM6rhR7KaBKZQfinpknB04LCzG/7Pqcxll6SGPWki7qLJp5DjluHp8exHgOUxW4CM08n
MtzLpKB7jV6B5swHWUbS5MlM3iNS/+L30lX6piUhiNEDwtbw40rhdNLqRJ/XPPYSmoJZEItlJSyc
JYgr1cQKLfq4wbkKWYMRFnxxJofD1dMepjmoD0vdTfsTeUDAj0dFK/t+XsUwXXbVZd2JxTC8mjl/
QeqJh/L5adbDOVEv4VLVTIcLqjwsgwEG4VaIFs0KtdxJpBzcL3/plMcBVYDbqwxV3isgtR7voDYI
CXIge+rEt1rvtR+V45yUD1OYJmvaEESk7OQcJnHDquV9qbQ2GRoyi2ViHwOilCiT090c0er9CyHw
xIP1Bv4bi64/+uuQgv3MmwcRuyM29HDojqFP4uY30VmIrqDWWa86TQXMuLEADFTG+wPJS4o1WHbV
Al06kEayLaGCEHJNyK8H+PbP77o+jeVOyu+AB8gxsfjqLjCYFIvcVvYj7Bn9Q5UlFFk2d113WuEo
Lp8e/AIMwbGonohdfwB/i3tWfYGUJ0ZhVO+rVST/3t4Ji7/BVgQ6cJf81lLUj1mQCZhDM6xUNDyP
7h9ch0JmCtp+LvsEZAMlRUNtDjEjn0s/hYtAHbkVBVffF9qtU5EeeOIwjNcuQyMnLju9mXh4xSF1
3xIBsy/QZrmWJfkDaug2pVizMdK2hh2dIGJ4qf1K9wpXx1x+sWuj8UhrgJRxdAvfI8eNciUnD0PR
T1+AmUEpPv/eUGVRPZDDVkiSUa2GwnRFgcX9zlGoaw8oywEwARwoZkHOGjLIb+gbAzgyPXLK1pRD
rIzb3Lxhu8MKpycugYLZzLh+fjRfMVejGxDpD/nEThB5Z1ajECUwkm17AA9hbTewVa2fchgV+haa
ZVOHHNq3f6GsQCJE4BRfkvh/wmbL1wwThKVEW2SGf1doO4NzTQR5Og9D3s5CMupvLCLrZfcKutIl
Zgr5LIWtTpoofW3J46yCxkWSDL9kZnZZkdGSnlQOKBktb513S1gUgaGUlmgVPZK9IAbxzzHG9R4g
PfS7MCHCSmei0AL3bToGcjiX+R8g3n1U8WPolp4toJYgWRV94ALfxDTYadlCxezctFGHNupsjJ7d
LbiVwI3Ws2UvGwopdEfySQFzFh516y621Ga/K3bPz92bvlJwxacxMUEVW8EYnTRYuB4sqVdM/vXI
g+Z3UMurZhnh3cCi4/N8buo9hvQGhfrZYDv1gADOsivI8xAwaAWb7+3qPOPtPOxUeBH9gWWxNfTi
iP5ySEKi2iHOg0x0ZWKuTDz7aEPAx4g4yEzD5yhym5xdhI7s+/vOEoANnK7kGl9rQEE9ChCDuvzS
9jswk6/6PNeUGLtkkn1ievu44/mJ6HT6I2WbKnGAZtO0n53U66XZZm9mdEj7O9oTX9uuAc7T3njE
aLRMhqnbYsxjWwP0sBAquCQJpxzQDWfL1YHHWEMiSNWqVXrXIAqpj1c6AI+M2QdjYPfofAkScxmk
HQDjbwWJIs2pUIfLKh/gr8P/b48ByZzA94JHrfulURq/2qYKKoCPZFnqeYwfvm2taVKzodJOWvoz
VKJ6Xe5ssWx9YwqVrlApsmbhcKCrNPxQa86VPYlKE8pLKn391hAfpY/GQ71aTSx/iBAMAA0ED7xV
xCzvPX4e+Mos0kqmIxkT/yDAHwh5s5txmQ3LH+vomTG5u2By3jRzzI9KQI+WxUPGWcCFcBC4tYFC
YSri1pCjuLlP/J/HDenWmhi9qpqFd4062eHUQmlDyUj4gxs7A4lrXDA92Ovgz27KTqQg8y9hHo37
6ROHz+p0gRLfZiqj4Bb6QASHS+TvymTZW05wmoWYCyJUmtNy/dOu3EfPHtCpOUR1HkFkMhkkM3I8
cpAqkbFBu4syRSt094ABPH4qaH5e7/d7q3BvHhD3ZI9FGu4LPPP6R1r4jgMW+wNM4A5ec9ZrUQF+
hH6vWf4HhmJL6jrKD4U0hIdJRrvglg8TU4vG2nKsVK3+TfptQk6m7b/edlnh85tLJTsV/4UG3tef
npFgHt7KgMT3GeXYFF57K0GOAOTXMd9+Y/XqJZwzUcItWPc1IybF9dBJ/syhZ7FaPv/y+eknbbGm
ViIwWYXKlE/NsSuxXj4NVnx9w1BCRaYJJuHEiCsqX3/st5zn2MaqwaUqF8wA7YHV5wSRSScnAukd
FSQqkqUQZnnOJUpKkvlPwfoBLknBWsOzeiAevrx1bU3FSmtl1SKCp4+pG1dyoHSa0WuJxw1nJIct
NEwhVOYG/TPIQCSorjs5vHjCjHqJLyA9FlnxY4zbB9jy/9/AdiFFwVor0Hh9b7dY8snZEp8yJH1m
jrm1PfC/y9fsqLD2/+IZcrG8KPsCt3ByrcNXwfTkJcheL26zMZLTLf8PzXtQX03dPapCKcyPFbNL
BiZGFXdnVhrexx5ufzMId4ZO/plRsCYEWZTMgz9mNaFtqkayrHcCCWzRQxnh7pofGO0FJHCFN0K9
zyx5jjRSONI9UlVpJJl7yw1xMEgOoKJDpsUGJkqUbdgR3RzjKXFOqrraqiYGQTICn2jOWxF17IUM
/AF1rAf/XTvL1qwuOQRLFZPOJ536QskSg7WHbiMMDbjIN9rgjQ7478Edz1hQKvyqyiSMdtAV2pUp
VabaUm+7pGryj0jmPK8QosQOLsAkOndAUbl5KhpqQMCQTxR3FZxXV5XawQSl0xhDr17IFN9N/dpm
jomvHgRvUPibHKX1AIXSTPzEK6z73VKDXBuE0KoPIgXPJt9h/+XEUiLrg5L9m2QcCMBbikD+J4Th
KTyVPJoYkiQ4j05Rae874b62q+06XZ/4rTZet4EBew9LsMrptrti9wrkUKcOy67D/Bu558P8aHKS
3VyebotSdWC4x+1y+IDNcJn4SdW3E9BaMEsp/HsxY2NNRjnhRasgkWIn2JUUFZ7QqKDw0lLkD3kt
Ei5nudjO8QGiHUcg02fr8GWGeUGMKXz1roILq3jXRf0SwCyf2+Tu0FgF4oGQiP3ZGOviKMVPGaTb
vQU1qFb4x0Igivszp2VF0v+q6vNlMaHK4LYy64iYFiAUNm0rnzxxsrZ1og2iNwWpHeJA8oZaKYRb
tIk54C0ERgfBYWgwDslDqVEiNkeQPBR6FjiiSKzejd1OEylEB97+BrsBf0XICSW+tAMsmoYofOp9
dorgdJd89Dua6e56s5Mz7w5upG95l7md5daW9P5Rz3oUSvYOxGSyDBfix//08o4xIjuP3Fdkoc0N
Xe2exsBssvOUdd9PB4gk9qrbdbLfPTiSFIRX6H+y+56r2F83TalCbuNpJ4jg2Z6wrcfpUVzMovXS
0roucSJ52T0lTVJ61LXhqbMyTDZuwH59MpxNru3vF1FPgs+n34ySrnrz5c5BBR5DpDprd89I4aXG
3rr5c0Gtxk2+MSEfMTsMOuUY3nGaVVHXOGEkEy1lqregvLbo6TjWT0Nm4zm9QDVyAg2dRROZsDDT
F1sNgwOcGc27Wj0jL04kr9amAlJH9PiWbiLufVvfSxH81YMq4VuNavz1NJgPbf77uSszi+cB4jpR
2X5MGTEkWdAlkz3I8wg+vIAJ9KB45xcdp6MONWiQlkEobS0G8uV1lhU08OGnzyRKo+m9JnQXlhoV
eydvaq2ugfAVaTISTufglaoFy7yRjgnR+UvGlEmOUT1eqvdMf1ZUsG9G8WWOVlNIp+kcbq9UhZkf
CkLv9rqqBD6BXoHi0tpjipeIQcxYYckT0JClUw0A/XAg767DIzhvIXaaj6sMpy6iMrBfzxAGKxWq
J5qC/qP2Y/djW2bnMV/9uNCOvaQ4rfk9OO/AHrWKoojHcskNrhZovdsc0kPw4SIQQdZQHEutpJY3
0Ftok9WbuccNwxt9gfDlT/eaHs7XoXrw1Baj3kG4AxSsgBxaigrzDSVhZa6Ql79H9a6/xjYpFiqA
EJyxOw9jHK87g8qaBHL4ZOQOM9IEfzOi4TxATACDIRrxIOwj2NfU8M+mQiRQSRWDvkwfiPLHIi0Z
L8KWX0OnSoBpS9nInPMjv4zMC1pH4WeuV1fp9zgP/pkyZn6+Ir942wiBTHHNQS6BNMzRnMKBdwm5
jaD7t2n47Je02aTu7Rxv023otdtP3BlGF6k1/vEL3BnseKEBWvZmvvzr9lH2aJoW+pD2RAMKmiuf
xVxUC/GGB7YQV/ov1S8cWz14D8dK/ejC0iQZTXOtiePokXij9tQH45/VRerDO3rsfMbY+lwjDRLu
12mktqFIlznNndVm1K8dfKVciEArW3II5okwMRJXZuEe0zHodx8GfWTyMYyXN6PYiHk/OEX94Mh3
dZHPPjukNtdZUOuMN7RtZ5cbMMTw7HuPxgUQYrp3tp6digvIgb3RmRfC7y7uyRNkZVM2+hTa5+4s
zH10xXyDyz+kT/1NybFcJVAGHtQywQoxLhcgX0lDy5OXbobsr/d3Xh+NoUFa+hdXEK9pBszIwG57
LsDjS49hICzsLo+79sgWInAsy2F1QxYCzxEwSyLBsS0iac1cjHCUMc6hzVfhuNCWRSjilIAhHDsH
iOGbstOoIZ9pPjg6uafWlQn5WenTAN8+a5Nc4D21Mpla8MuF/bV4oEyPP62M7YkDrT+16l+N6yW4
AcA46E4gSo08jhVBDhdEx4UDdLhHC8ksi5QyChoFxjn276qWtJJ+miNa76zbOMA8eEerSJ5NsUSv
Nc+FpSedaWQbdt9Ed79ScFIzTXgM6SJ0v1H4RPSVqsZ3j/zSJHuVoWB5n1zwo0g5qlT+cs8bP8kT
RK5qZfFNfF+jdJHpz89X1d0WizrurdrIm+DAnCMT2+9UOwru96BI1c48uZMG4pcAYXz8lP9nIRUC
1GykW5lMc6xdrxwJtGEeZYbh8wGzsgpuVQAZQaDBC4mOr3ypwNn1LmvTuqv82aESKDHFDYk+gbi/
cWsqCVVo1M0COthuwNwfSJtcssHgCqgfHVVp+xu8dF0UVkGNHvZcsg5wvfYrJc13A2Anxq5uWfzX
ExYC3dABShayydTyKPeJlZv/8gQedDbV+/7yjwa1vhAvlJu5+DdfX2ObUI050h7ym2ird4wvWFQF
LidIPFY73l4uxontAnm2yZKbVgtCQkjGe7iNW2qAddAkMpBWr07Vr0EGZrR4SMlRBSzCq/trpGY6
Yhz5gaF8FwbbmQic7VTzFXFX3t/kDhwstYPJgqxLcK9WeXs+CEN/9onTMeDlr8ra4PTg/reUPywZ
Ga+dObB8ChTdZJne4avch2uNhFJFu7UaLaHqGOcfM/eNkbaU0XAByFywU+f7RxuL5UKVa8iAxRIy
9WJkfjo40qUB3CbCgJYPd75n2us64gq4vYf+0toHkYhIRP75m3OD13+yGB6pb2SoEWiHKqdW6uh9
B6HmGlvKrygyqq3FRuyrbDx0wEGe5axtMRM2vKTegtvN38o7Km58noB2EF6JEQmMB9a6KRnus8cU
93f+LNFMCmsYS6DKCxGPD0hezE7BZ6M+h/+eLBSlXWl42G0ND3cEkVV9FJcreUHeEbH9s79aPRB7
UlLVrV83FJSQMBh3TWdDmr93PgFL1zNY+U0+U629eaDSLis4B7ITVgAdboOVZ72tTZriQblW87G6
TdhKRuWpRJLbdbO8eiuPl8rJ7kxOAo/gFc6SIEQVQD5UBuwiUKEQ0wUYQ0enw6LeEYf94Sn1nXOk
unVjtI9Yej2I5z1aZM+D0BJoKODdX9gMGevjEECUv7TYCddhXD5lR+qvcTkXVZvtnYMico2REAFV
FFyqXQ/bpbPHxv6KOyEGqVz40+oyGgw1js1SZqXPEqwMr6+vGx2ux3QvAOYsp3VLxhm9ATCx3PvQ
IY8pY/AnU+0eXMsYcvLN0FgqAiN5syNE1TAX/fuL1m/pI8cYw7Cwn6hWx3/CieLyXKwLREsrrIa7
cZcqrPUBmyKqVScguuzGurVsuVlbQLa+RB6krHOrczmXB5034+SFwARGu/B2IH6fyr9FojEt1NlL
P5F9yKh0Y/9smC9N7O+ypb+Tw7SZEa7kujLmD8Sa8f0xGKtCqje/RA35QxFN+Z000b3OBbYJx+0+
5i6e3KJpxIOtcZglVmi0nB+FoxGMQlOa0zWArHqbtr1SH7to7SkPouiTf+Ixrl/8mwjjrfGVpv4/
0mA0DVkfywZ0VcnT2HXaYS88VFLoqR0EniN0fPlHpqUQCyF+OylLrCc8px0ISHqR66zcDmzEIfkJ
8lqTvrx3oEbJDy0sbmmjmH3/xWPPZulZwtvCt/R6g/MdBdG5pMWdaLE+0mdI3Uj9t5zuzw2P79Ea
OMZZF50YppGJUnxhDW6FCEar6D2czqOc+7LPIsuvymlmHtDuBoH85wzS8hhrH+U2PxN+o/CKXpfb
RPyPcip44IYdCmrZfji5HkBtIUW6OiT0QZ017no8ysvLVgGqNiXSj8nySTbk7hZQixHczCHP8HmF
bQm0aksKjyoK7dMvud34Cle8PwlVXE5v/OjNuv5kWK14t7hfsrsQZOv8BLVbnm2BKdsSddMdMg/Q
9XED6jjNmaRhLegkGWoPR6RXEt6byFJ5NE3jU+UAGQLhZ68lMEXU4HSe1deZ5JmihfoJugE1d86/
uGin3tna5gGB0V8TNaCBbWwlw6KSqdgSzwS5JfKZmSNjv42bXLvG45YEpn+kOQFUhB+ldjhv6UeH
eWAyYU8o44cPDHssrY85adsFGhSsh04pk8YXe0j398Y1lRgFJELyWw/TB7CjZjwOiFZbLpnrSk9W
lMLXCoF2xCq6NQJHOvIEUDfZszVhzZGAtvijNcwZI7dTZ4t6Lcfyvor/ulaJChqLbmbC4ATKbcUI
GmSiP4WpSEF2kO6lr3vop01DtSCaSow0okLXGN4lMoTuWA5S4pmrB0kGLNYcEpIxYqIBe973deWc
44RfSbVmzJZ5RAZGc06EMxcNeA7vCZWVWpn3ty5skIJmTawWK7rPmZZrMATmNfr7KREmrxjbKeW6
i5P35me12asQ6SI2cOEbsWK0C5wvYGMG6KkhEHB/i+CTfWM3HslFY3/85fHWjsn9GHFHbhjwJB3A
dOTG/flIyIu90jqfTRJHYi+dfKNwQyKGOc6eNXG5LX1PywmLVPo8YlNM8qSBFDmZ6itnscE2vwkY
j2APm23M+jXGFVbyAWwZWeyf52qG0NtHLNwiUSS+Kp0XjtvtqH8RouMEkZu/73wa5crp3X1HjNlW
adz0w0CAUoW2ew3hLZnvKWYj3uhb6Cqyxf1wA2Sts0d4mpbXKzZmEJOTQSjDaCFyJP9bCLJvJ4YM
KvRc4rnTMMUxFHHaAQhnTq+NfOlPZz74Cdpp+gWSoxLx4Z4sqBOLBb2+npHqgUo1N2hCUKISnuqq
GAMltSnvzvIKt+LwdAwU7BU8RLhUpIExZKL9jYGY4hI8dNw4JKLOfRhLUM4X5VXqSZ+wAj9Je5hf
u2afnOQIKc3QtM34WOazs0ct/gQxiK151ZLI8kTFNOhT9Vhp/tHZJu5gbCq5oFOVhsO/4ktmbJB5
u0Us9OQT5PgVieUJZw+G1JnfG0bXoWJZCii3y9R42g6U5MliAAW+UTL1IGrC1T9jNSSrJgwdFXp/
ZEYDnoDfwU2ELG2TkrYdoBCfqDTBu6pKdZAQ6A2+JRyjWVGqAyPuIYNxBE7C5puWg3ktiSo/uP4i
sIIlDu1m/lGhoVSv/+01PxMAiJhi+TT9715KEbddTEqfS12UV9iSeM07+sPuIG3ojvz4v3gf+bm3
xKB+WbEnHeYVKMgWGRdmeCLp2Jpmq1wIPEOe4K95Gzoyvqr2Jd3BeJIJSIidPP4AmDjhld9oe+UO
egpn5+lFOMtqUB0+oEQZ0nkean+5CR1+SRcMaOTXliGwiGVr9xb7oMkqp4l+7007cpja4c8kuxOX
CEIFYMZITiovu9WKPKtqj0n2RCLqMVi8yuOQB4IxQmXBZQDb63Uj/rVxvQ/2bhc+skAU6sBMqJq2
Y5GzNIuB6hbUE1xAJxDQvk5KcgV04BhRBtxSV+y1H6zZtYMABaLLxupl800evA5DJHKpRFXJ4eZn
2hRAV3/UFCmycQedCrY6dRLaLuyQknyW6Dko+ZNlD156EEw0/EOUfoixYq5Iw0IS5Y9x4FJtFd6r
JmCd4Mo6NtAE4d8fH5y2Y62N+N7unF1ZOhM4vLKnLYrF3RUhnV9O/fspgKoiUdn9dDL6qcNxiUdd
fa6x6lNGM17qi+xN7Lv5BBqBj87BKhJkfIZeAm0jARs4eOkOsYMrMpsB1MlXlyCMJ5DRQVcBY3pW
mlIXJA2yt2GJPVRzpa6q5xZlwrl2coYcn7ZP03xH3xchF8hoHa/94QzT/4U80XOmOUwxQ4k6xuLC
lktCyOgc238ZKj1bKh8gkfvS6w2X22O1MLsm7hfA4ELAvhMjIqp0il2ZBxNc3a34R0xPVEhNSAzY
Qi7k2Jn1qzYdUcScBuAKrrlQb95Gcz+3UO7NMrIPYwGL5ki1HPHpKAJGiSDsht82So5xXGDi+8Xy
lWUJVMBWqKJQwQfHVIjUsd4/g2dgKkEUjpjpa9ggZgkki/YifdxgOrwGy16kJRinO1tVsrJqUmUW
A34BSV3gN5xDigJUjDC9wgXUvnDxpT3ZsmeJ+YPkfIiRyZ8P59AVZBg6+mR7N0Jwvf0N0NkeTym0
Gf4B9hYCxNUuh2M1qL2TK7QopY6zG/C8wrFRQf5SdR2v+q5q73Y7YlKBMcO9Yoa9KeOukRLwM/qD
odhoY2/5H4NMDIKrCzNyxbZTe0wO4UoDdgMurFv8QF4QH6JEYMMgSiuOJEPYFrL30U9z4blGijYn
r1ADXI24RhJsZOrx032XKuSmhJTodf2QIKe4VZXFGTZ5Fv53jKtIG9pEqtBSOn4aR2m0QGSfboS4
bTG1WOO/vVUY5zjZmtJIC2au/AL1N55AVRm/8SC79oUmcicbtunPoo7PPvaFILvxeTMpgD99NjXN
iPu7tOpbB51tjAfz56zISICuY8d2OIIQsoqNQcqOYXiqNQXOKPyOz7qrE8vt1c/YEwyGfoa2W/zR
oJY35uWtuuD/tEZ3I3szKoGk47yboHZ9UJ4KnRQghAiR0gLJ7MUwL5XX/n/cmnLYaN7U9UbaZIAe
zRVmWJnTCZ+e8QvmN8yJC/dxWsIyzfNxoS3qbjPpa70svC6DEP74HckneEhek/vWkPz7eCgPLPs6
21wjYotdgyeoCuQmXpOn73obmHAxYZ14mYkVRqtTaNnAzOh5GazXo41HYaI+sbhOLJx/Ui5vZc3J
EXjEZj2ORV5oNOosX8PULfUt2zxd6g4/Tujgf0PMKqgg2ImfJl+RRW/n1HOT2CEi7P9bNScy2TYd
nydaIPkswL6qpt7sENL9pGWaQE1tsvbR7s+ghT1ow4vC8jayVeBAfD5p8DC8kfZbmjf0H9zBTCdJ
Sqhpw9BoteQY5kUK8lAag3/iU38lNE5kXgA1tDEg85x4KjUCqO7StIDCoAPVWQZqiOKSctbT1ufo
z+3z/4gmdEK7Xo5lyUyXiJ3/vqP1d9eXQsk2Elqk9/MDJo6ROZWdXDMAFGElSToR2dGA/I6Zg8xs
hcDhOe2DfR2mk1YuDK56jbN9RabPqY3wF4EUH0lhjNNj1Z+r+HgS/mKDwESs8JtT47GMPx5/PlsA
OPFIa85hO331bV1bvWqi3TrvOD5q18X6T6Vg1b+YAVuRLx2j+4tdNoV8SMBxN3oXNkskbis+JWcF
3bAEJjylK830il6upaapsslo0tkQhy22HMo2aUdVQbFzG/bK6mhHu2mckfa280av74bNPK8mjENl
I4TsW8Jth7+J8AnOsNJOUh+76/kaxQYQhvB06jOLFRDizxdHzOGN/PjzQimxIYqQA7TSD7Gqfwxo
JdtppZjY9UD8XCxpU2054Jje+1JV47zveznnK67tN6jmziq8a91W5HIHwGw8IGjU20nOgEwldtNg
F5QDYfHpFb537F4X4jo6m25Tm+tzzmk/W7/UMfH60q3qTYl9M8KE2xnOMumjkGrWVvnGFzHXAk8I
b7ymtqcPrES5JRWmCWHWMpFhvTwhNhRlUYU+28C9R2jbxTcfXkqQfCa8Bx1zUKDEiy/vBEKGlkhc
QiLNADkriAwZhR20xM3ypGMYEGlIAgZkjt8RAKUFnrTPkuR2JKonSzaAmKc3MwIdyvGxUd+ufgKE
Wix5MFaNhFIcwPjAlzIpYQjV1BI5mSyELXSl8dBIoNsau+Ap/xSrVUORvWEB1Y0CvLEJMA5nuvwN
p+HZOSKJYTd4r2yBRe2XYfU1A5y89kIvCdTHCHHzYsQZGZaFs7pN8jNOTTPpKvpbgds68XZ7ltcx
Ix180lLarIhckZ6fKXRAKdiR4et3tVjQyIfnR3v3j8bLUKtHBYdbwfxe+MyHgXJfe9GH+dMzq9oM
e6ytpKud89bXZjK+jJUWjCMbToCVYAMOhmm75ce3/CYgdk6UjqYd4FEuj9dHa9+/o11TKytnUS7Q
voAzgozSGHlAVBoLIz/wMQUfZ1TM6tUZO1srKQRiIRfGP4VsxMtFHReCuXbBhEMMNPI73F8f98iP
aJyI6lBgIP9k6GQ12KyovFbiKul07pQzZQYUAxXcW1znKw++Jcis8bBRd4K2Oj2W1qpdBhBvXA0i
nAoWdR+IbUfXTj7U5FP3D8rDYahDKIvLpu9IqaVGAHXz+Ue4yYf8GrmPHPkb1um8fAV5rBOWQjk2
nqYu67v2jZ+KISRKG+BuobeMfT8/aZD86eSa23Zocd88b0b6WbGeIF0GbSFOAy5UHodiHyR4j1Td
fjLUNbte4PHsTCKai17zBeEzotWttmRtB8lN0DAKDGhzd21et5Zs73CQr18X3f6FxoYwa8bhlOq1
uwMU/Us216LY4rQ5BYfHMuZ6QfsQW9sG6uL2xd5E6pH3jzDMNM2/loPHNZyWvsGQjvacsx99wuTz
IOXubcCK8uXxF5+ircS2lqQWmeDuRpGzy1w0TczDogHVtYlnh9vwQKIRAfQAA/MzAEkj1CbdoEKi
KVFhDCw7QChPd8MZxa8y38hTXntzEGi0T58yG9mp71jkUuSUq6FHgYKcz+A9nRit7Tp59jmrNBQC
P94ZikW0OEDPSLaFAjVRkr6drP3qvZxfk+OwbxagsQGqwM8pocSORHqZGJcFRV/ocYrdXtAZGK+Q
c/fEhgdAtzRlSXuOjDbZHF+6KQD832rtp9/qZirzuENmaCBbHXBsg5AhT83J2/+Vu/KIXFcAPMWe
zn2LKZJm8FoHaRriLxupwsv3eoOn0WAGCYZaTlZHp5LxHhbcjI5auxl+ib4T166ZoavYpSB1wBow
e5qJLrq153mjNb2AGKpEf2mv2BGMpF7oXC/7M0M+92DJuIO0NDFBdVJvk6ckcbSRoGtovppLdXBY
Lar/P1nNFRPoannXLfaLM9QxUuhdLu45Hq16GtiBU364k0ERJ6+NFasegKJ6xq6c8UtdlyA+C2py
1Jyv+Xh98C1GDwwwL0uZhb1ITK7jqIzoLjDHD5kUHFLrPi7xngryXdZKPtXN0Ez2iu5R0GUu1VBO
2B9ihLctj0JnWr6p7wnE5SjlUL++cbUG79qsjg66jXAOV1aUImx5jIeRsIhyme9zx6SS2GIMiI8X
en1LFpr1thlL++oyo2bTbFMaV4mvkGgzaR5RliqhiBHXozE7hkRfO5zG/uWIg0Lnp4OA7e3+cu0L
CU95cX3n4soi/9COUfOAziOYLZ6vySZDXDJL50vsetzqmwMUylH/ofcMSPKQV1PMhMh2znb3Z0qu
5KeLZV0xGRg72Yt+NJPE0aB8SWamrxsIJBFUJCxjhDwNjNkVavqgUi7ZKMc6JkiHkVKQNR3jZ14k
nGWqPxxWp5GBQhPm1UZeDzDMlJvJxcCIPerYEBfAShTRcWV/O7z6Gwa1URePYMfy1axSan3T6Z+P
GhNf2I3hp6w6lNX37bBRXXiWWIR75nos2bTydJuNwTVlFG+T08rWIaGa2p/sMhulBWoa/L93dcaL
qG/E+tTTqyiTWaR8DfpEQ7kln8u4a6X40cYJPJlRv/GuPIhFB/nuxQ8Lisw8ePprfxUxH5R4aaX/
mkvAukzNWv97U4fn5x6yYl5Ta8bg/mPDiesI+GMrx2QJ44iv85gEqsrD/qJW6TgPmbnQrIW8hX5C
UsRvRnL5rJ2+dl33JiAzepGxnrT3z8YXlPv443WSHnMXvLk0ojZJi0iI2CK0xatE4ce14gUaemr+
nEDSjj3ckxutHYHhEILBxTwH9uiE2s4tQ7hVeq2Ms/brxlZ9+C3fzN0PAwwkqemgjyy1zVeuLv1o
cKbLWpsIHY86ACH4VlBMhYLPqgHj76mEOOBm4KMyfjp6J+WKMz0vJ9ByK8AT6q7wHz0gq2NXY0a0
jUMuX4f7s470idfbyVtcN+yfNI+/QoMhMT/pQU4s7u2P0B9xgfHpHbWp6xEW66wXP4LDbwRT4rTG
cM/2vr91eKkoNC/D/+3u8K1AEwKc4elL6n5OaaropleZfDsY8b6k8rBnHQy0jqw9/XEvK9DBIDhS
26uVnAscc/LPadVqd5wdNsx6XdBGJVHzU3OmG4Mm0YyBWBb3Qd5YuZsHkkyJfOkukDn17r4EbGks
ldsoMQIu5azvd1jiQVbSz1jb5di2hbMN5WA7fP0eVAZnQDCNbvsUBK0EvaevjmQ8KUg4KGQzNGq3
NvjC+1OWWEksMA1543Jjp6FyCFdhbwxxl6T3e/wdyk5LzRgwTG3sAZGHnP/A4a5w9Yx3Wzl5T0bC
TY9wXooX987TijPlebmdC8so1YcOHLKMqbo2bhNdjE+L6/eNuvv9uKcjTLU4rUWobs+XKrhbKozp
AM3/iOcj9m617hmfXF1LWSDhP9wjw8fNpa/cWEavejrdoUhZCkBeJUZ3uGQ+myjMZKXAz2K8PS8Z
c/YS2fOwJ54NQvMcVwxX7Q1k41hHdebxQHEwdEBZC80FJxeALb5dHbDadgYGp0X3ExAd/biOetzP
hE1mrBiyGgdObMz68fvQKeuVmEwFNcPPuIhGna/1EINwv16N+Hc09GtvBvlWmUDwcUbKicoeJt2j
nEi8nTha5KniJSPGwC/psFNE8MqBpZAazwGW1EHe3X9i7p8vZNSmGAnwc/xCeNEkFnwv/WrK0CAd
JOy9B4Uby3CzF0Jay2himxKa0HXeGkJuj+rTcC8Py33L+KihSadWZq6+34cHcc9jeCqyDhfLcJx+
jgFtdaUbtlxeonpLQKgeuJERwS/+fIZNfyFhxhHt7S32pS14bUegfszI6Xq7v2MpGHNshOMDi4qf
grHDem7KW5PARr3RPO9+cCUyyKJqUYyVx/5/UoMQRxJh3hQKDfV1NnPTIeL7KxCZIh4qPYSu+4YV
NX51oLglGHkX18OI+hAjpFmDeV8wrFbAeCOQ5KqCrUQMDA6rUT25+eoebvDLM2jPHpIgnOwMYm8i
PQ29mDk3z/tl7sWEBeVZJZ4w2sfXv4DtIHHnopk6Z7VJX/HhxKemZvAkKrG/SRyfGgCuGGqs/9+S
z/ROZeabJcvNX7+h7sbVxaQO2tKYkvLhwQvZ+f8dGQkVEO1mcQPtpphm/ZkfRgwUsrrEUZcN6K91
dzRlPYs+f1yU3BofMjAE86lGJq7T8FEM5v36vaz4EtYN9adxeb+J77AQhnOOqaODzIdJ5E3wqxS4
CR6NpgsklPZwwQiifnihTk7XwLXFB/WKd+aZRBGLz2aFiR08Dhi0HnGi6V+ztgnBitw7qs8WMi69
cDC0J0Pm61TB4BabAH3BwSpCwxYftdxFvkCu7jwsFM2d8ianoIalHwnPe/5toDsGvv1STaj+WP55
kE/OkYIfSTPWxTstNfosizpjEcnrCQVA0cQ5DOu8HDo/a4yG5GDIN7yCqsPtqOlxik/aH96EMzT1
rhCTQ54NnU9kzcns4dDahMaOv9QJ083brjqs+q3fErnBxDp01cNn0/H10+UJLUYnaf1/dkQ7bX+u
g0eOq5MxgpE211qCoFk/ln1s7tjbl2YC1IsVm1e3iyBf/tfzfQOduIy/z4rnREymUeh88k0nNp4O
YKbV4Cg1Zea9CxVtfUw6xBva6jYaeWQRyPs9Tr6n9CY/47o6xGUWIGfuwRvbe8m6VURn0/dTvwLD
XciXqVu9UZ4Vry/ZRHgrRXplSEvG0J40Uxmb6cC0KweooDXj5ejAt1MXyLQwBh4gg8lrq6BtHE+f
3oSNssV2Rt1/0uquA+XM9wh4kjWdIkxkkVkivuFUyxtcKhvaOJ2BoLdacU71oAyjj2pmOWwkuanM
UxPC5MkdWMD6rGbHx6vGStmOOyIl8Va4EudH5RNlRNhjFPqAF2fTKyzMoQg3qLUx4GK35Lb6atKF
UnaCIuIdzFrP9CpcHPPq3o6+a7AYAGjDJIeCc+tfwKC+M+IegtPP9UGtYi3J686CBqCrNsK3XNyc
VcdHPkTv4Ne1BwWeT4WdQ9/2m9FGRbnqr1ujFWfGleP3Bl6Wv4Nd+65kDCUNFpKqjBr1+/oJn0QU
oE8zUFVEoPZrz+0phOrsa5OsKlQhhgAyH7ygBEtdjTY1ygXN3l6/sPs9dzpRqaBRbQi5yZCs7kVP
bcyG+Ep6KRacoW7Yi1Op65I05Fp8zaaI31mmpKmDQADzr1V8tGxxwKZIXFdsU24lt56+hMs2bdRR
hmx/+esj0tAb+RKygRFEkazKllPGAuVewn8Kr1+6E71Z+Ps1kCML2I4R4V4OJgJsD9p+MJ1E3ktN
DjdbKbLRAKF/lNgMf/d3uIT6puG+6k9Szi8gux90ntQv+ujGVMcWr4Hk1tp1fiiiY63lywVSkQtM
pzWgSyiXLx01M+j4SUi+3IbyNSAmCcN6Vt6RVWIaItAjOKfj/VJyjAO4IBG/Nm0rNLxVp2vFnOaL
VSvQh1zi77nxSqxeKQfCMJHQFuJLetZEwpqwnvEVG/LUwEgnGjMGpEfCTVGnSVpYAYcFcyUQPe5S
d9nthcQWkbOgpeoGTfwnLz0RTnEOa+L1LRecNv+KgKIucnt9lYtFh04MKZjv5yYXU+qLAnTAdq/Z
h5hikoeUzs2QGUv2V2ve2EbDaBSwiGbkQAPFdywAHhKCoeAeDtdIsgilB57fvaY0HiaWN/jPL7lS
BI2Ha2zK7NG48m6m10nJKRjjE7e6m34P1yu63ym5kct8kOpsk7xkthgOGrYRAfMAYXapUMZioqQ4
PXgCxbUlmC+ONx4r4Y0bsI6+Y52E8IjavssdUhs5T38acYFiKuSGLd6FqJX5vnyluPQ+/JWYfyU7
YCEpQuZIybbEjPfVRYa5S4647sPb0//o+XZYf+pO3U8YfKvTrbLg7H4qVwitLiA26JYxGHjhFt+V
MHoXpOykzwnQb3UwyNDcyN/BHk/rY2rt2IkDZCKfX3+SIbtCrur/F/+D4u5Bwtlrn1TW+RXR1uAQ
lHr9idzzfpAzer7ftL+7nxyDrEO0UiY0+0FumFjVboByCKtGvx/7d470g/MYW7ZPrzx+lTeVn9C5
bZkVMk4osJLEEkbVWr/jw1yX1chw1MyZBmPT0q3hRlOlWwQnjHRG8dvLFpeLZtqz86gQ3VNi1aK/
nayMdgifvuRYZgnBjZlT4ZvTUFoTpJRgFlCu/E9ESktQF0UeQavlzxpvvuNzxx60F16pSoVZ/RwB
5bONX3lW5rWb1oMoywBD8HqGD3K42k81JztA1clHfrhpVNRSK9g7tnNn2Gqqv1uJup3vnt0VALPe
5DZAVoPh/LYON/AwWMVVtyJFsv6+Lt63b2ks1Rk/QZya0INo9QYnihilOAHyuuysCeYq059nuS3j
aTiOCor32TFb1azZ2NTOOB+VwqbHwr3yLKSRKwbVeTDuy2AVzUO32rIjSkFiK6tXGRnTsw3tkDtW
jq0P9cATqYLb21+rgw3fFEHxzaNmqvX6+FQbbK4OHbDWKDmWTV//WjM7wenlcJAD6zsLmGYFymcs
MEQQ9Oc8MqG6E8ZAI/9flFqni5+dut1KrE1psJuD09IhVKW2bV7QgsQD1bzDwF2OMYxPJzk08d5g
JB/HCy/jN56UYqe/WQ2hA6C9573l1ooW1N0eKhrB+5mBWvMnYerzSgljAu0OwZzxc4XW/o7UK1HG
QJmSANtolQ43mevHbCF6voQfEEL63WsKdexnK9BTE+0nzcAQ3Q29GxahSxaRiMEYVpeHb5ylPODa
LCvazpbyBw76iR9zVOy4qyh8e8uZchkYKwGu39kP156er7VVKzwX1vzFp66pLHocxlW/ibrFUNQ3
lE6tJ5Y9PFf7voNl9ZPdDsSYPn335rJw0LFygFjIzhEzbycSIixzGHA6FsWFIvtsjITaqomP18UP
u9tKirL2eQWTfe0JjPibn39nTE3xp8YCwKa31pu0seDOZVvMF8zCjjrJRqb/aHmkjmnx8WoXC/ys
AT6yNQx+dXAGqMD/W9T6bRy6la+3MpcRI9VdTVsBUghCL1W2O2X7LVrS0xj7KF7KQnZa2ifDLi9C
0SHrxn+TiaVI4IhousIkfkMsnFZOJBK5BmG8wn6V3fPPQ3tEsVSs4SOVGyVECfeHDTz6DTPkeRlT
rmMrtK/WxzL7Lb+N6yT0h3tR1hwkkP2gSiJvnGlm3MbQHJEplDG5uPkDsTHG2CzJgmPfbGlKhZcx
uqqf+R3jaMEt4BNS792DMEKLuIB8tlBFY8KyHZgWl2BjZ7lejTrW3UepEVIRo9szp3vu4jrS4LCa
Jngmm8Wt4kbcTtoJm5sc/uVygF0I1AnmZHey8flkNMgvJtTF1OCUewJGOwV0h0n1BzIh31ugxPYE
jXR+zaq9W9Ke44/ir3Upx3yMxMDaJriDdQz6VC33uWUCFqFchIIFpvdRHDU0i3x7aXdzWTfZolFr
okeQlDvVNaBMAg+mMPPhAbFjL7utzvZt6v1jOjaU5Jpl+8egxciDWvQZzxHAZ55SFOmMWrPcV+Dp
LVzR1dZ7QwG2RHFlSFiXMhqBGqE3C19CTv51jbWQz4K+AtLpKOkqY1rF/dZ4oSQMfEkv7ZAk/RmS
0g+f64MoRkxW9pn1clvkwR3IiKz8dAlZHx6C36dwb3USeJ3rZ7U4NXMcpJHjW5uiMSk1GSa/503w
t5w9HKWY/9mCook7igRQqK21opMojBn5bNUJP5yIbMycBO6iWmpjWPheHIgP6bab3WocqiWgsVsJ
dmAlC6mI5A0JXZ0hIY7UShsY7PxQKh2TSXl7Quegnze7WFSeHCWtd1wH/llKr7WYRQ+Tb6LCd9U4
P2NMhf8iuE+l1OuALGTdTIaWrCdgY06kguYIoTP1178zRrjMNjEDBNzMKIqHD1ebulDrQKU9ZvFQ
zhakhgaZcl2O19ptUs5cl7XemQhlDiIg2/Jca9V0rERsuvKaqcmuzCZdTbMU+41TkECojooSlI5F
ujnnsaak/Fua/L2/VReEg+Ia3T8G5oc419Vn+jTSCkEQ6Vzb50iGl8p/7Ml3C/t+zwwyjQLtxu7p
UvqC/tOCHJKwDQ1+7N5qpgBciX7+HyCMOL1ZcMx67EVZxNLD0C1m/MLZUlHySz1ghnPsofQuF3jG
4phNQ+xiHdD+UtYhz7hXzZzxCMHiBi1J0jRN329ETMvHJKqfXJoHGsnOIUZI2QQbvLj1IMHIM+ve
UKa3FsOS9HyGncem8+PqweFLYSC3GC2K1QHJq2odj/51V89PMhjYKMXFe8e62/5ijMIVo+gPLTIi
Lea/17oOz53Bx+l4YmkwKZfLSben41WqMzJ2O2XgUr9d/2jo4KSpFA6x3VE6YVJlgU7Fk1cvV9SY
7v5RibooV1zJTLwc01OdBUnP9TRxrvMO5qK8HOKZmtEhwWRZvVHD/C/utnCiIvE6ydAg+ecn8QpE
LpqN5yh/A6L2ZZy9yauWUecKrOmv4R6HzxKVbw6Ah/0xz7qstrEYPXHgKsNmhqQ1cPw9s3RzkGYB
oJPKzzJS1JovEROh03alukteZD5aJUsnjkXKT0TW6lHVOZbtR18Quf08SXLhrpowT5Yk7oo/zbOW
oDvYXsGhbG1tfy8qOpkZ0o9axVCP0fhlTi+I5SLSXURkn/sOEFUzzT9qQuc/pi5HuYL4bon+5aVO
yoULY7BF5MCgv9l+6ND1xr0Bw6t5Qnzhuf+JbCH294yZ9yHgnG/SWpa1+YtmOMeTBU0nhnzOCWu9
7fhghJK4zRlV8w94Wr0RdF4W0PiekmjGwMBqv0BWk8CM7FSYsU65PGmS0YdEwhoLdfRiVnKOtpti
876gKbeM/pliQBlvwRKcBwIRn3Utw17Sf43MVOJAm9as/HQ0aGe+kfQQOoArqqjXVI7cwejj+06t
G5bxtQoioBD6ojx/IjsTYveZHpiXh6OoLTIt8e2te4EIzxr80kVvl9uUFykBUXLclFnKq5yDe6cY
DCPvJd3BHWODckAFDLxcizUQSVA0JHowLObun0D6AD5A45iAqG27Ol95rn2C3j2JkL7CPg6gw+cH
4n4DH+yWWVKtzzGzQhx/67bY5nmSiHiqLucXYFvtynVvBLTMKgsg9XSKyZoGDf0DogJ0+wh/depf
m52cfQ9oGFX/TuRDbm5J9lwCqTm5dmO73X1XbGYmyWWr2yXstkLhhs8G7zKorUNu4SPkBrwH6CtM
CWVKQdQzr1AK3SjnKEOYpaIEmDX7BDwyFQiLlMCGRByC8VEpytzz6G6+5eywGjhaZyiLNxU2SdVX
YeZFsHc67fNTJ+6K57mo83asz24KI++WxPn0YF6Jws5hNAx6mnMgmQl65gR/x5BJuW7e1ppeOZfl
kxWu8h9vPcolYS5/DcFcE6kZm+9Ar1e/rkABdttoCY5WIYHh3wTFdnd9qQAb2oYt+qjSykR+1DP0
z6lVCPTX62AjsONksR3PH5PQBvM/uSy+V3hXJ9sPZCirkjrOESGdBEbLPTyfsqeGmVs7A+srccL+
G3m10m9g2iEpCKtj4zBl6tFVtL9ZP46rANdhUpsdx7MMk2RUpecimQLyS1AxmcMlLvR5aBjqt2KB
HQfvxQZanHqaoxfY+rbCF5SslIOzuT7YiYhUBDQXCcCNsGCx8IAV1BOXEESOBzLXMXhqk61Wh68h
CrNKINEm7itqrZ3Ay6jyRauLBoxsExvgwOd9t42a4i9yVq+vzBXGlbgUG0apAzhTIHA6Wdj8f4N8
7lIlijQlyJ0nuoBvWsJ75MLHF0fYvsovddKmgDafx/6okK3hh8dQlTT3kjPvjEEpxAWtgcvcJIr8
FEggANdFVA+EaXvhqv8GKPblzCAiDsFghuXDKZ5CYBJptVarlJ9eMYHrmZY5MgfJQ9W5al4A4das
3Ldndr3Z3YtcErQ9qta27HPhD/y8u0vn96bfRBI+iNsWyzZfHsAligaNOZF6kSHb5sqHwycIsxfN
LxRFmXwN9yOOA+Z6mTQwwuhxQhowQSpqv4wpISW9o4gDrcOy0A3gUkgHagFoZaso2YjSCxAk6tWt
+LZwxIHBg7hLPKU50ru6loRDkJDOcsnrrKH31C+R87SX+k+xgucbPBic50pS4NZmGIyQo9EBkf9B
y7lxRxJ7iKXH2hGHXiD1XJSM1y8x0IBxYeJMc95lsfZwR3AfdSxpce8K9DIRrclCAQFL6ZqmEgKu
tUqk1ANmUJul1XIZ8StEJ7fAATEAnZM2J6V3E3UyU13+Wl4DGAwWC+XzCJicasDeYHrZ2YP3CmV/
IZ0b1tHMlzp0xB/EeTLSIrRUFiAumc/xAArRxWyIv9bgy/zPuFFwkpBCBxbNtilKdqwBn4ipTTZ1
pXKjgd1NdUxNddPaKq+r7IAez+OmAb9B67ZIojVOrYgWT8VpYgYYIHreM5/9kZDguzpnhZtT+qsG
BYXgMznCGuvRkJa8TuJFcPMm63oRZCLWFVoHt2wJI0qzOa5EZrn1E2d55jlK/zlDqx4Osa9q7OH4
GtMv72d3un4h63O783lt9K+dWOzwCitcCofgPvywTET1Mew0L6y6PQFSRgYJeFnQSbiWiJr6jQ4V
okdBnrpZRV5vhpOQRwS9h+EJqdKB6k1OYEFyjtPLkd8/KJpBBJ3xxQ4sAJYuG1xgcPXMrAwrIUm8
hPxYcf635xNAtXd5wLcXBLRkmncw+Cf0WN7DaFtOPSNjKaxvz3+WaybJmfktbHOtyIgLA5rcH3/u
Ha7OlPszzWHkLLdoYWIWPLzxu08EbLUyx7S5+dh5ioep9AW9aUpD/wGnRUF4+G9zBcMXAc3XriCR
lw8TOR65bSixbkcyDYRh0Rou61tBnWI00myVUu9LlU+U1YAVD2cWRxZKWQwzaEhDmd2QhbmJYxtX
AjwflNoG7rHh0I82r4ycUolfQjJAmbu2YMfdYfhJE/3V69Y707V5OTQ/GkJ1Zhv+dIxMbtIAXo1b
IPirzwsq66XoF3ADSfqBIvU2korw8VvI+Hbm/+CbcSWkSeRxzIyE7mBI1nHf37cyqS7ZGuhEHQ9v
tDMiwOkWT4ERLMwvmPM52XDxKfPpCyUoMqnVXSw0gqhoqolA7CBmS9RlfE2+g7BPP2cscnTX8exw
Fjna53DjcexbvhRY1bMniCdkENKQk6i4SGiRIPvRkwg1YsdaJKQwdjm7QUq+MTSGmnJPblFJKWPO
Vzvvff/5JFDU/ztNwLjXRZ5xfU8yw0cPiPyfTowGpkIPq4vOMGJuKBeqBRuPhsdcK9dwPxGeH/fN
NZ9sWlHCx6V7WhYvCIy+6O5nfaTUuwmMuePPOib4mnvdHxtwhyxhOd88clijExQx3BmWsFvwo5DH
MkHjw8bR3EczBTaHG3pkCW3SZkCJaUdgcJ00pM2UZpIBesQ83O2RkWgRU6bCtVgcJ2B8FJMFcspm
5Vdo2fCfygM/bLDLZVBVl8ruXGl0ZnTExEL+6Shxl2SlS6B5tHCO3tn5wbQEavGrSz2OAsMLbfun
FHxyeMeJZQ0GSWzi30MiYrNQoMl7jNwEOpyURt5aKa9xqjiiDbO1GvqMPN4ZpKfu4hXGf5jkhd3T
8cDZma+bTqpomp+ywTTQHHQeH8hpfaVHGVRyq33FG7iR4zh1nwAWukHJvYQN+TJSPTN4x5wrV6RE
tkWCF9+xR8ghZ+gCkuYb3yyjgAs058Z4oVmc/2H1xWUMydIxIeHzmCZ8ppkWiNBOPfx5JlUi4vu+
b1iHR9PD6TyM8fEvGmEzPaVTXYJX6GZUaaumwv7j2xgFCJzwBqZM5foaKoYn3o2uGh6f2rjWMqRQ
g4FLSeydwoixdAMyoA2gXBgZAOheJMMETkeCQJqNLzndUxYjFfhLAFfpA9z+F3ATX40QCHBdIfbL
nuDzSVjvRz2J87SYgj8XwRtUhclAiPsyQjR+PVDXPNAkfieh4vQjl2JA6bcf4BBZ9tNxXm80o+/j
cb6GZHz5+Z9Uexoa1VkmTV6UY6kJOKL4BoDArPqJmuI66+0/XkImyww3kIssFsOHISypnftiGoL3
7Y/+FBtit36h4H1R8BNKrMNPIOit3LZ8MsD2FpgzNz0XdaHSqfxdba/zMHTEyvKBWdDqQzmxiBuB
FVZaQ+C01zHIcyg/0vdgea/uf9N9qhOYiT1DsJ3wcAAoCNNY3A1fr7h69DbR3bZAITR3HHSPg0PH
P+QVMZwRRkjqqZAos4Yj/WVNVfFgC9IZwMtLbxmaJo65Oomw271V4dnBR/07daz6+rKKRpLOOMkZ
PJMPl3Tey1t0RvSzjspTvoa3xbjlF1mKj74gy3Cwx0v/MoXwtZdSx47H/o/aIeobjrTwWmhmq2In
G73tUlceIDCbiwmZ7gf5INCfYpxy5YBJpu8aXHM4MWLUOIybrN7luDjkaH0dLYqNl64d+NoWSZyy
qVuNAcgejYTauDxBLk/jw/adDCveOOy39bvPwPWeK01oaXWLNZ/gcpJxIPzXRY17fMB6fVyB3kvi
JAtB1hIKI5vRgEscg9GErHPSgRheIO61pjnHSxgEt6l51FeEBhip5bQ8aDsW0LugdVLDqgPqmxHX
llMhmQtC8eHlsA3faXU8759P43YKnwymVkDXPe84sK6Cc/gNAtBd8TQALPqcwcEFpRlwe93vbsaW
jgsbYx3/DN7SF+fd8k596WZA9nirBHNEs8du+UcxL8dOujWZBXrO9bARt8cwAMfvl/kOTJ8X44nM
5onmA9DVbljFUM58aV5mr47rBmFyt2t+zdnozARqcmXPxraDyQFFWl52KnPIS1L3HhzUiZTXU5gC
UH7bSOTJmVQ15n+ve8/F3rYjvGas5YshgnUr80uJOs9OkVnn/TamB4L4etKAWtsPg+RuSbObXMNG
3fnQAthFvJtxMks/CIaJed5hlNIVk57VgP596sK3E6l724DnYrejTG8JfyKuAUjjCKbsK4wIUkGc
9IJM4fuJgo5JEAXlvfH1QUWpNMOwdrsShHGn5A4sqwY3OZagkbc8FEwQh/Hivf6ECIf5QOvXOu++
dvltH4aVpXqdmGB1j1zR4cGhgwxGohtHjIGs3O14VU5jZ1q+SwNfL6/8q1hH1tKEErgrVxzqLl8j
wGSKeoWt0dQTGwBQHNKM1p0P+9Rvu4YtxgcKOurxrNBBmH/pp5vYRGC/XlWCTX9yYuJ9vhv+3CNT
GK7g8RJxkpxcndfYyDhBptc6ygeyqy3b5czj/8vCK47oe3y7Vbh4j7GUyw0YOfz83GrttXmXBmSX
2p/6vWZfXAftKT1YZ0DwHtPUhefrlHZMZBkCN3QmRs4XxRebxKLe1XmWe48U1LtTIfQXfhBwXrNv
wshr+EYqDIG6fda91kV5qS5p2B7TLyhgMsuJE5WtDenME7TgL8qHRSxep5g9m40bl6aLiEbahbri
UsUy3mjeMGwwixfmnNfk3Rx8k3OeVb6UIX3RRZd1wSPwRm8NROEAG317yBKG3TKmBMClCB2+iwx7
hO5PgBhOz381eO/y9bUOZvCmW4GMdxB0/RqnEUyHXOtHdP0pOFbw4DyzCWZWxVo4mhJ/K7OxIg1s
1seNtEkBiTFNl+F5T7RF4bleiwKqgsb3F0QgY2SNdB9RbXMevrmD6PqpHSoOitTIPxDR0NPlYuKB
uo2Tof14D6ncfIKnaRr9HqyzLoyTPp4qK4iDbtfJf1QyrT3KTop38O6ZDUlPxKkOHsCyBiiUVUWi
R85NhhfrpWV9nutdZtTUSq25rkXHp+eceAHquNUJ6P7I2ar0gsm0nB6S/tKTGdnVCF/HIR824Yol
NYMG+TMsvqqqxGD5sPnTip7bUjLRXsZgPxmf7mmrutY2SgHMjW3n4np0QhtI0Xge46KNPU0Zvkpg
6T5TOpl0HWe58utjc/O/X3SRFZERY32k7B3pcWTOWT3bNcz8tqQITmV1fHtZk+RQ/fObjDjSOsJO
RhD5cEsxFrKWmpfWnsISMZ8y53pzUS7/FTvinpNymNA6NTx5CYOP3F+g9xTYh+zY1HcZi9fpcNv6
2sq6akl53GngNUNvBLq+vr4qmFZrpZYpR2Q+29QRWGKU1wvVpTMzrC+lW3I7MAZVY0fg7vtkGAmm
HOEzPiStX5hNd79t0fjekwarshj3W7Qo9rHd5p+I2DrisRJqppuC8Eqm22iR7x2DkU0yKSmkR8Mu
xMGNNvzf7F76XLlc4L6ulV32UnBtU6r8yLlVfzQ7xcUhF50jsxorKAEwjEaNM/OaKXCMpuOoEaD/
pTPDpzzX59MoCFvuoo65/mq8ZmMZ5x0PwWhv4Lgc2/g5VB8+lyeSWe5GQ6omBToKYy5Q3msoH/6F
7A4oggTfvIk4PjDA2znTNtoon4zjNmGVA24Xvz3fUWLHt4DDIpyUxd8Z5ipUWhLAsC807zhZ7RxH
+XeZDxBDHTY1XXeEPfe7dJ1n8NPKPOUh9TS+j18k3hK0+BMLaOI+i1AJTrMeBb4707fWXWJz2lM8
u9biZ2+KzktHSQ1raSY1tWg0qDAgx0Ic5NO9zFoNc2kWsOU5WY7SmtojQSSW30PtsxTdbuVvph9X
abrj3+x5DTcXfYMVO7AxFU0qRRSGZXh8g588eqAkJdAZzxT3dPXbZA42CxJhHtAeA+PNz/ePoDf7
33UEaFPzEQEKowSr6G57DysktebnevEtYFNxpi/Zc8on/RX2nOc+TPpvlR1Hlhc2ViKannXN6hV5
XctFSEqU7caU5yc7od9QRkcIVAV51TvvGr5ASN0kmteVXUMBrZyWooo9gQ5m9RVt7YXt9wd3RYJ+
WBmjcVLqXSYvUhhgT0VXVZXAWkyE+hXckfJsA69SXbCshEorlvGSWFY5vD+fL2qtnm/x8VHZOPal
HKjQlEz9ozY3nML8hFcLcq6v22Zpi9s7WlFF9TJ73DVSPF6FWxFCAlVUdR0uMvuQqt2uhjGvbIE1
GKEo7+cUbxLTxvKxGWbFNeeRtnFYARpLmU3/5NB70ZrC8hpPrQPOMlroLoWg0kQTjrzA4CbgWJfD
13oeZbUEdpOJ2gydO7LKfHcVCWMiMObec5WDfWWnH4HYeNYpuQgZ4+Tscf8ofePaFoXpdFFLB9nq
evo3PXm7ki9kNzqrcRRE1HG+wlz5nC9sFF2KMSHK8lNdVwgw3/Mg4EOCY92ahZu5ie1sx9Grheyp
k9ugY12BmGSftYIRE/xrQ0wqFXeQU+SjcRELmNlaTIFu0UUSh02zanb9S8AzxC9zQQMBssIoL2c3
+VyeBW0FLPPyqhIhQOS01qSUFCe8OUYpuo8FE0LwpwjWSxImJKF562w/Fokw8HuaswHNy/X3AtYL
GznVq12Peslci9JGK81tFniKY/upzC90/X/QEhi+diFrjkmew+ASdi7W/tmG8zwdx6xteZAt8s2v
34CBbFH8FWMkjPUyGivPv5hLbSvUWe9iI/BKwbj396/YvW7+TAHFB+gZWT3jYSKGVjbnPNmGNQSp
Ot0YAN090vu3pWl7qO0SAz8rK4JWwEquyyPQeIpfwEwc2awV29G7u/t9eNbU/6koXBFCDfZzVh0K
eRKC0CjNX0whLljmUb4dWLhj16GtWUDKeUI+hhXCh6eVeuSLF4dAxOgph8gasUL0sO3el741uqNd
n7hkxYV/4Mndwn2b1E6pAhVxgKOzGNU7b+ysraNjWXCfxoAKxojKAxcHcKmW6DgoOPn2UbNWoa+o
8ijaWxngB8Nc2j0TM8Ji3jxgl5MhmA9hmMlXtMHGy9VD1VJc3lyPQQ2QpQmbzPG1Bz+nfvMsM5Ve
B/R1I/SXifKPdR0ZXp/LmfKvNtRJcnGSb7aF8hYTuu+ZwF2Mln+kTKnc70hrTcDlqKItv7dRBzJ6
o/BFomrm5vH8oh1YQpu/TMlPdXF42M1AlxVtXR+lFOBYZZ1DpHC2aPhZBxImcXM2rvodtsPWAk/6
Hadi4teBXG2vOvwmPAfAo6QVRXgmchELQK724EpGpUw4bc48/eKKCXC0kaJaRK7/c4H5V+mLiPXU
x7JiWV8wZ30bwSzeWSoazsfFyZi+2mn7a0z7EH6DgE6MCxa0P37G+/eAy3TYyOd9HA2dTLcdl9M4
tdAu8ATa8U2waJK5fvb6aHzVSWHSwG8zVrEW5mHHCM18EL6bYZJKgNa4EAbJkHYOK41FAip9Msbg
1YRrT2ozEw4pB519YFQ49jGucKWgJrOWX388rx9abtuoOQzolu4OuwFY81R1w8h9m3wIqPdVperc
FsML3IAxI4UKFGRbK5IH4PJmkcHa0luV2yWlLVhj09Syp8FzCYH6crXMFRKfnn0+lSd/BTqjMYPI
4ZtTt3iXkE0PGU0E8Rpb4l188FpaT13QZKkFgieNt3gdJfOApahawqZj7OFG9KMu/m6gcSVGGkMX
swgjISFNcXu04BKUS6yh1C4hyBP0hO2gHRI0Igdh6FUHtiF/n0MneGwCeZD+u+lQfbAkLlfNEpl5
2qx221ymZoeF8LU418FIB7tKYjrj5KckzfCMwGFH+ZWkp/lka4Im86GqEGLHp4imBzfxeS7Ogeic
jxbklBhlRNyIWIE6+45PFPlsHxLF/5QK9wGxrdNVtpGfBaOVuE8nk8fyozv4fvGj/WjZ+ooB0qNY
9Qp1ov9Qf2NWYtSFW71AeeZxE9sSjzd93KtpowJPw88eKH3i7JwHoxlYF9lzEg0RKgyHb5WcpPy7
72XZWHi/28Q8dyps1Bm9UzwFqcKmy5e01dddWEAEhqLhqB1YHvgivOsGMAlY2q+0QBGop5dB/74S
yJd+M9+WGKuU/5c2rjULSTOuMo+bYzqWPpNq71iOF7zeyIAR7Lj2Z4o17uqrLLEGZrQgrGhjWH4/
qVnLuABWG52DCF9bYN+x6cxGTIwb359dK+UO3UmWQcEBiZdnzSm6SuanExxIIfpQTdNqzricGxA4
8daNrClbmtJdRDCQUtW6WTUYc9DnjyOxnnBRIScX8cGo8l0OwQmJBOKKe2Rr3J1Pjd9x5Qlr1O/Y
8kQeNNC3i8Q84mxU9FRKDFLnFrmosq0PbcCitkkm/D/KdpOgB3THHmJIrHHleEDMGrVlc5Tn47Dk
kt7yH/pl7rRMYmU1DpGRZGLRiuTiURTvVASuVsEP/aUc+0z1/AjpCvsfIcKeG9CDBnVsZnQ06syg
wVa/TlHs9BXxJIxeb8n85rczLQG4x6KHmDtnJDrmD+eZE7ksxsmA0+LYz8AZclfcQCPAFb/mqnO+
H2eJysypO1f87owTCclIuuco3uF7C04LesoSd0oD3JVo2l196IdfCxkNd2Uar4eKle9jBTmWhfFV
8eGsTZmC5t2sa1W+cQjmiWnPxwu7TMK3s/+5Fo24MjlV8/PQfyJIWBGzUVzSmjjYAHmkQGpuyh5R
J/S37NPLbwhRr+otL5KyuaDj1vr+QeruoKjj1VBnURlk6eB3OLoDnkCKDqkTEJkUd2gnzmYR2Eol
V+/R9EARrPdAl4LQbnNSMpwZKTNd2xr3Vs7gvGrJcqPWQsG4UnyPvLnVobhi/t8Ni2TDKIStGDbI
1Gkwh9oAlX9wTZF8EVr2bb4ojAZL4t8DuvB+pZTVNZ3YDSC5fCxfjGawvmVypwyAGNIFxBgh3PZ/
Xe8Z5XRysZqd9q/cOQ9M+irko3MSIMn4Ar4VHuZRDQloyKjOi/TIpRrGQ/Ric/z6N6V8cp6Lwvbh
OkwC7+9YQtCU2UxkYpLROOefeGyk512x4zIKPXCqOg5eppeuaI2oof6YiAiN3WGTa+yoSLTIgNy/
tLUE/GNKMGNaMdSp7blUheVMbZRIj0rXE2g0RpFMh+pZ/X4aJe+h9WEl2T9USwCo+RsEWICzFOnU
wrRGI88CgOMT5BNmllHMdQS8RdLF7TSVQ6Sr76tYI30IVX4oLh+ejDEBhlddyzlLRSKHvefVHzKe
LtKtBG5QRVqCQCo5NgpJtabkaNUY2aHlcsFs9/oAnAHtoMXKGfiroosNf7Qbk1gnkJ9OrC/rsZEK
GdFnMVGGWqHGtFWgk8//gohgxxRJ4xXFb6WrqliX2MzSH6PHlrEZl9K+3CGR8rnZCR16pIGW2k5v
44Dmopua4Q80vtiSQpEO4EAowWcREvvkEYW/ewW4bEUB48UXTCixFEX9l9o+mQlxoECO6NCj7aoa
3IbJpoBArciXNCLoxJUscopL2ERxZnH2Ert4JqNS7jj5TpOZC78fpk0+fvklZdXivHafcwn357CY
g5kq9OYlIPhcEKwoksE7RdcgSvO8+VV+unphznjnG9U3Lwn5Buc1Kupoa+oVuTHIOKkRr43Pi3E2
mNwbOo99p0MWVKQMTZbb0opngeszyzFc0gTq6kuDJERG0Gsqui6a61N0xOsKoqLDhWrsJoXH47A+
OQ08ShtCmILBIQMpO+V//UDKhKSZwjqipcpQ+o4rlb2mqvynW9A1A1SZj2dmj4MxZBQlJhOWX596
6HL4IgtAO54pCi2txxiDUwYpIKMFCF2Ig+mbIK1h6xq3CRYRxQbLChYl5iE/hfAfExaHhRdWCY42
vcwidQWxJ3bChyrApgdIRMoHSCVzFKozLi7IK2M20c3IMgzCAlOl6kZOkS4+GLQzRsMWnGsxngch
anGACyJl1GmcSxrjTPRslXlT5ZPnUp2QKbsfVfqTylL89BiVmBm3mHfFFjcM+WqOsftkvv5QIPcy
Imd/jxAra4veF40hYp4AA+koRnIf0jMFPdIdPNHkvu3w5T9bVz3++BGsT+2o+wIvLQ5g8rA0wC+n
YSgTKAw8mKMGDaDTUVoKKwIn/+QhwthaSrcIlTrc+4EWvYWLVjN4l0VUBwp1sislxHgmZynd8X67
xOeaf2yr2iiyRhJHzWx2Laj8dPFaRAB2thW0ptMBl04HhtbEcmzAd0XvTMcET8vNHWwPcvCCcbJd
8mBL5LAlWdnYzXZdQKCG6iuYXPxiYyOkEGQxlJekxvp1qRvt2Bpcsbl4ohSgBY5PA0OvfYNM61C8
TKU0Lpjz/fAC71vBBuSJjOJ4RXyC2Fma/A2m9cCNYKucpk0aO2c0rXrp/97vuFdubasaVlghVw+C
KYyzy06rGPfVaDEET4daArBmXrlUMzBPzkrIezOlgCI52MdRYQT5HaN3ohgn2Wdb/9uUBG9MCl53
BnGmt2jLRDK7HYnHc1NHRa7Zd98rEuY9Bo3B1+VIvisHAC4e+uYDeazbiTmH7VQ0rN+3vsMPosuV
F0l27UceApZiskr0z/1Ei5OKInhbtiNtPCWl2/hmdLsgnaPaEVyDDrBQGP1qMq6X/MryD9vxNmZr
POUmZ6EzFbGnFK7lkfznDxTeStvdf38mpjp3Cd1WjxPmJpRT3v6rdVgq0K73IHOnVl05yxSAmE+B
YRxYKi3IV+uIHjqkud7NZVSporCTiYqnblZxBmg+mHnCs5fW6vwEZqLmsI2RhiitSPDjxSwejrba
UHTJsma/YS6j9cAGQjH1WyXDeHzqsQTaEDcaaShZItLYnXb3+A0nwmjeGY5kapu43ne99MgtEYhm
HYOQox8ryVuAZFS0oYXO4xTItUCAD1CfIln+EPtJqo/KhKp4e8wiKueZPegnhoahM7T/iK/t5UpZ
x1H/Izt8gJ0ADPCidshDEWklc+0ss+S3xJ1n7S8BKgqLJxC1mjkjn+KFa3UK8ylZLiVkY383f+nl
0USNFzdC/+r4JDs831aK6HA6Im7QmJyAic0CTk0qcbuMhcTbHFRVgb2LD0Dw5aMTYE4xbcLxIQtr
9My7XXLEXnH10RNHvdusax0gBzaq+iaTD6do/76MPMqV0Hs0EulhrhDnuV9hx/WSc+lEjgR4300E
HuHZpWsDamGSz4wOaip0NELsqfZ6MjbpEGluyfMLnPre9mpGv9g3XVskPBTzRGJyeUlpzq9/HsNY
b+RMV84jiCz8S6Gyi4dH+nch+BcOrs1YT5WBZ992rXcCjd99wk06esCYLWVT5F+o2Pk5pBfIzLzQ
A0KNNcE0f81AIm0e0HZLccaDZ5yvKdsQFkB8Jo7VMlzr+9rbNbnfNM8NhR4onqIRgJ2uKjmNzWq2
wZiOBisdoEyO3Er2bGYm2JbFBTyEMX5/jBJLLpDTmEdM2h7YI7kb1ZccyDovOIsOVzvSr6ehvUex
JA/DrFhBXnpSkKa/WZLHSFGg8Tx2856HZQAVKycHYn9sz4wdMor3y/Qrc7MwvKQgGVpPlvweykVr
kYJVAo8ttDoMxreNituJkLcm2M3o6VOoRUGT9NkBGE/lJchw5u7YU3d5hiouXvb4MKD3r9D6U95k
yb9roVLJEmwoBfqSLEv2q4PQ73nQqWyvzhoL4AmzH7z3e9BTQKEx8WxLY0z3pf1rE2nAbgapnQoU
DqGS3S25skdjeUuAg92nkeWf+ZN28HdocGT9iucBFXQGsJpVZiZTZ6L/YMS06nNX2bt7hhBaYMcp
NseWpOzi/vZhP32boG178+PDRCytYVIBMfx25DiwYVlATua+1Xv4jhxGbkLu+xjtnaiM1YpzZHIj
Yo2sUaZEGc5AEeLBDpRMzSqjbkqKOlCGO6BhHWBxeM/hEt5F9mIURudpLP0VeULrFdjEuSuF75q9
k4gF4/LvIZbrxcqRF7qIDgbSg2fhLQcLWdiNbM9eANaGzzWf8srcLW4RaXu1bb1zMKOK4IjkONi/
IxCZ91aHFNY0BbfLuuVfCaZ3qKp2OcKitBqv0V5NklNktWTtyyjZKn2BG/UCCMaZu9vaWcgE01m6
80476vqkn8BficcZ6yW7T2UeZaz79QGhAgQmffZYI5wiotRL7nwpurTARl355emtbrgrjTsAAwfh
f551ufdd7NNipurgYUiE0IAYy3URQUnWJiZfg8qSWMlUk72UpCkGtOVX0DmDxjDKW6c0jZY0IRR+
CNU3+P9LjKDEE17oKz1oUAbdX5SExtLFqHvLDm7/wmMQlmFw0rrXxkAbChzVj5NsrHXzHn5eTAa7
qPdDpRtWcPYuBUUnFf7+nh+X7lGfhmiZX3nHnwDuVCuFHt6++c6bt8UcbB480NpqfJCjTPmmQrTM
X0OK+PXTliIF3Cm7tAdQCes6JczuPGVRL74wtpwtWmAuOyHMeSDZZkLLJFTzuacxZ4HQ8Phd+FvK
QnQD5xqM4j3d8+c0iTnn3ZF5O+vBncLpiir5+EUMDCIVHMPw+Xxo7869loj7yOe3GEeiV6kRg6Ad
hCHOU/jO0QnYJl2V5fxcSsDL2/IxsW3SlJdc0Dz1B6BXAH+PeIx/A4tUawXM8tjbCjljELQnrMMl
XNnL27HJiY46bzsVsNa44843/tE9WF/REr3npwDQ9Lq6jdxiqwqJMK74zfPHnFxXORQSJZg9FcXC
g2vj5kS+1CgUyPwbE4iQ7JtbYYHpm1ipkz9XNEe113jlSkI9lb7C2ZOGeW2Le6NkmYUmvWprbgzx
vinOojvjQnZgyV3gjMfSTFJzAwAgIDPeP0+WWDqIQHt0jmzUGlWp6Arj491zdsPOM1L86T75xAcc
RN8DbQ3Tqvn4+QobR0Fz77UkM5uttWlr7BakQga0XWUOCoKnUbqZBiEU98+JnyEH+fnuGwVPcuhf
ZhLDM8TESGAKWfaActN1UCbYyykWEJQ5ytMK79BgIIM/sFflphFjlL4J6QxjrdNlXYJzTbUL/x7q
qSKzypIqf0p1bEI49mKBwFb9nX/pC6Krvy5Nu4BChw6RDWNeF8PaMp5agBxAvEl5ls8Rn/WFqYYr
7kq5oMpzzYcSVc+UucbBMDjtj9d1aOGUQHWh1JHATWh810qeVZIN2bb8vAexlt0M4UiXdofHN21H
pBkK/kdRu4miCXiU8aan0U1jm901K8Ja6G+5zktUIYBTlK2tgVnBHd0W3Ba7rX+1m6eoxLJBnYTf
HmOMR5T7xET1Yf7jiGr+ix8uuFNcLVjLjLIYz/fESRd2fGVlhjeY35fRz7KUaj/cqrTu4SUQP6go
ivJ+Qk4pWYggxrB33onbucsi3xBGdm90Z4FSZ88oiXgQ5W50NOnoUjkuD70k2cE0gkAuncrXclUA
XRvR9x6XtW9ykZcrepTlVKgS/+/pLKOAIIKiw/8ROUfA1Dc6hng/vmsxuLevYUFTSlbsb2n/JMfb
2i9BoF2RJ5wE5O+lHtM0IS8w5y3SgauORgW8PWv2DOh9CtaEvPkG3aNhHJropVJMR2DEkJsbtN7d
TyWHfNZue2GOcYyhGRMyQ3fB+D5lvstCGXoFeX5yWfGxdUrWZO/ZeJwbL72Z18jtZHd8FEaxOrzl
V+R9iV38UVCQoby4mvePRHn+wIwh2+UTwbXRsKQyKTcuATWWA/C810i/miSQuwlNS3YFW9QOU2M+
zvMx1DldN7TafwG4MJJBTbQK0kxzkDjyeFjZWYF0tNFCA518VQwzhWVgccAyTxvyZGjMEXBvcQLm
2A+Heh1pteIYqnhUDOBCG3ZWt/FmT0dCUmbzhmbObaoI4SSIjvfBMCrMO7p4nqH7E9XZ5WQX4JlO
4xCo53GZtxkf678xMCSwR7jVRKxChXyjJKfzxmPXJ3fdna6t1dynOA7wDUEu2kAiCP2SwiI1OKKR
JVfZkpgkxkBCFqvG836VW3SwpP9No30RS73KxDExi1wTsoyQ8Bd4REcC+IEBYuPoQtzD/3ICREBA
NCyyC6eMIyLJoTObdX9BXcZhTaL83kw8omd/+FCCBcczhGxtU2yGAfTseFH3ExbH9yNX9Sm622Ek
O3qLdpU0vO/SLZOJoo5zZcDqQSAAJLlUPA0W0Lku7DUhy5I4DUNc+YixlUVfYPmB7AXpizbDmKRd
p3ezgoikvc5ky+tfZwkD11yZId7JDB3B3TVss+U3qNWKj+DTHpclGLdjE6nl9o3eR0e2mHvIHG9D
6fMo3MOj6rAMEvOT2ysALM/iHIhVhoS0LbCWV1F8UipsGZMH02gcIIjyL6pKTLsmoto4o5QcXGlA
3/hhW4X4ivmMnhIp4DBGRovFfeR7JW3pKlsQm0dck1r6sK1pB9FvzD3ihUHQ46eZgN3h6fQNKkrO
ghYpQYxupog0a2t2m0N8tcNDEQKjR0x1Uz9quOQq8o//0OlAvTPFudPNsBTLO07FBpoImFHCUlu2
ACsM5EgGykUmunmAVHZVssuOcZMlPpH1anJKov0QPh9DP+S34pb0/63G3lZmViPMcJ6QJlG+awmT
SibhLVRat1YD2czar0fpiOfptgs3K870oHzEgA3Erv1XpQRlM3LUR3A5+jTH5w464Ke3pfNYvnV/
d6e5zJa8RBqdMLFgwWGaYVQ1TYHrc4W4rjigQ2tJJmnCM+Lut/x2rWXtTtpn20X0x+qU7m2A/BXi
3e7ahSVbo7VzlolZQuqtN6Rif2e5HWsKmgG2MuAp3vkCyIqbo9T6PM52OGEeo5keS/eVpHj0AvnR
n1RuKK8xCXrKskKKTfFanr5g/S64VcbBukqF0Vcb0k3TejS61T2f87N28hHbnkKVYT3XjcIhGaOG
o/rM7+UHj3dyJO61z4EwGbfUJkvMRMfU5u6s/jrSBL87B3OyLXfQBhJOX9EVZ+U0fLi/gmOMTnFd
5MMgYndqR1F7632zAoOwYxPLGaa/CFyTeEojKDLAEfwx+vHma1XLECU1E4B/ZbK5ugF1klQohLL7
QcwGpvN18li+P30RKPXZ+0MF3ijMpHYh/VPEKvGS42+FUT46TGzBFPgJXAMkrHwUTGtHjwQncN2D
D+NNEuE6JjQA6mU2FfH7ETjw4VWdUH3uGco+dgu7GmCtIsEB9WrRbzyHqgVDlX4cUKQTrL0mQe12
uBp+kK9sSKpdizM62GTVqSAx2EYKVWrdVOSNkrMRirksFSPGMB0zmSD9RenqaSXXw0kp2ycEgW8D
1v4Njk0OCfmBz8KGLJMBk3s7SDI58GfWa6XENndsCnnTkFFaJYdW9LN1UwFLH+JtWfBci4dmyKzb
C+dZLWlEWdr0AIDqwiW1jOEXCRDxrOjmXIe7xGpS34MIxBm7MR5qjyCtGzzv2ue8qbmiWFK2SCnQ
1WR/9+58EyXH5/vVtNhWnyWVhCsACFfsdiQoBTmMSvb5rgthagoqCZqdvPinmA942geUSCS80pYR
xFz8JvjnbZs5Uyy42vT01Pa3ENtkYoe0WSep+7fDcMUMgXzlJohYHN4Swhj4dcM2hXv+u9ag/513
bGvJ4q5TrA0SPy4sPhxsHENAe8ri7/Jqh/C2vDLvBDclqM7XvKVO8WFKaavuafS/kyxkNj6rviHL
97dNPAn12DmFeXk6f+u7xMQ0nnQZV4uzBvK/NYEhLG0ntG4zqmnV7ZVAOT7Jfm4ytBGGVeZx+hWM
RcmN9el41i/mD5QDTmTCqOiXFxsKy1AnfGqSO4YPkjkOXGLeXK7A+wCKEe2Gri/7dJin3MaP5EoA
n1Brznysx02HCqOxVhjOuk/IxHQ2LOXFOcLUAZ3PcqUJuTKGvYyge89euiR0edPRkP9rMuqDHcSx
Xam5vmcrgEc8si4Hiaevz2L048wt2kz2T422ShuvEoz/XdY1bcmBr07S9o5oEw0wKaSrtpBC58uJ
nhSUEa0Hofs/X9uHaVHtkaCopF0clpMCEZQpj33lQ8KyQwXNSOTfnwrQ1bRUp9U26/SRRtmRV2zu
6UH28ud1FLHlRmQkbrYxg01mpMTHzGmFxSpdJpzJXuUsOdyrxVLMLZ4PYyOD7PMiwfeYn+E076No
xbZ/Wbswu98aVsyh+UOioeV0IKUW6L++rBJwJm1kQAUayTuJ0hANKmxm/BwjiX1s3ecBi+OO4Lup
RyAmLu3lEBW6h9q1USgqvI5J28fjUGPY0R81Ie/ENjH0KwBWV62wUVU0w9DKOyZC5x7yW8kPlRBb
11KlUSJBPMg4eGg4teAxUy+xVFsYwc8tjiTxTt+hIGixlO+dS7aFD0N3RfZ6XiM12mgNswGoKCY2
Bq8vpowQeYU7sCIabibAROEuePQi45wAmiaGo8SYD+f0zzNf492Aj67mVkGM9sm/m7YCUZK0xJfd
ODGHLCYk2Mz3AnuaMfjv6x7LVBRWryUX5FzW0zPs4oJ5L9oOzDeUVOn6fjU9SArULIeKLJypuh3z
6Cgy/j+TUf0f+PUqvoW7vLC5Z/SJQw6lo/R5a4XFojsOxWWs89bviqD7zYogCIHAL3Ec/7MbWB5c
t5mh6Vq4/zTsslZI4ANn/bQHBVdlRCxBag2O5wTIu405ffjVNo3SOkDEoiRRYg1Lc0LDAr1c42WK
Tj1PxOY+1LTwiShbksrtXC6hedkmWEg0uzeidCzyeRZMgNSJ5ePKqXeoFUjKUjE0Rjw/4gnff447
cuhklfLMYJZQXvNT2kXdeEMRxYKlUXI82za53hjvmVlFCXCjHr//Uq7lvw8ny4vX/C932P/TBYUm
/SdPixTJderXNxJf2RyTrju7P7NLwFzb8pTWLPcB4zpHKXcN2rHzESIyuH/ubzS4a/EMGvVi/Ind
W5m4mgVICK7Iss1oJDzs4K/F7j7MiR/VWUiPyfZA8YHTUD6AQm7CMfbAEhtqfW8xI3g6N7VWBFoY
xi94XTX4h6sRYlO2KJuCBBVfM8t63QZDavhpfKPHpoHw6qLX2p/LBFEEUe2YQdh/Y2KE8jL1mP/s
6sCXI84kb77YlevVI158yymxxdN6iRdpK5NII1TrxL5uyQy2Sf53dONoBVRX8TNMyxkm1YCq+Rw8
SkrVVVDrsZPsYAWkknqhvm7Q5otmJDeEUgUbsdJ21ucF6LI0UAYVtO1U7czCGsXzwxRxiBTUi2ue
IXrIAVOf98YFun2Q80xew4ABskn2dYBy9ytWlvy66XbOREZBu06ROXeoo2I/JpAHFzNz+uSRDNml
r7nTYX7MQVUDIlWqEVPkmDtlARJdgDo7je0JoJ765VwEk/VE0vaL/XZQ3O8B5lFYTpOHux2wNOuS
3M0N2fu0pGkWRMUsRVZZmBOo3PspXJhJ65sg7GeLIaLEZHe8bDg/f6Ww4hCRIF0g9z0UJ+YdaWi4
lu8kE4PYoUMkz9xVk73wh/loPhg02s5vRobgv67XcoYlpaZH0r4enTOHEovZ9afGywZTuTYErE5c
DqD1CGZxQ3txRgA7QK+OAUAUXoe3+t8bPeZpZ47SjdNPo64kS0K0uUZXfduOlKlLx1TAGvk0q0BH
RIg05247r5WMVwMO0jKsCRJ9H0inqwdcx4U/eRGPjNUoDI1qZJI2tIGaWmnWxCbfKxLw+NPR7EoB
Z/mxh6lsbEo3iTL2eah4JH+ZmY8PCz0KjEt1rtKS7mJTpx8Lo0vnvwcXCNA9VZJY9DqmBjRZewZh
Ms/enoGlfuxA1jUuQL6av5r1UjrzxHchWWacZlFrRV/Wk7O8ERxTVUQvNttroFAhZDjMUblltbDs
k1pbOquoWSXfP2e4YvxjvLlFKkAJhQpP2nxpxi0N6vUzS8n4W8+ZZ6kRIsieFWT+Fvu/q4CxyfG/
8vKJXgQOdIJ/3Pnu+12+vk5iQAZXmP1RUT+IgsudTpVeTn5DBHOe2bHvhkp/hepiujuugU6YzwXF
Z12s1ckBcNR2Cu+MXeTvAn+GwhTxz2qR2EqBRnrInWounGUGQH6V+jkpz+fEESwu4pPnmTDJ3RQl
ZuC1m8kALv7zcb3toeGEGLzN9CrAGjiecV2CWWRefQT9NFLB9MLnvwcq82H5p3/lHY/yrD2/ejUP
1YPrX/GbBJVxWebhja2VuM1tHEd5pQu8NnQt5EMKCAC3lBsIA60iWpdsK0YNlbKlnRfre1LwCW3D
TULM1hDZ98rdlgwpn+hK0TexEHsFhGqEyi6sUhx1mpF3p0Ss7eKJjSc8s0wCIUVo+a/ztVBAK4XP
mu93uPDAVrvQA7L4+DSMylh9fq3LDNJ7GE3eP0nMBKXslEV3YHJEezI7jSAv3q2A74gDqo/JTaXM
1LMONe77Tkc2YoK/c2s85yX+EWxuCrlH/jc9cpw8Vua3dLHdCqHeTWCMyoy77aWmg1eGZyq+QDvt
IzLImDaq1XwzxpsCI6QEqD/IVad5NAA2ZeqowTMoGcWBGPstY4VUbRwvW5Jukg57Y/CW0xiKKN7n
ZLiRU8DUEqyoRMtL2g6vAAcVoS2Mloy3vSs+yf4CjIOpFe2LSiUkToNxfe6WDQjvt9e7bjkEZq9C
uXJ7nPOfi0w/Vd0y/W7zH8BjF74jIrdwMeEq/3grTWNyAFdsqD7PGiLm7+NP/ZdBb2AO7OxS66GX
wMbMp8YiY0zy27KmPPLeFBV+sB2sgykIsReFnujwG7X4DuKlg1fCKMnEB+vRx/r3Mmq9r/uNbXhX
T5l4zcpt7eeKA9A/hKJvND/GqIDDuR+NhQ7CDXQLZoTsTnXdAkO5nH0v3xI4qO2PNgxqqqba+u1z
EYT3RjJN13fSLqP7iC8TPkV7y8lNkEuQ654tl7VkVM8KVX2u6Yiyq4eS7o9puFM1+DnNZaFXNOae
saO/RpQ8BlNrOWjDhheS3BkUEc8HYmCvW7S0KZhfcsZO35OryDn9YLhze11VtpfFW5cuViasKPbX
g4jo0w7SQDTZXcruroWbDyiSHLs0GMOU284UtN//yUfzBMc7ERiDW5kYXpQBtP6WVhvrhC2NdIun
+W7FKcc2Q0/s1ctvJO2+5rJy4PGYwEyHlQRSP/8vPPvy2ZddgSCmNkEGIAHBFFdTc8ofo1HNGYuK
MI2RK/Z2S0pVrt+mCm3d9AFNzJ/HNrayN1hEaAeRJBQbJpUKnNjDf4lyUkTvo5psX+hzJCUFhIb7
bhNNicloBrM0eqjKm7CvmUWtfNWewC7XI/ljPUEAqQcYWifZDyhvq8CEJD4GxAmvPEJpugXMLzr8
1/JgYPXsIZJIvSYgKK/kX9VJOofxj2cNwMH6o6nS5YvI/uZeDkxnugmsq4ng5t/gxktyAsYs9HNE
etndiHHDq0ldGzcXaMkR94JsTobaPNW2FjtXGrMMJmvLnLEcbw1NdLDx28IqKUVZQEazK9m9oQ33
I9cVG9VaWniqtvtOJvhsUUqehHyW9S9yQbTM7Hshj4VdkVvSBqNl3b9qmNwGWbBXgmP1FTpgTDxc
ayP0ksAWrbu3jfPh9qBXKsDl3Jp9jcpEF3/ROCsn1GxLu3+vgzUALQSJbBBv+j5ui2n0Z8rDjIIC
R2DkpfCvtgtoLaAH9ULH+RN6EdCY3lT5LKbry7RKfw55Y2otc2KtTBd0mH2GxotL44CJ3Dxxtx0s
Yef8f1y+aoLwU71orHsLUVTO7Su7HIhihStycRdeujsxRTK/n/uEhJq8G4Z427XC4lTXqGUxABxF
iTNX9WGofZDHpEmzp2yi89Zn6V/U+r9WE1GsR+BtqclWvBZ1tHSXwCQbqRIWXFzrQJaW+IqrG4Fj
Deip6qL4zRfv7Qf3MdVUTRFGj36ENWVunbaNuusvmqB6z9dJgpsO9SQDmVZY8GzP8wrUVl+ajMs4
le1EmtrVJH+Q+oX6stBrNsRRwe3DahE+p0AV1xeFgZanNaoKho7X0TciqH5zesMpxbAkNLBWoBhM
h8lD49SsYhZ5z5TUU6gSXjlJkAeux8eqz+hRTR4E+40mtNNfpP+5LLsvYSL6SVXZGwpP8q7bnHuE
hnb7PccKVLqOxNiSl+BroT/kJbi3+Wq39iTAvgzc8LHonVYjHunXVIGTwJufBc1Bpc5mSrrcM1W+
5K++GMwHJkbYZFl7VIXuMud+SbtZ5dzG4LhO9H7snz6Yqie+YFI6tnOq2APSuwqKqrnyZD4fmQ1V
/xLx9VT+g028GSWrLAgo7I8ivsGsMcptlz/jDsOUats7XVjJMSy1dqmOJgBwxRxx+t5E5gsRQu/M
DQ/6z496ANTo3x/HJ4Y45VlzLnhc6EfmjNBys/gJyt+AjYQL7voUGg/+M75lkevW+LNBTb7CJXvK
eZhFO9LO5gC6wBYo+8dDabbnBYwpfXtzFIEdRw/oPLy7svA8x3jod5v++HBMdCVKqlavuttPUVmf
J4USoHvfV5s0OfLouMBIG5GQrteCHR47Rb7wXdbiqmaaDXTOCCECui/8N3LByuMYk6GKorjCVCjp
Ce4MpYjeMUdKlB6I71wUps1oi9Ofs1unORINlVkH8+ZD7PO4F95uO5PFKErHDOAC+dQsLIxnG5lz
9mdXpAmseFZ9KfgRrBVHiSrbW+kCuquNhTYXjvrsZKBjYOKcWhm8f3NOJk2dFPPQpTHDykyPVfyq
RAK3etFmzIA28ljaXYqbpLxHdkGfnwx4X2f+y42l0EdmC90TnWqpIMFt5q7vPPv8dKJrH8KQ4eN+
lviPARfTqNEy+tM1upk/BhFLzs5UYNU6r3GHeQskkiJECzytA2GJ2vkWogmMF/wt/DwZeX4t73HY
bEfGri9V799Eta7qbgd3H8q6NXO4j/6Qdm/woW/UsSN4dOu2y6XFIdyPlfvO9ybGBmH9GgburJb8
0SbqAltDjHdS0ttdj6RF0HuXDMAEaz8N+t/HB0aCrA4TTzWTl4Lr2ipp2aC9zYbWIDzL8GY//QHY
q3IOghUMtGCBKxhf1oq+brRbSziL284VitDHDztWzdmS8BU0qF60KtG74f2uIegtHHcLk3Z59IHG
GhtYlBdKMKO7xg340foyaXqfIeNB4lybfO6tq4TA2qz/0NtGaB+4Mx/4tJuPUvAb60ORPnPdRDje
HDL76Usbd1s/HCg2jDXFIFI0f8bnWgDLee0ahobwWn+2L+lrmqLCyJrOx/Sl7RK5UEj4KYpss/CO
X4evr1wAEU0PHR7s2odW2LQrN/FAXWS1GD3dymNac0yXlyqUEqMLxlnQRHyd4juzBnUHjFxgnJG3
KcCgiygHSi4vcPrF8XcX5aLh6T3IXs40X0FOZF77/4gfJxoDQB4QTSUi3Lv7pcjvagJlKlsZA/h9
bYX4RRVJHiWc/bsK3PBdYXY6yAwe8Xz2DGcp/xNf2v3XlbXkVnfGJYv+uFnP8kyARJ91iUFt6loa
Xrs81sA9CFpVAdedEcb9/BGxkQC0YNoAhiRguxSPjBRzkprm0qgspeIoz9h7xwXOi0YSMkOO5pKG
WCU9Y3ylbTCv3gtVk/mHQOerWQwaAqsvGdMXTZZtTyLxooagiBrxSpxC9+nZJyttpMJYt3PyRKxR
bNXT61gRv0xAdRhs9SG6E5rf30u1o26cXDSj2gExrxVzAG+9zByk7NAGHg1tBF4DFbBHhxQ0SisN
jejylSZd1qi2ilfO8w6VhmBusrFo9Q/yzvSBzhvCwplhWImWNeYFESWFcf4kVGvcld4ZEsG4jTYo
TlEjR/VLEkAwWXg3WIwJI2DhhFlME14+vI0qlHFqM5zK2XE/wc2YeE9xB93IVdvWww1N17syxQeQ
ekAX6l58Dgw40AT2FFJ3vouhp0rg/UiaUAwQ8njdIQ9FnqVRNVw8LFz3u2Fvr0byNOiCYT7Qc5w+
HxyjvsWoHDJ15aEdgm80ZUmMwPI25b3aAmgVKUhfBeWlcpbWIfJbMreuF1jFjmxUL4zs3htWR9QW
7DqxF2yKeAiVti2104d80pGHTQC87NjdrsDhjwrbFQhNei02DGp22ZIPP0uu/p56FCZP+FqXlQK7
u0r9rOmthkvFc2iRgIOgg2l/4rK0yKanz0IC66uHdfrRwEytRJZemVx9qMFRbhJIeE2gi0MTY/HT
JBqy1suj19zFKgxuBmjjdQhLSVWVf2Zvi6Ndqp5G/V0y0TJG40tmJpswm9YDxSEz8CFIfZVtcpWx
Yo1mfDw4D3G1MwgyXQNidXXKonC/qZUmo/cFpxIBiHpWS6ky8KXt1+Lvgfya/l9ztb9nWh9eEjep
nH9RkpX3pTRz7q/KlyBqxttyMiDDTWmHD4OEvIbwYF5ER6Rv5xjn7zRd4d6nYeo7zErcONm55VNN
4Cj+NDutCvHd4dW7eK9HFpgQT4QYNmKI0R1z6gN6N+MIY0VoA8Yzyu3TdGk0ER8bX86FeVwHL2AV
xoUxm8I0hPmLNHhdn6wwJHVUam903FnTNgXfzjqn9buijqXKjrGlzIFbwWr0nPMdbZxplWkfjKn8
aQZWnBYH6nPLzyspE+WIFzVsmoRuPWgd0kgXRiHmXoByBcoZGyoP/8eL6TrQiHk8H4hJF06pjK7d
jNwr+iWNOSSLa25TUBFVDCeVKsjeQAOQbS2g7NQCHnu7clWXe64obacigh1rpo05cJ3zFWz5PthW
PMngsYBJWii7GjuaF0qhDXnKdNtJgi88CvFqIBIiQnvVM0VsY1MA9Qb/R6X14c/zINEOoYFJrhGI
J4Boa+OA1znw9HlhSawPqrpzy7VEuYWvdHs4H+1SAsQ0CuQVRPwpgy9mqEoJut6WeQbUXVuF7bIF
IxuIlMIvP57mcdblz7n8R6S4TU8SwXfbQ5uvjIwaQkSwOugh/UF6LToNuVqi+mzsMycjJFgdU5wD
6y0HNUyiqk1Oeh+6paHQZerwJLDw7CdJzev3pagP6BKzICCkysmf0KPdoWtzK0ZsOw2Z+RApEvWj
D3HYaikYmmSglP7UJnJRrXzUoWrrE7095y7QzMK5eKM46i+LDLAhWBrmurPvuwAA8J74tkQOe+Ii
D1Xt+fuMqamJHN09oCLbPIrU8BIkNofLbbD6KMeKTB5l5q+RyPH82wd9wM93molwbrMJqiYYe1N2
haVQSYT1AeYD5nBeRVY1Kk6Krhm+KJAncaLhdbAifJubSc9kn+0FfBnVZlYb94pgxQ2ahutCMunj
l/p6D5RK1j2R3hLbliSXbM9lvoyouNdhGKhyNX5ZURllqeO7ySO6HSRnhb9XqsnxcXJfR/WdKJ4C
6WkASjm3MeAm2crgADp1R3UdgnaH7gKwILhA3kOKIn8zsNIhHNaRtCPK/vELrBgEAA/VhwqmzDe7
hFN4G7LakYtDEg14t8SnAYwJaGC9X3yJXIEFEYRkJ9zY15hsx/AItcrFXPbf/Dk6Wej4k7bgBkSP
kr22tA7/x5yh54ysh/cXIgR8KKjpnhigveJpcwEuQsXrTAOFGfzpqGrr45RdsnBLxaa9wmcCs+Q8
u6hCZ97iUImGdv1lItgV+iFqcNl5cDLfzhOBgshccM/so/rgzx4cD7OqEv/WWdvZdeUQnTXqnGjo
OcrhF2Bnm6nC9kZ79MN4O2w4HFmqfDzCg4PVmMQmzDeCoAt8lNxupefA5vb8vA0DyschsormYs0y
ycmDbgON8K7JIUclixfl0KMnJ+Sr9BXum1GwHJ1BdlFN8TRjr/80y6iFuO3V7l0kCErZbnWDIQnF
2WgWipoXmNylF7EML5svNpEOKr76HRKbQmVyyI0Wj0D6gQmJ+BYxmjjTZ59PCHsVeVsQVvHm+xVO
96EmTcLRoFitnp15TcjNiLtJicNwWvcp1ZVZvcGOt26N91gPSC/uGGZWILaGzK3RzmXdKhx5t9x3
msMDhz2zse9VhXkY0NQ/x9Crw+/vuBa/ry5/0u+w3y9kIQW/GC2Iaes5SScJdgLIh5vjc2DCD5u/
Pcj2Yl31MTVnA4zKtFyHRS3mCuLitTjPOwEyWQRm2wKAh0cTonO0Sy6gMetoVcI74ZPMOV7E1Slo
IgUU6EISxVvqDS+9JRzl8gF+lV7JVAGCK/kOdSf4XYlhHwstzATuTLCvxqZjmGqWOgM3U7N/yNHg
2PSu6yqnHk7AaTgRo5Wc/2/Izky1AuiG0S7FVrfJUDf/eZePW4YDgnB69I9L5bXtOuCOvrSKjvFd
eUkbWuoy6sNmiT/cVPqSzW46mJ4FLFYOGpo7xvKDEdTdzFryKnrBLe6NFUzkou+V9RKGevZCckJm
eXZiI7c1h+IsSixbymzDn22NrE7Q9XuoRTgnaVEQavBFcAM4gk3xps0q2tRSsKclHN6kZseIusVB
DbimIJFl4N+zjryc47D0IbGbb7klvCKKb/UWw6b3slh8Y90omUxx86haUBjGyEBiZOACymn2GnlO
n7cRFxwikli7gW2OApAygb4LdO0zLEtVQrlKsHUPi83R9pWMeslwh/1dXeUfFoc7AG3ANbD2xSvj
veVMZNqI72eaE63oWF4+5pRBI5Zm+LgmzqIsV10NsTPW8jk0u0lgNqYLj+KQJjaQZtNCktNctHyU
T8WMKcV3+etqD97CAur6C02dCXZXm5yflYbwCX1fGw1VBYiSxDG4TfllEvQrIcaBV0NjZfMNVmwl
nvTM0NrIm1W7KgDDef47rZR98w2HizY9eSiuXd6rtkM94O8SNO9uksUjMHvz9qmNZg5zmHC56X8N
Aelv72+LhUohrTq2iVGPJwv8vPhit12XtFh5n7rSmmSBlANdyOiU0JfUF0d7YjcGeGNgT1j65vui
Sv4MIHTicBFCKkU/NONENdZNEjAHJ8IlCno97PDW9/45Pr1wuT/1AFg/2+/DJk57ZYJpg5uYVK08
oAexMmg+Z8XKSouZHUovFydLS3EkzuHW/eU5eEtzm5QFenD2dSxfSsDcpIqOTIGYsmZ29WmeQRx6
2A4oThMgH0gI1zoRXRrW7E2HBTzacn321QELYJLFHlWPOBJClZjYsNlDnD9G9YRQSY3P65NTXsu1
hScvNsrEo0v8bu42W5ywykPxvVGoHQZXz06XfPEhSwTDssd12fuS6PRJO49W7g7l8g9u2gN/nQ4G
Ya2cznVxABjxKODZ9u/dG5RAZspIh3uGqmhmKelxMich5BJZyKtokDgcT0JKYXx4uSgWzgAYj6y0
5n+bem0bGCw26wDjavXTnuK5/L4Epx90STl7QCfzGJxaU/ObVhEPEHEJz4X1hPHeX0jSpe2WJQA8
ZC09+ih0YtI9kQp/Twk8Czk3SefnWHaDHBiQjKgABYz9i0AJM8/BIqV0QGD5OUgs3XY2J4BjrR+0
Kv5LOXDpKKR2g1OwIKNMP7JJ69PXcBzIlIMzdrbDe5RAZbY6exs5fSs7EJvG3xVN3CQjLtpVORdb
2T7dCfPpNlfrf0yjApBy16PFnIlx3d3lyTvfcesiHkWTlJnI1oglHlJdhyQt6byyP3TY3r55SPRO
qJ8fje90L0nKs/6J3nFioZwLSIfebRPKTPjgPk0egG9Uvvqa16q/y4RDSpoC9gAKknLNjPoi/YgZ
/Xy4x5gUFW9M6YDxmMeqyvrDy9/HIw3ASY0xSwC3VaBO6hYDUr59soh9r1efWDixKU6amUjMgV2R
jHDXKM4xz634zE6XNxoyyFfZmRHygAsVbYsMPBqXFnSyT4ejBhv/jgaghOTyLr7qHrMzAZxm8Lm+
TuqPwd/mDsHxk/K3nKxl1EyJrcwxdEsmHMPcwbHjP11+Xy/BTbwsO0x1xBwmsG7ClTMdFNmnjF9U
cCoCD167eDWkRH3XVir+pisOzZLMX4nFQLnCe0uQU2mKZC8X0k/Pp9aB1hpH6Dz5opmFP3vJI7rL
vfjuHnSV15sCA4vhJtcK2hQpzzdfvrhx6g7NCVnxNIr8DWRdvPf5JLfkQTWS5AJpuHqph6qWgOXz
bDkXy5fnj74cM/HewVZ5uDWQQqJK+HL+mgu07KigMVvRC5YsXTs0TwMSpM5LF/ekmnACt9un2S31
YbjKZYx8385YybPacBAYrEwM1F9WlLkie2UYOkRl4NpYYOAY6LsyXEYWb/0oCzE+D/55ZPJnmB6o
6J4mVyG4LzouPvqMXAUEYHxR1TERFJ0unTy0Mcgza3T4zd2EwAr49GpQab/QbYZTNa4Fjxpv6Qdn
lXf2y71xR5Y+NNRo+KdLAE0vwn3iDV6ijHVFah9Vhf+KO929Atdb6jhRkNfkzF6HspFntcfZDbWj
X91KPm7hmyCivOk0Nwhq/039sTBndJUmR3Sl8GDgv4qIdyjzIr+c7B//jBZO48+svHU06auw/Q6a
s2VNmVPt277BdySG/fMdNlfiX2g5devsSPmDwfayRoLFpZcSWnHYGyEIdAIA7JQka+wRuaC9bz7k
WtSJj/Xe05ryr0MnhDmJQ573kDJtjGC4lKcD4PtoLQcTuK4Cc968gItNsGUoqUUGrx1oyfYLX88n
82q1LHtDymOi0/bOpA/vYmPPAvc7VdsARYilktbtOGvPcfk/pWGgIB508Av0Uq6HI7QCNElBjkUG
+oPb/6qQx9gcV3jL1BnPmTNe7mwW8KgV8jp1QyjHcx3vWXb75ok0SBDmkr0sUM8PVRazk83E0ZH2
2Ilz1699tT60l/aoUXQbuPgj8IWR+OaQWq5iXG6lvTbtNNMmJrO/tcOzd6QeqeR/wf4zXGkOmavf
mVtH8PygjuMHQ9Kiw8k0C4TTZjkZzxXFKKGy3ADG44dauy1WCy0Zrn/z9vRV53zrLwxeEJPDb3ti
12Ys2rmVhje/jmsfiTOhDv0z2XT2ExdS3G+qF+efebkemoqu27JDhYuviKf4DFSqgETBNQ2c3Nha
xXQzVr3eFrm1p9frAf9ZIZlBvpotu9JuR7sJvIh3zSBFT5blgVMdY6aVGf7y2lRfWB8EPt7C812i
we3e6So5ssEzxdt/RJJ3b0Oi9NNskTzQOM0Gry8bK96eZ8FDHwD4xOuhd506poZf4JG5Pvo7r1uN
7UUtzDjDYlq+LF3sFCUIn+7HYBsko+oJclkoh5vj1p1WNOQB3KCv9y4B0zTsTxNoOs7Q3aCpnxSy
PtpvLsqTUDP7EkS10qUaPkWe72/3i36QXap/tNeU2vXjAhBfRuXGTgaMExyB/ML5Wd3Cgu3tE5rZ
L1nM5CIujZLaYuCnqpjmdloKcjAF0Qp2Vyox65SmmcIyQteOpLHP29HZwDeOYBe/03+j30Zz2Oiw
v9ipm3wKBEshjA/gUlFkbSXEqC7pjc2qrGbdvcpkb3siAIPP0gpXxFfW5cUUHeNYyQop1n0vtDDs
W5Opp64x0dNC0iai1vwi9sEkSWeJhegQaxmcbdGNGsynhB78PLQib9CSz8gSqHbmEqQ0F0Q38UxO
Hdafu1RsfR6FjiRDWdPvI9i3Nuis0P+kHx1zVqCpTw3Z1VjFF0z1VkRihebigEAu6xwdmSyan3Pz
EMinZ5N/cE+HAJC5IiHouVooxueiGVUWFH8iMqnaggasBntdH0a6H4xh82bcvlANV4pfkFzMMmUw
9wmZ+7eljIpaj8xYCHQWntgeigps0NWlgKX2hY6KOID9K2BgF9zNU6txpXsHDYQfXu8Om6IFGzP9
FcBTqqYMS6ie2uaeRXugyav9e2WPbPnJn0WvyV1SiIZf+qAYMGaDU6A5Ek0nB8Sk5zRCniCjXZwS
6j71ueFOOBkHMVekxG6A3t6m5j8zyScIszTkOPLsGbk7JeaX9DuIilW5LpeMmwZsaqU2YtX2w4fF
HRMKOjTm+ndfI44uudRm0W7bmSY8JrENi0E7tpSZ1sDy9iaLGk0ql7/IBOzub5C1CzEH/nDq9eJu
W4UE2OOv3yAVLDVJgXTYdfFPDCpH5mbaIgzz89Bk7w9lXQwALXaQ/RerMIWTbvy//DgZBMtAIXq4
OF1EsEJv4/TsuwGPnTk+YbDA3aZaRA1Z7O0KYs38gm4u1qss4PEu2ML/3KLQwBwuzy6SM+KEJfnH
G5EPgx50621flWIbQxBpY3cPek8cZNT2IqXcOtGeHW2Jgj0e0P9D+7UW+9WSIkvsBkTQoYlluZem
0m/hDHp9yYVeey2rswglPZ5LNfGuwcqH6RbR4LXwXJxy9iwQRMq2fLsHcO3i6HTft9NY8hnQKBBT
5jW6UftpBQOE6TSUfvSc8pEnR+w2nYn2Vpj8fjGlq3zvEM1fpMaKprlIFJPYzg+HVzzlUnMuAwv5
Rm/2WJEshumCV0nBnyssQ2KqBvtxm1rIzhpkbOELbMI1K32+57YFwKZ0aGxFzqnRPDTyopyAYKs8
a/pKHBzUHkrNZFihNN1WHMTVmazShlmKy+gwp0j5QzBpEZzwtDpGxZbpZHlFFU+q6s+aaL4utrOB
ZNVmjNQvs45r0jTNFoM0GZg4kEMH/5y3BZtCAfDyaujqnaq2EQ82N3qCEJZLixtFA5jLJadmVxRS
DQ4EqTElMwSQUDSdVHBYq5j2kodN7GE0lerBHjkJOsqlFd+MHtNH8B5f0SRUrkkFjx8SAWw40LAm
atV48w7PtywnEEXcTGFRWcmwlPXnNtAzkQmpLal8uy9bxaO4kCysVdohSapvA6FP7o+VJ6KFAarn
20gh4/QxgB28zkUMfiu+iNJWqkoLPHSAaUXzQBglTuUGpbvgcqspSMPLSEo+yvlUthj4apBlnnRn
l9TTLGHVDwode7VKuLW3Edf4XjTmL2Jem+wBxE2q8ye8xdfCzznM7c4bigika5988TCEHWM4zw9Q
ow/PU7NkcO2jakQfmOG/vqjweWVt3f/DygKOFtIEXtQ/PLaSQICxPj6C2Dm5+t3Ya4LLTxSp9ACW
n4LK7T3gPQtjmcKi8F0ktk7Y8TwHF2CwUnWGmbJAf1fhW0opqzvRv09HBU1W/VvNiAh1N5e9gDts
shH+TELjaxQ5V6xH9JWe12rj09OrPg4Sl+VqoS9cYU1ePENdgygmQiDlz85KSy7fKnLpvrHLkIx8
/KXDkZ9DlBWOV8/oT+dLqldDkgMNFtvnFUBX4a4NGXRFGo0Vnh8Xu92hIu+/IOp7LU2TpXJHIhPL
7M6OpzLzhzC5NHPmQQLWwsE7bB+60E4BSep8jDfFy45YL+OwZMM0D94Z+s6swp0MULy3HL58MjzU
xQODTkH/VAcG4U/egn7+m0xmvy80135euFw6pD7TzZdHKTCoSoA/jGF4Qzo9bB95urr82NlSCDwi
+tT0RmJPMtzcdOo9dEOFvPCaaCtZIUP6WoAKLvTLcDLmHe0PM9XGFzPqY0A94VI1FiELLCGzuoja
+ycpSNLL8JnrHOXvfaBJLVGisTUzlirUf3A9w2Qtm5IQoiHNV+1k+iunj8zEQYEo5Ke5x22fYzbj
se7p+lZPVmTaeHSlpcyfL4EEMoRjGLI0F2Daxq1GaT52ivuY199mmsVv/ZowUTcugZUmkK2rBPnn
fgEQ4u1rpfs5r934LMojNXXQxaYIFAs89p0oJn36mvpkvlKb+Lw58gbGpfwQ3U3NcIUx4ObEI41x
Gq3Q2GUXxdhFZf73hMtSOo6DqMBd0uK+flHjOJw59JIpPITURDzuxvbTfNwjUEo7S/bo4usSoBeX
Myu7RAmKMl5Q7ZXWxPPFoVcdScKdpgFc8414/2ucGieW1CzbsAyUFl6FE/bgCH4UFUXwcwVQCFDY
6EPn5OWf/EJmVDcK3vKn0dp+lVQps8CW+RCjVtFJ0jU9lsdDA5fabJLVhvcwgq5/EGzY8qYp2c3b
u5g6+VSz5fLb4dQyvuEtsc7I57yG+bk2A1OBSJ+GbmVCDC5d0eRTjABY/+ydXxzqz/xS8TQSwEO5
M56JtzRr3buoERimQxnQRGQ+8a98ZOsJuhgnNGG7WS5azMcpchudSCi96f6OQXHoxb8zLGSOWdkY
V1T2pbZzzd4UzppfuXHKYL/cAAaz5jv7oWHbY7CpFeaKmlAMuySpFO3xep4Ye1fFCijAgGgVUMcW
5rIg0l/nQvf6+humAuvWas1mk90KH8YYadV5BPkaREWOzV7PpXj2G6RuWAR9/Te3ZYF10WmKcv63
LDOuQzPt+yLRXzNG+gXJrc2j5UDAyk66hxkGpm4WzBQQD5beB6LdYWvTGNkSrKu9CpAJTlKBBCjH
uT5QRk5Ps72YQFkNr9Fegh2ZrRseNFAbxtqooEke0vRmR1JqKyp4vClhlpfpmmg0uaMGP2h4y4RX
8M8PEfOmdV0Lsx9GWvodC8d4UbZ4QpczwH5aZ1/lhJRQciKFHoyKIGjTnqjaE80nYHKVUb3UsLJ1
/qYf5PY2Hz4nIeVecTO0GE6ClQg3hsrCnQroya8nD104XwW3tj2lotKj5FE3+uBQcKHqwXr6srd9
7VkU1NmfKlRjYrXkeJU7NaQX9mqFWn5zN+554FvkSBPwbn7ysyw7dsHBCzWkhfD3L9Ck0pRpRfCk
sfFYiWeMar3DdFdcqa2gzgY307bYGuahMT+4x68Vbm2tjzA2/ExwzGu+8QPPpsj4vA4c5UGiWxl2
iohWI4qdFixa/BaQhyPz11lHq9VF/ni50E0YRPc0W0MeSQqGd8zCLVddLedg5JLRjx0EQ0OTQAJA
03ZtS9Mw6ihHCJkjDy4QWe7OqOsU60vV9BJ9vt8zMKTd4LcW/3CImuW9jkm26CV00RkGlJeXm/bx
LWWCjeetLSpXW5r641Z2lY6S0k8gY4UwLcnGrthPRefqeWooTdN4LAZRgSgFVg/+9vUtzZm0XVTT
cOPyMwZ+/o+HIvU1pw8IhVzw7PPNtwh2PNQnhCwaVdDe8wxwaSUOA5aWxZEX6iirjQI3HUNuoTKx
0QuP341C+qkWgzIyduk+1SOr4p7klja2TF1ir+ra1QaeD3JEoBB3tE1fw2Y8BoP2ZkFnFVuCshny
PG68rQE6sCHjV9Mfg+NF/3HFTIC7M5RCpW50lk9p4MCyXxbSvQmaoZdvlIzGrcQeEVvLbNA+J01c
UNiUgHOgwqI4048w4FBZQaIgWNEhCVqBlUmUiDGxTDPJMk3MI+bo+1EssQpTFxXhDm6qHcprz5nz
d8ZhHC8+uBC0BWmAZ5r7Tnl9wEp+c87uTspO2vrpxCyKbhOSKJJDoIYvdENWsuRuSNOu6ZlM3ccO
ipKcDeLSCVHdfnXKzLldtAUen0dUm++z4cQg81uvrVzOjOZvOfI0eY9GImllE9qz2kTc14n46Q/g
ril4h7gyMwOpbtkQiZQqCfnDszuPVyV5MY/al9aQ/vESMKw0QUi/lJt33SzQ8lpDOZ328/X/tEgZ
GZrGTi2Ke9VbhBHcFaoaOwmQ54OM4wBu6FlDGvtHsIf/gGtZSBQlS2mFdOZsZwylzFsgFVpaRT4z
pn61nTWZJ88AmhtF2hv/Oe99LMEYT+hw1M7N4FhF4Udpva6WAInmt6rvoakCRqZNd1KTGVcE98Af
qTmbHyouf8DNN7ix4pWirgdOHn3fEJNBPA2Wp4vBW7lMNIHJlqocSzoE8M/8Mf5fPWIESvKNIEVC
B3eEbwg9OlyEXRG9x+ssK3PS3lgjhmHddv6fXaYj/i9stVER3o7ii7LgS9UOQ0I3vCQeDqsiRJ/a
oIduarMjCBpOb5wWfryDoOrNBsVRMpt5G8/mcrw7szhnI6RXHbhvXHUYnM9hYZkStXGn5SgiS0Ej
hzCaZT+NJVhU4w79x5xiP47menzuOUIx+FegNJ+BCwFUdX4vs+8CWcipwJZrHqViggMqjDMn6jSu
m+9fOVozoKu3vxJ37t8LMEDnvMrA4bcl3sZbfdXLHMDZdAa1Vq5/kBxxkGMLN4HEHACeaQKEP5GS
6xVX7U5RkG3kG18Elw5h0wUVPf1T8uEJazktU/b/mHIpSWoyPZUyVJmq0tF6pEqsEBJ/zA67ZqnP
MqKK6ci+81KXnL4NeacUgycuuD6mD5xbh0+47fGPzFG9/KXeOIG0cWkV/kP7RhLLEFb90Q39AxXI
rucmPjGEW9NE4c8oVwFF+8oltSDO3hGAMyki28htVMwAtsWNLP9Gs9q4bQwPGdAsSPnFH30uf8zq
c+F+9iTytTUxid0vVxyEPIeL9FJLqWuc+4myBHlf9zzkF+LFd7VWpZJCEGcagSc7R+hWTwcGoOBp
sq8am7jSPB9XBFcajQJhALCC/kOw24eN6041HckgJd9RWES1FH0C2s6VVxEMDh+6HQ4xp3w9LqK4
mDEFb8NrgzlRXpw9Y4DRRf7KdjhoVXEMAvsMVc0JlKsgrl9l2dW8RWqB8hh/t7DnHGp8gKE+OE/G
0Wr68TYaHup1m+x98W9C6XyvRag2nAkBr4SR2EJK5c1vMieQbWAPk9yX9SLsst51uINgBh8FXdlc
iQErHf39IUSqIBTYSSxDaBhIrgnTKVDYWjCSU75F8nG8gwHKmz9re2jKQRk0Uju8CFPm0InntJn+
okHVC9upes9uzmm3QFf4HicCTrbOgSl1P5oQlmkCh7vb17lkmRStRrotbNDzAwzoHpvIOU5PrfKx
filmD12qxozEd+l+3hkiP6LTvcRn4Y2CHw4y6xEJDxclwoZjE8nxAatnHCZkb6zjKBkJ322U+X9O
jUnEsqGP4aYDMXs2WnTPRgurpZHmMOoq3QPxx3XvrKd3/vsJumQEDq6aeenzUbG3vCFXl3V/jmLw
BWsp8vw36hnlT5ZekMytrZ99Av3O379bPwLren+CIe3YqSPzcZyBn+ADOeA3/sztc75CdJy+8y5w
zD+1TG15kIxI9ndD3qjo/cUPo16U/br9n964LtfUYCpXgGKACjTw+Vk3HRwGTbN2L9YK46e4PMDu
xbal0ncYzTMHVQ568RchlqG7K9Rw9BWgsx4RJf4DneYcRctd3vSRIJ78ath3iZ9sTUzhd8RlY/+u
65Z+BMC2NsOMpnjDOCkOF6fu+lyTr4Fanx+b4e3Ox3+gox/WsIY3UiWnslchLfygNsyO8oI6sie0
RerSqkMoRLDHll4WV5LKJ8jV7WR1JYfI2+IXXY2ucMEdgg3C3LNW48j3N0GCWplqDG+Bg+OJy1pl
fxeyZX0Bf8j6sqsJ0W7xekvP6Px5k6bsZ/1CyRsmfv5/wofnryWq5qFBgTBq+n1QyYDvdcQ8Npao
43qB/coN5XimaJexunm853LsiHiL6hc2BWaPk4YpbL+r2KXOpN6srb7eEOjZpOxNjyx9aFITumas
7ERC+ue9ugynI+Gg3JiSsLk3CU7Fjxqy79PhYB8pNMI/V/cZ8oxU66kpxjrl+gAfn/deWSKnBZBy
UsF+cOniUFTuRv0hkGWtz5WO5+YZZrsS2tzrdnR+bQRamFAYOPCpkULdbXBbpwambLNF1Si6E8DD
kUTChwd2TgC3+sPjrKWIhpvV9TOGklhzOnmwrFgwgiG9BQcIczqp8rMWbXvo2glh1zaXw2sFj6TS
+2hvIZjQExcDmcUNa3tYvpBXX7cGXorrD66w7xqP0bwQcu1g15dG6wogaKvqkpwSCAFSZLHvjfMP
0E8KW0pboXTXNFB4aqzVM9M25R9wqpBD3Qwj25nno7kx5KmgdeGR62GMackCMZr/38m72CM8WYFq
GO+0PVMd1vrjqf8ntXLjrSqKLD75hLtD05pKu/uima/MJC43E/zIeXX33lI1tWq+az8Lhz0mK4CD
5maQjCSMveafonJEIHspsZF55RU9zJ+w/AOyolL5rYHXcJLcRrOzCpeUJusWJd4p+BTcMwGbhMXD
rVw5xVs1Z7tWZJPqlNPfBjnAcwGeA4gbN4W8mA6zvUQiVnLjcr7LgOjHExQQ8YhUJntvWcT5PgJ1
MjR9Qkcmj2mCDyLTmfAihN3L4g14pEphjia0cr5Ay+DYTMxKFEDzERy8uYTEPMyYAW0rTq//pW7d
pgk2VwKNEhf5posJuRZ/DXM9zGOVH55pnwCrs+pwtyYfzquPqHKBH46qQSCAy72xwVgBbjqehQSd
wfSYiqHTzJLvu1k48H6vb/Sl86yaaqze+F/Uu2m3uUZQJ+1HYveoDDtkpauz9/Lhtc964NTWAN6s
jryYDyzPXTcMvDZ5uiYR0IVrtjnyKXfXLk/MQf5gIBmJ1pfiI9tBWGUC3N0+8u6e+J9lHAqCPb8o
GOTkT0K/rg0mykQj5RcO6+1cRoba351tkt+aHIJy9edt6lA37jlf5eOvprJX0124ohCHpROP4Yuo
X308mmuX+03iVenPbiFZBgikfslhEus5flNn5SWBHVQd/ouXZat0JH0rkv195DdtjPL5+c/cNJdc
T1gpyND1ktf2a1wop15cjL2dcx7D7sPzz8ie49znLS/cz2hpO4bTQbwZv6l4WkO6J+YCR2yuekfA
i0afTMHCUbXMTrd3hWwu0/IkZCoVyBqq/eD0tAWdZ7yqM4rtUde+VqUYbe8Ka2hwa1u6n0rwuJj6
EJCiI0t2JDr7Uc7bu8B6zT2OXbLBZFgtpOwTJVlZw9aOPHUZQFTtAhn46tNIvznH+teu3b5GKULZ
POyNlhcD93mBU/jSQ8VougvHE2Ego4g72SFFd2n8yncXEyPnc8ndyZVRVvF5/qZEblaAduuEtCMY
05Ge9wHkEF61rnSlHKxDu6GhT/dcDhXpibf8AMITOikDMcLHlErVfy+xm5o4spzcNzn502U8BZ3B
hlZFEOHvIOetRxsXuOwG7k8wsXxAOVP0/Br6ZNBApsHMCkh3a+PWNgALMJm8gA8k7v6RCmXep//h
GYl/bG6Naq/FWJW5W1SwQ4K245eAxESOKuJ+1SZMAjW2wRJ8h3Qqi3+aQADGLXV9/5V6DTS0+M9L
i6VAZtz6QmNvwNkb1bvtL31IF7WED7KWzOV+L4BM0/fpjHXS6Zo2wxYPBDdBD8YcdTyJh42D2rF8
MrktRrE61VYX3ykAbJtcweZ/JU0yT77gJc+Y1fk+zWXVYeaMfocP4bzUVR5Mu+MfnlTN9ZxmdYuT
FScsIzaIeUYvKyzE/X4/SzU4IfpXFot/MdHyMkraURJBWActxIW1Dmxb54qYKZwul9AIw1IaFstB
3XhNIDYz6yw0JaX2ZIfyx7Ijnu4raIbg3wrUIObRlbY0Y80StyShR5ff7CoUfT8Fcwk57SNydULH
aH20OxWaRk3DbeWoxPf/gB1pOeT6XzgdfdT42q1vWNieHczk9nkFNpumnIaygUhx7pO+iJRDvhr9
+jvLfdTt5Zalxqq4yxVuGTEz/i7aekVKaJSbg0eH4f8c8ZtPHjMSbn/rMi4waR1ZztekdYUTR/Ui
VsirYAp4VWRNro/cqP5yS2v/g+Oq+uytH3ApZ3295GnF+R+pl82/HV78gUrilO3c+KzDWPsDh9KE
4SmyHKMY2geruFCmr3qAAWDSdmhHRI9FXfHJQRKU1rci2GTOvRs8ysZRikHYyMHwN7aFNKTgWUgR
3bk2ukGoHGpwZ/BEHcdSx2JBGV523fyky90w/aQibThQWnHg4ImKrxNqKzCmnDhXjnL+p+jYTe0I
Iba/BM2iCApGwfaS4I5qIIsUy25g4PcGeAZ/V+HFAJNU7TeDWVoR5Fgd9dml7umypNKk87SVHjCP
YYmYSqgDNP/0rPy0hkmahBPv4dca1sGOSWanYPTu9usTyYPcHg5NgU7EOGxJX92Lzp8woIcnswls
TeXh/mNy6v0xKd0qjmn8/cpt+ZiPRmbfhfcT2jmagAx1DRy7ZsJgj5tZJkEWtQKBsceZcCjfUs4j
83BwdAiuWuwwWLDhJalpGQTVUVQMoqwyDyc8aosNyOtA95n5hQYbisGJoX9c9RPhCWig32C70WR6
gX2GAN/DuQoAi7JwRLbkzWU9t86HtLBfoZjgfUDWvoxZSzwFwlY+YzaoF4uqBXuvgtvHy/06Rm6v
Gwe6kIskB+Vld6IbgAuTFhaqanZmwBnSEEowZACM2bsbP0omBXzcrTSRcIYv5h3k4KcXk+60BCZG
CexXwQo9+aaFjyForVzWMQ31xDFoh+9b7Lwyyjj9gC0MpdyIM6RgbBbQXwPwh92H8htM/KGiPUac
TLwE9wbMpFnupXiteaN+LBdd/KNQOEeMApxCpa5LjkPDcdW6EMnmDxLaST/e8Ebnf0AfohBGkn8d
pgYdCpPsFchGAmfcSFKzpbPqSjqJv+OUaEKtYwugZgbGUQART7trpT68gPIq+7vaLpFmi02YgOEp
jcwHredtlyLq0eeU4KT3TpPkoRYg9t0afGM7+48wQ/yGEdQTlR+RebPlWcnr7IkdrOw/YXAVXvER
oRKRnBfv29HLuNSWdivsF81PMDayb/vJsr4JjUhQEacuFLDXL1vGktGl9hkWJ05XgaUsIhNLG0a5
M1RFRsISCIcSCC1wisWz06cMu+Ym6rp9exmZYMGBModXIzZZN6zxWLstdcST3SblOMpnKqF22gVj
uxdNFxzkOdoJJM2IxbqmQdx1XfdcWgXI7mFmmbJvZQCLhjIv+ByXrObIhGOCnr2CN43AV6z5lWz9
rwc5TG79CefwkaDrPqRmG9JqwT6nnCZ9ISp4yDTO+ov7v1v86bd3u1J+FXx0AiEPpotd4UuIyRYe
zH7E9KU9VcRD3TOluzZFgSyAmqbSBBIw/y5dIwT9O3oOFEWaMWhQsoSSdSFLFJiqYzE5bMt98IAL
XavHkTNd2lPJgrFcD4AM/DZre+05zx8jisGnIRnAOwLYK21Cg/E9Xvyl1oWnTe/Og4rkkxkjlN1N
nS3vFPuB6CrDR/xaK3v2Qh7ep2D3thpr/KWWRqcM+A8KJgWV9LOvO2gezIsyhBrDW2RZGea++FXO
vWt4grrYP1s2PZzwFLY6sW6ff6+ooYB7/Phe1LaNp+cNHb8uoPDKJA7NrznabHWCYc0By+ehqtBQ
3MQitxyQAcKaEnNggTlxDvJilNrS7XLhWl//j+7Zpl32pRGx6siT7PKVuUVR6y93+oRmmiyFjweE
rhSJRGqgSSjbL/5kgVe9Tj6/JSkzJGhH6IuPvz/YF9an3Yw8+mwnwAcdqZskAq8/AkjKUC2qIhV4
WMWt9eOvqAOXJiigt1+F+MnyECxAYhM/uP5md9e10el27Srue0exJSZVeT0Wj8jZ17Ba+fj9LPsj
rJygSaobGXJDZysVIls1p5CSipxfBjFcSmpeSoRpAirGUVA82Es3G5OixaSquVLCqI9impK9Z+YZ
0tNpr/Vxbt8JSzdhP6sB7piGd9ykA255Z333ZSACsrnSZ8emF2U8oaT6LiMNXU4VNv97jUkug58i
RyAa4J2MXqy7TepMcfi3tK6z5Sqrjmcso9i8gaIzz0B4jTeo3r9WkxQ0i9D1SgMfaIfgaLabbJ4W
PVOQqYhrC9hbOz412fm5PtSr+9KRl4JgunYI/cRcl//em4QHHionR3s4Aaf7l6A+X+deNFdFEj5e
HUIhu/mNSz1Av1cvmukKTXwMOC7FYanbJq1mMhIgrgp88KujfnS8w7mAcRJVzP3uUTdZZuwgCdw9
snPkGbqTWBb4hM72Z+Riv6juMBPVe+biqWdhFh5gDd4PFHrjT22u3UMc1bsAR0nFSCdJx6pn9HQB
jrI9Ohg3NpQ/HDx1BY7OM2Mobwp9hWg52/qtQGdkrgBsvHBUXFuiLQqfQIbsdLfI3Tt/xcYFPLyH
47JWB0B9t6jiTy4tbx076ana13uoehflnHn157gAA6Kztansbn+sry8PvdPQ0ux8nbfqvSFJxHN7
sflL4fkIUBpIEPIqzZpnUXi/HUqg531UcC3VqJa8QmVpH2KILK80xbZ33XE2BkMFovHpXAjqSB3i
47Q4wSXYkJ6zSl4xqHSfOMDJXB2HYbYYqSIHYGLsJCZXq8RiprIaLbgTAPbo0xpqJo7U2BEuPT7+
3UT83/Gvntz/DUMfkX0sSWPLpwL1wrzdsMSsGUJzBdz9mjCHcAI/RxPFKnVWJyU9Mkjp5xz7aEeB
X1902vnJi31AgmXkCmzYZTnOQyeyNSrAmMlfNvRPslL84sec75I2HDxV/hgICNY0L54sZx9E1som
uKVql9ccF+My7LwuV4fLCTbTgfV8oHsAfQXamdaaOkRnXdXoWpy+uaXEvEFt1ByfdJthdkdD0I1u
MYzRi5fpJ8fIV3oqXiOEztTvxVFxcx+tbkI1IEzYhj+g3Hokv9AgKjFV5Alur9O2t3L4dgHMMD6+
2zTcl/i7aBQy2WDDIXjabDkmsWKzvMaJ++eyxcXxDCUHDHVNSRqcM0jAvSBEiWU0p40WWdZLn03E
fFGTE0H2/TEW7bCxY/7B/wgriYtvJyP5zR8817nHu3XU/wafBq1dX/mhx5vhXkw4HyAKb78YCt9x
/ypdZMIv3R1MXG5kBsk6iPNTlgIrjg8D/Pow2phKGHsSxeEFWkoTxORq61jUjqs1RT3plCheXwnn
scbUdm3q7gqLaZswBuplGBgxe05K7QW/MA4vREoE3f1WhLP+5yAwB4UEu9QfJHFzlDCy3IpSYGuG
p7ylz/XGdghEG9XaO7NkRvqGsO+HQdMkrLYECNBAyQ9i0MEyTfgTSODjmXi4GHy0ZeXMsZaVRtvk
AhdPzsCd7vuNYxV2/4v47mHaAC9gFEPRkf5cxukOR68n5+Rm/bBkERZHgoYVfn8TVHQDh9sHeL06
rOGc01pog64dibbmdEvFINDhTHH5Ube+bA+A8x1+5pImGbM5Itixnev+MnmoYLX9lVp9U2TQN5Mq
bUSvChugOhRUFqJOiMlBBf89JpPuhh/aHkBBb8ty9sDAaoVXW34sSOMlbUJ0C2cDg8MDnA1jNtWf
RnmCbjS/TIvQpytqPU/dCLkWkWFw1g5Qp97tE8QJbSUO7eC/+Zs5m+aSsoUbtW2uA7Rnq1mFnkWf
kBxDLQ6+1Rrs31BPR4Cnaj95QC/e6/br71DWLL8HHgAsX/VPJY1P9g85XGFsYaDIxuC6OO1S3Ugb
3OFRG4o7XRj2xpACoWKxbC+ikiayHuNrh10uYKJlnQch+mW09W6KKYCrPltFwiYXgEluAtf11FQ2
pKr0Oj76x9P8yp0XFgVEoBiICEnnyH2YAyOyECTlm4uzVzVZIQlVxT/iNJ5re300+5f5zf5VG7F1
FjpIwtcUeciWAZwFse/7Tpg3BTSvTW18yZrUbubNg4cm2rTXEZYD/VkvHPDAtqXPPp1P3Jbzv/nG
Xdnrv5cG1P1G419I+1aXdWi4mhTcZv+zonkW6u/xbg+HLozIlgeENvBj98VG33A5W8U0qRGVAlxn
j+7VpqtZq9AKyvY53MNZy005+929NQWaYBQt8OAsRBfdR2BOVPSETR/YQSM/6tc/rv42z1g4vnLl
9JWSKEpPDC0dY5wBTyrOgfI2kYNWYBbmSnGdLeGpsvXbrO2HHsOVwMYbEKVv5Z8qOjR6VtWDRDfh
OTeyQN3PR4WzJ+bmrUIBTeS2pzjijR84iAcmc+jmNj542XBrpCvPjGtI1H/PUWVrC0Tmt1mYCAjA
PChhsyD2yLRTdmbEbbvgeVM8ayN/3TSIdjgMdp6XUTdY9C5UmHuT1f68qptxidEwWAkFBA2FHjxE
8yzyCvv8rlcp+kyCSleafNgPzUylfP2rUObp4L1EnzbnoSnQT/dvuri1A3cK+YasGyKD6GD3l4we
tL1u+n7FSbbUknPB43R3dEl2U5hvKGK0k2qmSExfBI52fb9gsBjAv0PjvyU1vNPCpvLtAxJMyhcA
AnOOamOW0Jnu9EdZcTVAVnA4vwDz1MPxWumGCb7r9b9d9ibQGFl9Xm20sEjK56M2Ir5AL5emoYep
9WgCGVnBh8iuz3htvuy39N+zV46Mo8pvV6lIW1kxfBMl0V3vS/eZuGkaL8sdrPwgVCELgPWZn9qz
J+ihW77r7W3MctpOMcTVpwB88izcsM2xifU8YpD940P0g2waC/jx9Po3UxVW5Ku2TDZ2GmRP5BdS
FBYE1al4NJgtvdwd4EnV3T+Y2FDt3bEaxhQ6bxjBlmpbRjR9OpohUOlS3Ch2jXkJHMhQtumx1h6D
C3Gmsw+WWo4lupZMc8sTsSmTEpFimqGNiw7Eo848bO30E2rW32U1SuO+8jXxybbryo2TvFaYL7pd
7q2aiztO6A0uptmxd70f/pBA1SbQPq9Z52JElukPkxPwvzPYruQx7HmQ1/o/2RmywIdh0z6wbLTX
OTx+ztaEPOG1RCpj3mm8x0j9/IrsOMl06ULR6/Uw4/ynUApoohvScTiKM0kF7d7zZaFGILnTkTHE
NjgFakdCcZXUysftFrHCYXBl/VuTxnQVa73NAwiPxBrtRGDcsGE0RWqP4tm9LX2044/yhxxk+6lC
9w4Bs7TU53nGrsu4FKWgMnnaolpLrP+cGcMZ9a/0o1Vt4fwfiHN3MZXnAvos3aOnSo4iIIyNlQmq
2SgNfovE+3vSjo4NkthSfo8Xs7NuSRTaORiO8KeHEy1KQEMfV3K+QcsypwbfQhQVeaA1Sw9WU2gO
7yMAkM1CyXN6Cvry0jQJue1hapA5WhAtpESldBtszFVqI6uyfSJnoeiySIag+TcZn/glMQetINeU
svWPxfihGll9e/SYwqaTmQ051D6brFA7FfjmuHjVQIzeJnSokeJourQfVXGpqs2e47l0ESiKwSdQ
er6ebCztAbj30OzjIUMZNjxGqlo2aoez4tNJvRiC0R7wAuNzIUquyIMbO1KbXRGhWm8lZwctHILq
nWhDFrd7r1HXnZwhecGg8fyRq6G0IFVYgrd90iugKNVSe0fmwBDKV08p6mW8rlbT3hnIGlOa7r0g
fqkuGXOY5IHTahlgUGgRC3A8AtGY+aa1B9XIDuCMUFr8te4Uy6k6XzrO3zYg4Xor1a7E+nG44WOx
4+Be0R+NlhDWlunANSWwSWWsSsDQdOZwOf6VqMNmxDavGGS/2UmnmU3PfKAmzIDO3saJZfjR/TPW
fMllLwJ2mTxCwg3TJbJsO2gSUDZUK7pdBXZeN2VG/TR6iSz9cTZaw24SPQJeesbSma2DF5xVVMYl
pkEQfFsJ7m8fiqBgNILdeTxxZxE5JeQfJ/48BLiOWZkr/Vhwb2sT1L0ETRSiVO+lpvqHbFp8/vZk
757ApVMTWDkjvuiCfJSgm40cSFUFw6qUQtR6KuCK+AQCe8jPu7m92L/72xCxooyUAhLx8Hsoq4iF
8ZgMwmCdHYsF1xBuEDzk4Cj7u7mkj19j1GpA8AaLUJO9Zg3Vukig6V1Wxiz9Ss+WeTsDvNEat61s
DRKlhVMEcYSsrqlI2yT0ClYDhmbgO6dyzMWoSAtTrjFSlNwPfqcZElDr85/9W72qJa57O6uB9zEd
+M7S1+fAAp/c5X4U7OV+QgyxFIMd51Z9MlPM29ShIm1G72FYi7v4Q4jQnxs80h6nogC5QfWX1GC7
IHvIB3TNxadPtbNiN8nBU0tm5zFFrX7SPNOJFcq5l4hAAqOSILbPVAIysM0ulmkiwfwqrC+LqDyh
ALz/MX9V+AocYjHobmaEI3C8OupwiRQjr/aVRPbA9KLV6fu5+hbTkLVW0lfPKYN/e9go4QaAY8QE
xri88LZg7BrNCAtV14JL/0IS6NvIRiDZcR7cOIRtClXbbw29o8QI1ego/kJdOcOTa6Sqy0r6HLFz
jh+2JgViGVu1eENIqh6hJS2y1oohJs4gNrbnnOnCPh7BkzNYDlJl5GaCeyblxgu7GXIXq3tgxLfw
2b19aoAOsWYrTyP1Wy9HacaR3O/OYaVZT5EJDfdURPREPOTnrPeomDYrl1f+501OQ+gK9dqYRTGp
y9njRNopyYjivxaHObTMhQIXg4FPofz/M2XmKmnDr2ZE5TF9dYPQoL+1NWjd6NKKln+GnUjbn7NA
XESPpg23fVp1COgl9+KgqDLfhuNP5j+wrPpZi4yPyd4mA1ObBq5LAMZhHb7859te5Z1FgsY+noTx
wu/Tm6EQN3K56Woi+AvtLBpyKtt5l3hea4UpPlBWjNJ5bfF95T2ZidW5rs3Ad+41Nf/Su5HFIuC3
3Zeyn8Gxk4Lj5Z2T1XuSRjMVsWO9tTy6uALcJFxl4CmgUH4aZHO7WPU21eNG00VIEAc1V/7GuzI6
uHGRZYKDqThUI9M/CPY5auoEOsykb2HF0/oNEW7TrAs394XmxAD9Oxwjj0KeHnqF/lo5hTUSbcwa
uU0eushQVm+FkjczPormG1s90NGOAf2Y50ve394XWmK3feyOUb2rkf8T+/6bPfQlMJkyj8+Samz2
/AHnDTBavGmbq5BGk198dE759u/mMnBhOHsN7GBv9VfNSZA9BwA1iZXeBwjANqiOEcxyxv3Pj1v9
uZ4uUOiL0UGqfQ8tyE3xmtjUgmkHLrRl3S2UPVvthtr/70DBVxHdRMuzAOc94bwpM6UrnfxvZEDv
Tag7AM3rb9TKD8Mk7Hut4fJaue2SjfCfGVCMIPdlxQ4QVfs38u70MfqlZjrn9oCcAM+l0xC+2QuE
GQmgauN2qVPubjGxmVLckvmAt8QS1b1g+O+AQKkrpktOQ/pBKaTFml2rHlDXO6I6Ghn1jewJlpcd
dxTuUnb0ZmiEPoT2+qKEGfcE0zbNG2H86MEUynaorIvrcRPtGM7gVsHGK/kRCxFo5stFq44R9Rs5
ojxhPnBFrCAndo3wubLdowLz7xCclioD9XdD7dKHgnNYLM7QzXZq2PQxXgwGRZlLu+6lBdfvJVBY
O95OOFc3kiB4Z+nEVYKnUjgnSMVBRuM/LNWcN1BHVEuS0mVCRFqOAsvQb7tubJrUQaCbQHINdH66
LCzKtWIIhZ+8FXWMkDhndy/fwpFtC4v8h++VmCWV2YTQ85Oiig7Gsxu1sIT8uzIDgVAdixEr9ki3
fhLDqoyS6K9bgyO10fKsXXfgeJ0Yi1ZvT77b5jB8iu5fi82l09mtl8oP8qfP77ffXWMZIoGtrbaK
JdQmuRSYVeHhHrlrLzHN5aUQ/AX+j4zOj7HlRlW6dxpys9H9ibGZUo8JA+eUx9lRaooHlbqWKH/U
IcjAVzjstg63JqwRMd+FMcQn/pu0bgbCd5aDE+KphleLCK6PfYknanI7ObE7Q4Zise2dvwW9CxAc
Hl57Xd8xPZR2h5GFM9nsWC0rpcJqyUICSouCoXjUl/QMopyqiLyF6GhmwTsgmE/qk8JpPzM8Rawo
kdIog10Dtpf9Jj8gu8zkmCVIGoAzq4TRGOiQ9FtwNiF1txs0VicF90VWLyX+bgPAlS/gWFYRis6g
4YVKBH1tuvibdzDSA3xsaR46O5HvboY69R+EUGLHOhE1EjljtTH83Jg2tOlLMafxlTHm2ClX7lc2
qhKAqNqXo4ehs7pTYp/pzcHSmaDwBK/uDHhd6ezcwPtjfgb/wKvM19LbzssFTpKolwzZ8hnjH+mg
UITVuDDm/TUo4NaioUJMScxK7cwid7B9nGsxXBEAja6kcEIlqw7ywxd9TJMthoTnlfHUsti8C4tW
JSYwxEYdQS791VaUX6Y2xUv3I/EHb/gghgnq2mgAXTuG7MWXS2hQshfeHxVbDiCT6qXDtFJmhr9b
qNqPAhF//OsBdSfOG7FBIKjFddZO+mm82vEQF9MvGJoj6IUgz5+PjRySBzOfg77JL5l8KFHacRMS
OyojWuFSOf2engG3iNqvwB3xendQLKzeDeK/Ww1sAh6+aeo0toYByez3h94BDSGuJRJCAEMX5t3c
nfm85sR3CZC8jFPzDTkTuReSklOlrpAg0OG680aurHYIeybs3J5wBsSt3YL0gZU7S9ypGoCqj0kt
tOExECgQ8MZSiwgOUIY8oUc3apC8MX1pxSW62GNAQZhxAeAgrK8WVIlHawQ9JEU53yZe1yZx6PEX
n+P99tYCKQswjk5pnJsLHmbZ98hknUXxTaCKGENr9hnlGNlhYbeFs3x0ZBoJTwFGg71oJZRE75zW
vhyiJyKsoo5E6RYYEpMqdMzDoKrVHlesyCtOAp3FHBL2/aVmw85dDw5T7ArQzlurHRSvhl9Em9aR
G2t5/E7VpQ1Pkb1C6b+L/KVwWgMUkt4JgEDMj1BG3+rxtwm7z8n9mP1EOyyAmblk/sl2ugbu8PHi
K+OzLSqVic7/gwablasE79qYYwM20Ii3gbN/EvuzYPCSSUGwr3u9s7iDDK/TQb41iVzOstED08oT
OLpwxvkwHfW5AQqp2iF+t9yq0FRmDIvWMC0qd3Sbn4x4+iIBxOD477mLLBBa3paFjM7C8pwQ9Dbq
lCsvIlRfu7e9RtnMtxSCo9R1b22Bjqk+UKaNKxVkty8OyFxkabJHmxSn9CYeyQBKLDVlkUF83FAv
W8lSwyiMy3a094n00etA708V8duTvq+Naa4s39vzSbZVyrQkCn8Tv2fSz7NBdTuFMmnniYpP4ytz
05SLn6Aq0J4vCIQcqsSsApotKkaMryI2d+c3HDnz0h3gvoIr87QjQMnHBJMIXiIDKZv2Ubb9tu5k
s4lGC9nBAEgAKOCJerTCqwEprBLjjL3SuIViWpiIg/NdIzXEfsA9HpyXvn+fM6JHaqg9sBB4cz6E
RiyPRUZBALh5JCps4Cj+F8C181+jF6pGK0ppfbNWPOGxQFT0EF5peEEhRNE71dVbIOyT3saIeKAH
2aDiiMaDa2yEFPTeq+XxF/2RuXYGYn251rcbR5fZDEqEdUmufWFjtomLOrmzL5E4P7T64cY21weN
NAIeX01R5Yfnmf2sFN/Gbn4vB0WMdeZrgk0AZHI4gePGxf6gUymci6kmiCJ+Jsi3XOqYmCKQQmuo
UkIoc6NGp1nFz3b/ClcRlAwpmMkDZhER/nG8/Oe8pR2BSe7CTW+hQoHnd6G2JFCcEtmyN0FTMvxS
bQXtS0A0s60WTRyfrWH+emVMx1qyvqGCg3Mel3V2OEXGxwdsS6c/swCSC3NIIw6b+6OiWZZU7dt0
W9O8W/1O3vU7cQA7Fbu6+A17WU13kzZwpWLtTTALUcLORG3/zw3h1S39Roq/SQQe1iRtLx5B9p2t
zczZGLqVMJXn2G8CulArYi3pcwAytlL7DZF+W7O47x51UnadPaBZgLl1rj1J6M0SUGRVCiUTaFha
UZLrnvnyT2BJAqrRlRryxXpLlrdp/l+Yv5AEa18xl5RTnmVdeLH6hQhQ+BzB+hkYb2Quqvykm6lj
8xsYyp7D/FIzPgBZl+X50znr6pRl2l9LcXsIkRQ2XGDZjTIvzOPx+llEEd3Bqq7HZQ253C3V6/hP
ChH2TCMhjx8OkqA/9rBDsBcMvSmut1rXWH0g7+pm8alHF7AXdA2XHOcLl18KK0YKb3ntXz7MIaAU
MozH7hko/qbWBaxcUJXI6t2+GFCKAOkBZvdD7NThvYZ/qgsxMAb77pG+9nae7zrv0sPiMKnj+asb
djP+Rv0NKxOyMRkhQeNrQfiK8TbFl+RL1wRmBpQNCWGEfESKPt92Fn0gJA2hwfbBQfAhDFu7nKpd
gA+Xdj6RC/XVGz2y/ghPkw5AU8r153hK15IPCquvj7JzZNlUP7oi7X1Mzg+WXhhHECuLpt6IMuxm
7wb+Au8lxq0fnJRlczFyzXZZ96DN79pmcQuSvcV67L65J30mEmsXj0y/6msU+zpswO+YXLk5qMle
BIFy2wtvPezgTR4AV/uHR2neExMOjSVBHoFCxU7If/5Oj0baBQnQ1L7Fpes9fkfV+4agBbHWZ/Nv
Us0v8LZoJeBwjD7ljxUWo73Zq9tDeIHPAVAcfY0ulYp7HK2bgbNMm4E4RkTW1kqBHMYM/GRUinM6
1WBBt3q391/K3B6Tzm7Q75opcxDslK+xwomBkyOoyhoEy89uBoi8RTRh/Zc2br9ypt/6idTlk8oV
WmxG9as+C7/aT2dx28h+kyrSr8CGtEOrRggBUKIQusrMy9bODcoZnyB0UmP/zYyBh8ruJ/hmH4sr
uJULHzhtpBMIjnPG3EXND5ON8Y+rYeDsNh/rdWBSAGKIyM6CxL0MXoNBnKF/jb3WngzQkNLhPmDi
+Pi1r1xS2yAmVE6xXLkc0qpdyjm387tz9DFoKe7revrlsknOT+ouPJodbWbyVgpSzygdOzKnFvv6
OV9h2gjjrguR+JgpmrKPLHtq1mbTyyqb63rxrRd3wb/CtooqGNBedCUsBCiVPUhguScCA9gKPsFD
mQQSXiYv6C2HVLfSDJYz0dAhiP7iU9nMVULy8xVdmp7TPnPUukcbjmRBfGwPdiBE7rqykSUAtvyS
z6Pb9K5E4M77MbDz783ty5oQQTfm43ftHEBqdlOGjUKWCLjuD12kPSA3g/s+VNMCaWw81wztOOk2
09v22MzYkvGNq55Qlvo3Js/R6djE36bD1YcWuZjrYrfZMBCHsTYiA8g9mAtz0I7vYVjZy+ofKrMA
IngH8FqGtbIip3pRkVn/u2omGmEtXZuZrlJQsGX/axHEu6DawWnpkM8ihRT5SMD3nZOIAcC4yAlN
UB7/s0+7rO7qB8n+3X1MbdJGrWMr8upP/ItTx5PsUtPvdmBpWj6QJLiRHOQScjFa8vsAGHlChnhM
9J7qobiXds//eMeFwlYdx3btx199LwKe7BEVVttbc+rmOZr0CgB7WMk3/L9RAVtGijrKYdPnhAb3
Grlo4krWYekUq01vvkASUU5KBWfmLMUCoLyV82prmsW3eVOEdWAEgbDZJQW9avX/B6zH4IU29m5p
y/DGX1mI92bNiuphO3i4yjYOLdNAzX3+uL5deU9ue9aIIZq43wGOijcVWQGT2GJoWGqduVaV85vp
GNCmYY5WVind3v8BGWrErIL2NAYynW8xHZ3Fxcla1ePkQWkbDE40pVyycZmEgMNLEH+Hy3cKz9jN
PfNt+oDOcmt2VDN+nBiL9I6yLdSlLOKS+KmdHAczmiuCROCTuh91KmoPnGa0P2S1g7IpijmMOQcB
RoqIx8YhUlL/Z0/KqEcLZd6s6Z51GnZ44LLRh6YZmStnnhBnIxUwBxCeTfpoydurJKYtxaLZG2GK
u/izOVAFUGzZ2LJ4teLEtwWAdcbZJuoE3rBtSom9kDUBZ3WBW1Y9AarpFcYvv4Wa/HMUuSApUMq1
L1ncl9F0swj0qwc8jolfj7oX6gbsBGC/FveYqs0+LYfy1EspkIpxGthJYwDgshFZkFfG4f5m/vP1
qQHrEdBmVrMWmpj9O5W3IXeqsjyTlIdZUNFnotTbFxK196R+9FPJJA5BM8q88T4ZSM4y+3ND6ZqJ
GOsyh6NTA7DIB/WfDl71j1cECNEcoTQYyQ/0jEhKfs9luBBDWlYpuiqGOO4LQGPTAM0gkoITAUp8
0nHhY7er6MrvF7DIVxn8n9dSPTARTywObQg5ab0FGwx09kcImyW8KPvMWf7L+MxuJd9ViYJDkzdt
+a5Dksk8aDF/8/7oIBduBCwXYzoP+lTxYiX9ctaZ3jOz5vROoKvXBT8u+Mj2j33ZMqkrvZe4CXkx
sBr9gObqicZ0KdwNgGpAwrFe40/oEpqZtHIG/RziqiGgAPOYBz5YINOy1BOUoHRLsLLGyywPfWb2
YBq+oki8vQ1XScD3F940rCnEvQLMbmPqhiiEfF0AgOeeqrNZCTKzyQ5QWV/m8+g/y9HQazSmbD5k
elCRytqA/6E8rkaulUAFAhdJjDo2rF1ppQ5TsXf64fApa0Q/RvLXqf8+JjVkfLLYGQsE9nkewoc2
S4gZEE0Ezlj4kENi62Ofh6GTZd/b0OCAnoo8P1xrwqDm5yRaZ5irBhWnMcAlczg6Hy1/kT2UNNgD
Edq/sx51jz6r/rvnQE+bbXo+2WisX0MtqvqsI0phM9mhMv2d2UhnKPAmrv9Tm8MGXM7rCr6p9dJP
H322xHN49FaRYGNIEB9cp26khKmpGgh4/t+5vuTa2Uo1bvImBoLMZmp2HuTDXg2Op36aXK9M4caW
ROYh5Wyc0/5Kc9EB+wrV1BHJj8t+vcUgafPavIp/3fNvdb+x9VAWNJHmpn84GhBKMvk6w4BwFx3V
k9rp+EQacDX5M0Qo/Sk0R4N4fC6+XX6UxqdnjKMTNuMCnwRq5QvWsHnaL3FCYaQgo1b+RDFn9NWg
iYXloqQeA3RUjOTCYpKkptOpeFhNXWTAaNYSAreBWES/10jgY6CIsF5UHC9XxqyqB9O2wgclDPVF
QGIRLPCbLESXMVr8bLtjPs8T9q1p0iF2UA93rb9g2dUXBGVdFY0j8Y/1c2M30sHe0DhvfKm4F2NQ
YUTSq3X2AvvngeZZfX6FTlmvjOo5o6E9UpPVie3bXCXM/s6elOidFSzVAzJgQhPEA4qs40qoz0Gw
7EklpIPeaoxMvsbOa8p9qTsDoGE+mLdK5ZLSUGqfOBF5SA3yq6AWR3HCTh4GfxSUlGKzWvr/NMnI
SkF+sb8ceiqchyp/bpZQUUIel8SghDzXBE9snyDy7keyPMAY6WydU2Vbcjg56eK5zj6KP1xiWRZs
PYnse1L7rOGnsh1jq7MwuIB6473NdnzAnJmw/XZGAOovHOi/HACRBMXH656imtLGhC5pDHcXcVCl
htLldYiKh1VgIIGOx+E5R3BLXcSa0VGTq7K0duWwp9TwlcGgaXYPim7ZM5mBZr4budO5D6zilN2B
SEHc3mX5DPvt46GEHkGvNenLjU6r21wHtqpHhB3adVXQxIJz/QgypszPUrj3GCKEIcPF1ZbLZnRl
gF2B32/vJJ3C9TeSWwf8hbcJzSBZkWTjA+aG7Djsd0fmp4qTjUzmrBHlPg73cAVb3x6WYpbfHEbx
mObqiF1D6+oIV9qUASanbwEIeouXg27X8Rcp2WAS/D6f+0nSm2Ut9frKaNNRYS+/Fk7jf5drOVuJ
+0IP6GJWotPkxm4feccGehw2MrN5TkLLqLKun1dv7jQ7kDO6WTVU/O8yYAMvRG/4pFAtIqGmBSf/
+ao47LD5zQADKOBoNigAx5IpGhIM1pD8IVwXEO8wRQFoziXJpPcEd3/BQk//0YQ5HMcslmaRjKrT
JudgLT8Q2eVHp3IvPALzefGxy5wkNBDWOsJgZioDQMkf68QY8TtKufibpa97sllVfSR0Y/TO1ABc
dhn0bUMcrA/G/0rC9rZAY16DLwOMjKaUs+OgEwyS0AvH3nSRnoyTYJRElWtMRMxxln10EoJQSaH4
Pgc+T1NtpkTDIGYv1dVhQSS9h4wgNjBkMOfew34MIBXQjZMYLmnlc/k16UWRoNotBW2CuG4LF1fH
FJjc8rVAkRPR/QEWH4q5JzqNzaD64DFF/GlKF0VXcGUhQmq9Z3w2d4FAkENOe9fkCiBaMRvLSs8J
zsvaS+BZ75dkwnfYPLyWu455xvBcRBXSjuENbCXIhqt3bh6VVbmCQS321dowE7fga0SuSR+HTuA6
GTh9w/Weeh+wcbLv54iQGrYhZsiB34A0uyZ1mEqtuaI25PvRipusM1pjUxHl+LVIaRegpAFnMqvU
UqlTzIGO3DrdxdedgXA88v/7uO5juY45/PIwz+dBlPr8XXS3Dt4BdpP46MzEngbeOZGLJQopOp8i
stJbhCCSpnG0n2Ld0p+0cigIt5UQVQXbTON8fyrl37Gyma5ooBff/JTJwh8DKmr7Y+N9vgYUlB02
cLnHe60z3c8jjdYlwGNmRbDyyZLcWfbFXrUM0YyYlbj5FR2dSi9Ufron5ys9Q+hlv8W2uZ9I+2Vp
z79zD+yvBAMVUpw0sHKJxEiLUrruE1K/4jEq5njhQOsafd7wykV3iu9UnGJk2YjfrN4mKel97KbD
erCbLcbbfzdfqBwCuKxBr/8MEXETFtDKhchX/i7QLyb5NZ1ySstsbZ/cwFSmi29CqbK1PHgV7OxK
jbe8QQ3KhA7tpfcOmXdnqcY1taFV5m+MW7WgHs0L2C7C/4Afu49po3UfYk1WSPy/nELKoiEW0SKW
83Y7OJ6qEnfXBvq0OEPR7DjOZhJvIo1IvQHAaOG71qCgLmXME0WfhS5H/nCTsmnrbhMQLOJfbUWf
DxAfJZFk4B6pHwHlSRmwh5+WQ5o/wz15TNeWowaPbVD8cpGo2dG0sw5SX7lH1ra6yixxXnqSzVd9
/6nfxq/d3PP46EV6PPFiny9VRLWbyn+MvmhP2r6M6Jxajm5ucSdRxvmZAj/NqIU/zLB+Gw63vlZR
1FG2vEjHNlk0OqaCxLVX8BcYOS5lqOHGR9ENvNUdwsgdbTOUVT95XbZRYbKePiPw8VoFB3xxP0xg
wzUUflYYj6GAqX5VETXaWAjQiri0t+6dxlp2ekzY9mn6h5/Ck9d/syj7spxKHSqWRxXXsWDjOYP7
U4QaJ8039X5S2Y/IM6O41HJN8/qPW1T75rJSWIh/8JKE9WaegqiA7i0l2FAdPcNOVXPlGgL06jBy
avhScZrcO2YCgwq3jMd9yQyfCEru1D66znd8HYNhT6khJZ8Ac3/dKQ5poiyBn/85zrlDs5Lhh337
rawhzBATeaCxg5QXi/5C9OWWGd2p2d/o0udEZBAXGg2lD6iQ96+/uk0c/wbvYFexISq9TdDBbYI5
HdlJOdUV5M+M5wBUAsbz18ZO0D/GejkFP2MmCoJJCyFrLYkzzg++LPJDQzwywK3uWr4572ZYgsT+
dBepf21TsORZbhuxQqSlli4sPfdAW9V9dJU0z/w2y2+/YzLtqynA7ujGm+pEss/85l5LAQC5rdkq
2pcVPZY1V4l8IlDy6XCGX9Mk1Xx9sFKoVUaDpsTWgnCCI7LQKVFTPoRdE24vOLDoPkCgjhBi7zRt
HiqQcf31s/Jy/Vh4azffNmIH/ESTpS/KgHxAv/Ok5ncvSdMlw+cRIbO9tplg2ZAK9FaAXKVEBoW9
m4jLN5bNw8Kj1uEhbeUldUYPmK+z4CZitYTMxVAuYxb6utkuY7nRAL0FW5Yyw722Ur+/M17EIeSh
bpcMSgnKBXYXd3myIZb+b2dEVVgfpPtrEm2YenQZjAQEST4Fy9qHsutwW4YLFllLO+iEQHmEae/P
jkaodOV4klCMuN41I5OKGQ5ljWbeHPRvlzkssLq3j/uPsNgM37GFuwi5PZmEuCp3W/2r3xiEn/vA
22R7cZIM4l+H505D9WxjIm2Gl1nb6/WAWMT8dSjzWC5nmaaMqjzydAt1w0Oy+XGrBHGhmuNXh6+1
vIWF7YVsO9pw4/OIRb9/SKLK6xpmcAb7dAkfGKzaFyjs4KESBE+emhbAo+PjXNyyKK76G6Pq+AFz
Z5QvppDhOROKgkYig/BBJ6seo3qlwNmCTWotjIUy9T/rea/EWrZJPwQPFS7jPT/bXMPNJouz0ZqQ
nEg8LoYzGNQ/4zdV6ZOUiBw5wplGVEWr00kzTXrXny60aMfQ0zwzGXahqJJMAOAv0Xdl1ATceDtl
cm7vh5sVE3EK2KrAJ7Epe4o2qZ9nyBpI30mhMOw0XNHU4USTkTvZiSb45CcRpg8AQ69DiCSO66B9
fsmwIJDpOv2z0oslQcTJBoXhBMVXkQArfcrcx42vyeCeaTspRluWbLEGsVr4wdbahhRc+/gi03XD
/FFwksPBdLO66HQwwbuqRE4dUjzCCziM/hEe8o4+Tfztz/AQet9gSPvKwbBd+UQMciCNqadE41kb
dTEdrBU7re35qcWaxJxQypo12mAt2h0QtPx007FCsckZb03XIt/mW54kDkXNQFhGOt24fbm9hDrk
lQLN+VG6FOoXqZJvt0VmeoMaVwLu6u2tdZnk26cqPgp2bZultrOfPljqIpZnxVpT6R8dyg49U6Al
ZFlkvGlZajaKQKhN3+8S63Z+IYMcc55VQShlUGSQC25Yu6hzV17cex+Dj2M+m6BqmvDKbGf4px0c
staa1FAiJDXOH6qFaykKbq46jCPpenOiRmwTNr+HecZzVrF2dql1fHYeKVwyPA2a14aynUR4OaEF
fjDEonIU6wxGYvQivmC8Oo1Sdl11OlkMnOvt48ERJAMocnVpIOEVzkeVitoJ80GkHKD1RZ6mOLkF
lrUC4riA8GaK7uVP4jjKwvpuorji8Y+7ti7oNmsl99qMjzwLvYT/JQCXz/6MIIAHbTBiXZbT6DFK
6nsBmbgdCeaN5aG16LO7fEIYjDvwbuyjZHzbQIi/n5FM2e1buG92kAOniJqnvtdUNI032lpRg2zi
fwHXReeKML0QdTyl8/XTuezDSLSRpDV+hURHByH8wbAuECWJEPFVTbn8ir8u5cMe+aYCLPJYlrDe
w6HsJIPjwv5IoLdqR12Bijo9S9TjEzO49Ahz4MFo4BeJEdzQmBDVA+OguMC6HimpSyy1MwS6XPCL
VD0b4sO4+eEmCicop1uYwbHt2pfFeb9vF3oLzXa0uQwfB2P4wDh9cavzd11p3ccjZ2JiqDddjWF1
BOIw5HRxJkksGKQ1s0CKU4KBJ4UUGRhtb+xhq3Pzqb9J6/w6uM5CzhQuqfUb7SatKzmjTUJ/Xz4I
ACN1YhV1lA6WOfYoXXrd32/Bi5fyyBt7uNwmIgxZw0wjrw8EdR1p3+l2weMbGxnl71xCb/TrVeVJ
Dv8eQFGW4SoXxzzVBjR4Sk0zR/QjF0ci1GsxJndqoXIVNXqhN7Q/Wzc9pG4uJKrLpd0Lkhkrv8VB
1Je6j8gpZ+IrEmhxunVX4+uLg/tXRKzPingkmTMJXzGb9A0dzJvtXlkCdpCAlWAj/Z1KGQpT2D4f
pQG51wSH4PY250R1dUOKLprEreprqLnygQtz5Rg5H/XHOSwKW+/qDJNpG8Y19GXzGcjecjDmIHy0
ONv0g8vv9qTOCAMit/ZQEUNO1A0GNlCBAi9uUiuvn8pRRs8osAZkODPptD8f7mGotuYYQOIGSHRv
jTdqK8yiDEIKvBkd9lG2EGOYoKWdNTuOj+X7ol4w64rCeeuxLruDRbGniVojlNPLqIqG10R8ZHsx
V3Nn8L5cY1IOu2EuJXbJrCAs7k6Yd/ZrqTyYZV7bmoMT+VCWR4WylicFKhI/mF50fPV//T2b8uSQ
SCr1WRFxvpAxt6Ih6MheTs4xHhngKAVq280gQPxGVrZPoS8iAS3QlZ21Xb+uSViRWTswF0vnGCOE
XLz2aCm/EPY/d5kzBSMl88rvVj/AZyODTkX6qaVdMexHtCKBBJ6Gy1GYtcVBJ0jTNmLLLAQSaGKu
YzGKzLcHNwJaQXwSNlDpVPypJGjcuMaOFOk6GWh+ZtGhSe34wcnDXNUdFk55zgH+6Kg//fpH42JU
HQ6Q+8yGwmN7xHt6rKLK1SGhiAY76L+GngtsZK7xHp02nEJK1D7AQwXm1sW9x6Nx/5bti+tynERH
L8z1alm3I1DOMu1htAwZ4cY48wvgZn8nAlEAt/rVohGrUlMh/yLLdJl66us/YcGqmaEJReYnJeF+
L2e2510EU1ZjKHikuv8y5RiRkjbLj/1qMD/usPZrB4BhHNLyO9WLnJlb8ldwiZa7XUuWXIMD3yiY
mDWNJlE3TXBGKQwHRZoYVHp2UFbYMuP5bpDr9GjJcN46VAFnNCFylLkHmvHTlq2oIRf/js7wqZ2V
2d/FKIZS9zk2++SFrDBv0RzNeDcIdUfIAhXUGnKo52nDsM1kS0ed4r7PKKd1VR94mWhPAccw23z6
zyDZzAfXbaeW3ZIWGMS53/55GSuq2+e6CASaaExblYSKn7Z94qGksDDQ5i/+iE4yqqn3P7WRuJVc
w6H9ML0Unphf+U3JwY9iJeLj12V1sm4OiAsNolt9pHae5RJr9XpkpisiaHwVgmhl/frHoS/RztHA
Qo3/LF9knWVPBMNj0YQFNUECJfZuFE+wZeif/wP9lbvQKLLrZoIow/gTPOVeQrgXrw21uBTVskth
AARBwJec+pQeDsLuPDwMmqDSRD8vdjZhWYBXjxx/ZwTd+20ROjB8GhEMcYvd0KNLsks6hj2WcxWw
YdMEi+LXaQt9HIrvxTveBruIClSXfB+WevjsQ3UkvDvUJyRFKAC43jG7zKVvbH9v0TcFV3uslIhC
/j5Aob9lkJ3UM5w/TGDLkqGDFblqucrjbx+h9fzLlflZHkRaYLuNqLT3XH37ovHlJrjb0YAGiOnd
rCHYvNx7OXFciNKJ9BP1ShZDtAKyfh2VRY2tADDfvBWLu4lhN6tnnqC3P+3NbkDukdLtrZ/SvCJO
bAbiyd+tX6tp8DHacNzXxCM0xnrUbw0SU2e0NoWWbeAlvljaIIqFmlnGBP8udszt0n64MlPpU7LW
9DPXziQXG0/clgb9GzRVnZBvgsyinaafEim7B1OtuZtVk9kFsgvzWQOwjhuQb/GmrqzBB8KS/Yga
Srt8AltirRRmM3oFIWySi9SkO7jCzbvpFN1Qy8h1WbvA2+fLrmuaBFDVk5duHEYMXjqWQJjeuyfc
lKOcjpxk24v07GStApD09VCzK81FBoctLulEIiJFz0X5bwWkNa64+H+38zE99xxBv2pDEgFg+tYV
YAmDMqRTVHZPIYRlpe83nWaMeQ//QgaaFGFH91Eg9HaleK7D05NugPdAL3FVjjytRD/flj2nat1E
8Vp4avQ36f+Zv6wtIvrF07CbyYdv2Awm3NZeUQOsLPbKLzFNke3B7VKkRdCJcbq5k5lqUnwsvPDd
JSp7J+h/w5UFhCkXPxPKSbbUl09ISNG+mqpT3P6XjNrvXWu0qy/fQ4CuVwGqxwdFBn0ZPJk2YIto
/hYuF1g9UfQTFtzCG6q/sEFIEqIg1EFLJFqQIuF2A0wVzcFwzxfxTMgXTUwzs6N0U/KzvyF/oC47
xPgVT/da1uHQaGg2kiKSIeq+pHH9yo0DCm4JXmyJHxvS7J1gqg9+IY6VwPNVvC2CtAUxAF8HGdil
EJ6BnXO4nmHudEmr9osaAV1SRBsB7caP6bqYmy5KvR0KuU1hX4HU3lt0uXzgesPeu5OON90taZKh
waybKNmUNcLUW/fcHZDAdMNeA6qV4RmobnUYEiTNfmd32n/mARiPE6sbC1krXNMojlxu2MFFtsaw
DiO3O/To40gX4HM9qLSFZV326Dtc8X/BIAStienRkbE+qyUBVmlk7O5WCqD9q+AQn8kvItmSZTkK
JqI3H8fmPLj3lcznqH3U6kbp3daC8VmRbc+2WLYwyjb8bzb/Xvi6wCWM62u+kGJX7wjwSoaha2Id
qQFdHhdXOucXOG3b/i4FsBGPpsLM7CO3vmFgNYuLqXtZHFcJ2ac7aXf7+AVnBZeGTsgUbu5P/Hix
RhqREF82Ku9KyPaQTBZH8ntABUli0xNCDz9Jat36EqzawbkkinLlMFXu42Bl9kP+cdKRkLG8bSgI
dkYsp66boHDQZepz2XW7EzPetmoZNtpo5DEoxyI65KG1u8B4yThlcEezUu6TOstk62dQcu1n62Kg
q4Y3iG5bRZYy5Ja5Y3w/a5b1vu+QHvmIrLBdscj+KAQts26QJJfytWJK/sQ0oGbF2BzEE4syfHja
BGoCLn/h/Pb5wMbGYEpiZ4azPb22mUB0FCUgdqsXv2oabqv/Ct9sg4lpb2Fnjw7N7PHG0Y0lsVAh
AFEYYZ9NT0gyDDYvyUyAP8kaINpHqS3Gg2hmdbNO6mjDhBSMDkZraVLRmAfuvW6ArziOd3YKcbou
jUOMGk6hyDOnhgDM2gRwUd6S/N/isqSfyFZJCkgJHnfJSVG98WUGOcCUDc8u4GPptYvndcpd1aEf
0ZUWhsYKprRbdZuczDd054V919G/2Kjv6S3P41hycXP3Vn6ruHlQqg5/Yu4zB2Fqg9pCzqS3L5WA
6T7Hf2MXBlFcTW+vg+giOEdisyX5w6cIXUgDyy3tDz3NSykpDtMJ8zCbJ3i47uJ/i2cmu8AmHfj/
tnLi4C1crlJGC5ZcDZQMNfdspvrG0dLthUTPJ5ptHfSJcZJ5xPchdhdQlWdRR2IfNAmtBpDP1vjc
C8Qu49qRgzfjpP2njaxBRAMkOV+TkOHIV+QGFG3VHrA8Nj/qJuv7HY61iO0d9xsCAf20UOXz2RFq
XXt84unm8xfKlzRPDGZ/vSQMkV7YMhfFkDywNKPSQ15CrCFQSnO1DDEByCSqvEL0sAG4nRKtGqlO
W0jn9h1lvAaKF9WhGEvzOP7RRCmFk+PKiPj1TfXWtsWneW2X1csjX/KgwbfIYnzKdrWF03bWg+Ju
EazFC5/eyVQV1FwAp4wrKra29BXaIU47Z3DkWf9Cc11FshCO+lJM/IAN2ZNfAnieO9Mw4HZTILL3
f651TLTPKMTibgRXwMgNM9mmjD4Bw3J62iRZpOL9ck4umgVSquapmX/bxqSpmPSDHZuaCCnnoTBm
KLxXAC3ST/B2vCKSfwn3JNzi1avQR1xQPnZgaTuGW56Wr1rwlzaRtWcqMvDqr7APEJ8xKMGNJ1Ks
L0H1LxVc5JtYrDYAGSwo+m2vZOtJBAHiHIdpJE6ZuSU86T72CTV7X8my6wnB5c9s/lz16wiRvf64
u87AY6cpBuF31d3DE5MaSRhXzr3TwHDTrUj/5foKFXngRYhRvzz2MWqzq969KpT/W4pVKRUGY6Gz
glVWVq4CQGeuqlsRxz0j1aM3x38K5Rq3NgUnlPgX62KlfoVede5Bt0eIhJdwyiPS4pILPbraC4f4
Nt51hrtZTQTzEUN6k6FO/U1QzfFMgzVvXQSSvvps3Grn4t9DYo+I1JbFM8lQDkXoGm77a1zSV6FO
UJxqZqYiaBKEZ8IQCk2nBqtVV88Zn+If00V8h1DIy07d9MfIPu3c7W5KvkS3eVuBuZF0cmJUKvDz
pfzpUUoonN62A4B5BljjAlUK6fU/8LU9zZuaUVW2FRCh6YJgZut+9lje69N3Unk9YCk7BgKj6XIU
CDAqB4KjdYtErCvTNx5toR72LfOA6PqnkCX9cUPJb8In53dtpv9ejxr+x4mcz2MRBsH5e0fL2SMT
XY/GvWS5NtSlcgzdvsBesC8bVSfle2GpzHTEa4QRR2F/7xUOYul4cRHFM43aAgRR0XQZeZrJGJit
/XRQPPQdfyXjg+XUDs4lGLSaEpfhy71yX0sEYrJVr/XXCjo4nXwapgZQOC61XuNmtW8nz0tiqHos
ociCIaSOnr5cXQqkmxGg6p2SmBzCpsS4ElKkXKArhdiIgeIyN3z6KKI1GaZ8ZWpik22F5+9nr76y
qMfbOtdBGRdbK8uTbuMHjOO/x5u/Rt4VzkhY9re5FgTuGhcZH2XJ2OBySNIsGezVHGimWntWGycb
mhsOuK6Aptf7WL8k8+kERppmAh7DUFWPfifnWOo70X1amzRKIYk+GCoLlyzHybZRNvlKSiDG2dyA
RpWI2JbIpbOdnLikzR3310+nFoLih3KBpsBPYjgHj2jbrYh4JFgM0+mMiuyCS3Lsl0NCI0WWZmW7
bSx3VZg46vuPineG8lW+oyU6Pbqc1ohUrkudcV4fv1V7pAvj7QdBVA7F6+79+JDGfrNhRUzO24Br
8jLvT75vyGDBYcXwC4xNsFqbJxir78OHrIt2w+kFzTOMnb8wyKqK0C43oYsrF1ttjNAd+11be9kF
SsH0OnWBD1PVCyc2CMGe/waDPQZcqIFcd3KYuBo9Tf9zQAiLLbhEJWzSYC3Y9wux1bngh0iecrAO
9ahTHyWtCY2z6PFI2QQgWr+wzkE7hIFW25kerevPVBYBshuHQQpvlfns2gTZCHL9907MMzkKsMUr
kg6HGZoQCNUMlamdCLYisXqyiz7NvunVsyivr0+ld+KUzZC/xP26EATdhqSIq1PjZAgRC8yPOLEj
8ivb5qG7Cog6G+GXknXfTsNNYfr1iSCo1yC0N36TYUFln25lm1AhVdEzzMluM82gkszFYVeTJ6eu
XckY9F+xLIRAvuZEpqKFnSy763cxf1wuWBdadQJXppebWeHg5s10n60BPeocEzgAw/O6SvlxPJMS
qgailALFht0eFj6HN2Z+E43alkB6tSa1H5JUhGkzl1/NcVn8a8OdRHN7at1F2ZKQZzDXKEZ3kGnx
/IO16ivmFr3QjVxXPsbqlONOz/36x84wzlHG7v/yqT3I7DppmIRzUU/DqQWMBCHkvJeaJqmydacp
r2mOTrVRt4JzEkFIPpki03oqcRdFUP6MyqJI4ETsBMn27Q/pRKDV5gUvlZ7f1bd0sMFxTe8Gjqgw
smYMR2YEGXlxdD2dsQuczgrHNmSR5NhdxODd6GmEWy4CCbcFTgZeW2Mj6WVCeP/ZvJloia79/oE1
xfixOEErLtcIJCZxm7WqmNttat/RJErPBOUDyMU23bQvbFhU83WBBXcjQcZ2wWVkncoVfC34vt2w
tW+vRQtVnM76JC7iqSR1UZcZBdYcE7BCTcO44fjvgjSjDS4AlkCkP2vXWchRLhlf5ntJf/M67WTw
eqQFQfd9D2m8eR/y5u1P8q/AQa/pAXUsIIo8FL0RWSZ50V+mY+r63SZ8yQYhG30m/6ojeAA9aUyp
byvc50GUOvWr2kdWNV2SWZbLZiX0EZE3+kwJmiZH7ZVPZ2ilCDC+tSTRzIS+iYJWkU1acG3GcDkP
bPpw4KkT8BkE88vcxnmhhZAmtaP9XDcifDwf0oGHPOy18tMBx5KyQiTsFOwRlj0m8VJmqcXFsL0G
2HXvzPUOPTIoQKuCpalNKlfmY0V7TuHe5GZhHzq4h5CuJMeze7G2wD8ujKMd4LEbIrcGi3r0k6z8
BbhtQHoPCfZJvrbAMvUkESmlJZ02teS+5AxN6kQQOq9yUsnvwBRcxQtBJ3M0r/SiyUlla7HJ8K1+
3s0dG9nhjlQ++X6iQ/aaYUCg5zJ84i2IKifGkbGthxiPROpQur/8OJiKdsY2CCOOaQi4tKtTy2fn
zUxNim4bjAKGeUElxQl6wJqbgwSsMnFmhLvCKtdJwH5ZGhPeS4ut/KdvcbzEKwphwpFNbUYIJxXz
DeaiWEF4BvoPzfVpxbpnZJQkjJ2wy857detGfkq6+pWIxOe8TTMjBQno6Tn3sT8qm5G6dkfQsK2o
4x+HBIk/3faygTuUEV1HTy/hOEvY2vZEQV/Ztr+c6Ch5NlNRglYgJYXMSkSYkiTOjT4RdDnxh5zo
yE2w+AalOcDp5ZVQANGkZPulVIIkU/+7aTJiCIvL32EQwGuxJi1oLKfw78SmSDtWBts1Z1G4499E
VzcisQo4ubUtbwRb2PLIvBQAkkKxjbfXiHhtyEhB9cSkmGYeDOYHezrhxiYiAao4hLFIzeYIHrQb
LXG2BHKNjE6aFEd9ZY90s5O8kcVHFK/TUqt9XdxDgGtkh3B2ylXd+lkl4OcBzjc20pwVYR2FmEpi
W605RAkFKkAzwesu9qPEqASX27IR8aALelGn7IdGjBum/F2n3pxalY3YrS1KkI+KcW+9nc4CE1mI
s/QYHTK38qiRvdmt1iP9gfo7+l9KZweGjtHY98+TKeKljHhawTry140s8v68Fno1QuHAvQJlC09Q
lRLqoFW1bRvkQl+3RnO/1cZtzbxh0mbdsHpdSarqNT8dVK0wkiMQTdp9FuRjITMZrhvHB863Zd+3
wublO7H8p3TSxtLqssBs9rGVxN+nCbBfpdhpaMinVfbiWyIhyRe1Le+vKxjxWpF2Hu0YObafW7UA
IC+MAdnnn8EUHG1oBL23Y52Pkm96YDyL5Jhc8jodsCQK+EqEiHhsnCaCHNByiE4GhTCksMv4t7wT
ZgLA2Tj379uJUsKM3uteXeviudW2QEm21pxm7TzNpneAG0ECNlCvUN2J2+AI/ocQABP47UH09LTP
URIYdDV0lOcvuG8wYRpHexajLnaIbkGUemWvY/Ga4Xei5UnD19UzFFvnDg10Q8/dHY8eF773Wf2d
DNVchlkLdrw9tfvRMSHdmJo8i0zopWFR+kkB0q4w4717W73r3emOlqGtIaR23Q2tjOIdWzAK/jeh
mi4Fe7UPwbGgmW0G79g1QAgBXDOxrh6rLWB50iE7PrJY9sABA3UNRIjGcwRqIRHUgccqRxKcfCUS
N1w1OEiFbozFlvu76FIowLDmjAtXZw4jyxecyjKlyGu+OjFMFn4dQGHh0mpiz7CgwB2UwU/xeLQp
PvToJCPCRQXosqdnFlOX83F7kMPC0bg61eiaerZGuaSRLFZuVbrYapLtjWko/gxhZ1BvM+wwRUWF
jhjois940u5WW7wWioXV+wZr/Q3RiRjumJY9UpiALJ2UZtvUNSxk7x5ujeE4ZElVJMjshMXkMhJU
D1FFLmCAuiB4m4ZtgJhLP2u6JEY18IlRQ11Kr2vCd3VykVxZWIDWTuEDjpxT/4BTt+6HhufjS5z9
a6RKHxzjnb+63N6OOoUhapuzlDp5jBSSMHBT4b5Dbeylm4c7edcdUic25UReqPjk5Iwr/7PVUUgK
LCVokYD3iiYm+rvE0GDsBgHYfOP91th3RuWQV6PyLTKwgrKfIZu3iiI8MN8gxJX8b52DuVONGqwL
y79bJzb8XUHNbvWXnivrLF0GiL8dCNnRCadZAkwwNk6Yt+w5BbnYbZOv9N+sNmNqkyL+cN+yuJ3t
ntCRmssSsklpFeFo8/ylhKPOrrJg8StesozApU+MxbbXwsRnpvdgjL7hzsKwnUGwm8sEXWbIbSLc
gdz5UAyIF5NvM2ztTe99JPUCVTjB0MeLMxN5bLfqysWKQY3qbAVqs4qBAcxAFNgtCybldpUD7yrI
1067bk7P1Qkt1TNHEBxln0t2GCnxU4q/X5pea2p7FmHGwV7srmJSSPyb75AyTHMSzTIGhU6C2PI0
vVZejuSW5dJf2eSr2HbvzmB6r934UNaWuFSO6n+ijLH4aOVcjPU3IgzPE5gm6+AJaExaLVF1TLMD
n8nD5sB1S22BieKWvWnfEuQ5HUE/bvU6j6T2IjCnAUVg1PBAfLuEppofKHBjzWhvil5p3AUHvzrm
i9CPGx4l1W9vWD6AR7GK/VqU0Dt9bZadYhxUnCsBoln5vDKZ6ICK4AAjceNcRcxj421Qbnn01yQG
9/tGc9LyTrg2jL1EGmTvgvkiNVrp9wUSayawv39xFMY7Xr6oFibx7CncWjTcansQq/x0fw20sOq5
sXlAPxAEMEIEIEdf6lSX4vdxe/tyO3gk6wepNIGOv6Lt4zb5jiWUQv6fFNEjEsna8Y2LFDxZAZJu
Xcj7RHk6GzTZpzoSuQQvxnjXlWrN4bixKIke7u6XF1vcN+coY6HYrn6sgPWp/fyqOEoAgirtP97r
F/iJC3hIM7uK0mn7EldJKXS+SeXiXYa7NjgIq8cmlcX8U3L73CuUE+LVkvoLgCBB7nXgPjgx5VmG
lnrQJBMFoGOlqRKteIJcy7y3cCxBOn2ZObvqSTYdJwexTv4zFX8iqdoyoFg5cIjMaEJriCQa0j7n
mmH77h2n3COAqiQtugVk68qD2jpRkK1WGQPJFMXG8P7o+t7U9jqjvYyT6E6QAAXoG42+C+6L4svu
gdm4x18ZVI6VnhmuO80QITn9AvF5WmfCseXyHMzzu/DG1rsMdy+ghnsdO952Lb5t6TAVrWb6oyJD
VLtIPPyQtQHsawiddbxmGm9LvX33HVBEBWlKlkqyPkfat8w3MW79/pMaHX7x13JXgWgOx+xXOXkN
E8FSsUGIclUeHMUNfrSj/PYwFEISzpJLUmr/+xfcWY1DfyUwap0XZKx1gaOzbdr/ikEXSGw4UJzt
U06pPIm8M+BganT4SaYkEGKMmI56IebHbAAbp/VfHFxqFGSpHNBk1ZzmEr65ZhQQ5RQy4BCfqj0x
WiZH4Ds8kt4lhbVlZ1jduZma8f2uG7Fv0cjmdAy3dBjvEpjqPixQzUwSHvNecJDE2TOpKhOF7bXu
smdWmU0h8VMq7eEdU+1oCpPIR2dypYbkkdFj0hKvz2B6EiZYF/vqKvxSWUkYTEaYdjX5gm/KhpWT
D999wKFyJsBrgeFt8DkJxiL4iSsv0kwmZOE9i9ZQ/x0/bqkr4IuQw5cyQeFJGJcd2wg+dDoi4cSM
pgoxMFaGqoCma7pULv1Jv8wlp+WrKt6P9Rjroy9rZRQiNjZKEj+HTFMPIEvohPVcsZSFbXfmgZ+i
oHxntAoFL/C6BZxMuWabVXjyk5aaBulNHl1mVa+9Y49bOv2ndgMLy5T3nfCouZlFQOfMTZYRcNkh
2JdhFGeWCzqUOOJkd1MBe6+kpRSeyiEN/inUcJ+xRlRU9YkepoA13qzG8Oe/1+6RAsHDk9AruiL5
l7rA4T4yy4YojyLqgewTLzEAJVGULy95+2GKca4Ij9WQCzKJc8Ya3kt+w3FVEDGrYEXppTSP1wKb
UdU091erZxncJvQ01JYYDIxgMtqfuu97m8Ie3eJhYlNhrAIl3jdibsEYmLgy6vf9AOUU6UOcmcP+
n0DI6i2HotQC6YZSA6/k2XrgL8zOYl4ZIUny0NADq8xhhizLhj1BiLp5Oq6y8i1/RZOeuu0OTgPi
yydqoI/L3cFnfewl2wPoo4BzliLWRBJ2nwpqXoGA3iHOHXpS5WzcSQwgKNHmHnzP487O4osM67ou
11PRpSaYGiirvN3ca3YvWfnze+Mlo2TXt8Lqj1IIHII5Ou2PpC99XvUAYCzdJqyS3vVVyZmTi3jK
sQEv1HR4kTc3l/oFGNKUpGZc4IOld7oRL/622fcTSKnsCjMiy+xL21aWVpGUDsDlNk57rQmUItb0
nkZ4BIt7uvyxIvcokUG6EaW4bqW01th04JUDYM66I+MrEYkGSstFd2w7+Du44yiLjnH6wT/cXbUu
NejTf4BDwSQLaHiHLeoDLlZAryja+ehhLf+tGdTj01WajARIrWeGzBBb2fYGkcHfzcs51G78bow0
3J0rd/RNrkBS0kxYnpRhMI/HlzB7AjO7kIaUIfpMcQPkqBXmoosZheLMyLIuAgErvB1LQgIpVb2F
SzYyIwQFzslGNSDy7IOH7+4jZGdZpvx5RTZLNNWiOlNt7k0uZw5VyvSl8bLAfT13h42YbuH95BgS
RmigwKU8ft7RTriGHKSzvvBwfcs1gXQd0LaJq+wTGVSmD603/rPPgbeoWV52wLEPaNKFtBK8mphx
WvU3haKfRVrpJRq9uPIV2fWZFZb0O1u+IoxPDC3kFb9Mbas7viuDvCbDG8Ssx+cHXUvaDdpaLLYH
PrZCs0X6QWk3Zy96tBBiY1qsC3rCtmmLfUHn2dI+bm+f00onRU/NX2p6aQUQ7fZuh1SuZZwyFnrj
jL6KOrcGPxEmYWa/NhADxEfwL+djc8Zp5kOGgiFREreFj9FgkmTNO1cq6IpTvugECqtylMXfSTvV
epRbdj9vnG2Gcaxvq84eTl06yRZ5TUNYTMxczB6V4JT4aUZa0e50cmV1DpVuK4W8GhFQwLrjDbie
ph+NPBKX5gSllvBOYxXAPxSXmhJNJ2JAKnpmiQN9haq1RXMo0RtkErgUkyp27Jd3tKW2Ak+u9U22
fjMW6epvg58Zq8jUClxC8mV7Sd/5PxKlSU6Od++kBp6trVza+4FXpH9a/scU7rIXLiX2w6W23lOj
+hd4RVmYSZO0wRpCU4c0/XxeVx9O524He7DzIMEnxgGoEwRsolzOTmL7vC8KNpnV204z75vjy8bm
PzWTP/J7OKmTfbKTFfNHyR+HvgR/6Z9A0QX6kHhPJcW7H9mVUEdzkgKCjcTHAxhIUZkEAoWIRJmO
kxE9K9lODuaSSgBjOIG3len2fjxUYLBef8/Nyh8oTcs+Bmn5ACPy2oPp/oMV5T43ffqyq/e3UlKB
zOa3hB5XO8Ux3/QYSy+KtzwW175/IiCJAvf4VLxmxpZM4XGF795jo2qolFcmRbrlGomotp976Jcf
lmyw8w8RsX8h/+k1H1pyj88hUkKQuk7tmtxTN19BcAzsAC5aKKNNhYp/y8de6lFkviUSKY2+eQxP
RXGp7ltD/osui8sT/4V9VKWsA9Kgv5vMb/9SODmaQ0ALapIlEJ2kolskdySAW855BEEbQSb1P84r
2HpiYE4DPJlmKHXOXYVADlWy54xpAe42juPrLAAcJAUlcNf/MAfRg+3Ry2OJB8IqipXTyNs4H/92
geJk1M5REEkuojNHjrOFX3ZnMuqlbm5jIYdZOK9GgmHv1HfHKIMQlJmtRo1HEQvTVYekeZLdsZEd
8UCp9g6SvVjoTjbzvG3Mza7iIGLC2xHcKCuvIiiB6oKio++dozUpdo+H/f8ff1aKTWErfq+8cE96
k9ZlWUZN7v3WmyxOggZLahSqJ4dnNRYfjaFuSL2Hk6g75vsl1YHRQ1weKJ4q7PRv7hvJLryyX+nm
+I+Gp/Lu3/zzqdvAQVI8DNLzkG19rGlA0eNq5i20MBxLPLAg8EiSqhJJdfieuSamnX2uxVXwHa5y
+BLYEguGKYljYI7i2aVjVhYBL/uSczGzDB6nPmeW1tHbXDTZycZw8iUXyg5Pi1cW+m4jUzvSV2er
Xt5MzLnRQo84FR02VBDblzPtWn5yYn3ayypInWZzBSWWdgXbCituQVuKRq4RfZnDK2IQK7/GMrXB
roS1ubmFomFrYuTtsgYe8Xd6KixHenr4ctuynbF9tbDAaN48TCjqfEs3r7B+dNn7yz2Yx0brefT6
igBZmwYZnXN+3MWSab9gzEZrcBeW6YghDe0+IlI8Q858X/IqDGYje6wQOxvPTTOfNAptqeDbOSeC
wpuS8uyUwgrDIqfydX2lP5NEB9lhT/zZl/MUWU+wtUmbo335mW/swUK8TnjaExHLr92YezEGPRS2
cXK3zbzCZKTNJYKKt8wqn/0vAOvRe/P3mQpwMySOrzmmUr4TwZm2O2OtNMT+3+Q0FEVs5jlSjX06
IJ662Y0ekaK0szjJuqU+0OMh6ddVUkwelgZIU+LAwBO0IEMG/8z3hVp3Mv+NJ4h61RWRR9+oICOx
hi0Zzkywh6QZxkN4MnQEjWIazNjNGoP7f5kFpyYDwelNnnegY6LQ7cBYu/NZTUYzMC7kt7fKnGtU
AfLpwTJ2LtCnNSMA1x6QqqQsmUPGgdKFYQVkiAs0aD9Oaeb8TSvTr2F7mfmAuE0h8NZ6CwhwiVg+
UFiKKq6Rl5CY9uJkIYAuAjsM+Ltv28XUuq4mG3PnI6T6ag5dW8iis6CoKv/vdvnn6tWlkWGFw4Ky
Ytc23u58dltCgxACUSDvR49TngpU0SxqBDx1Cq0hOjn28gcVz3pB4xB0A0bt2PfjpRgp21HyvEhY
SCmeIFjKW2WgSxk4ejUd59PNGm4kFVZm/0I7ozWAlYNXwW9pIWcpscajtRQ84anPp3Za/tj/mTBE
YuSZUuZIvi5Y8AiKq+Jiqbj/TjJmGYgmcHGda+M+e0J9EAIO0RfkotQl6SJEHqM5jKjvqvaDn/Z5
N7PM7zUgE1u9J9MDpZyaSL1VqD89gDlHkeu3MY7+QOZsXVY6WAKMDTs3flXxNXEjQKY3ioJbzmmy
Set4fxmz2crb9jTJlzdGG4Q9Jsm3cyg4JfrflsN9fx0K9dvnHdiKko9OgUAEqfDJAn2TFY4xGutC
nvI2jMWsr5VoO5tY63SFTDZ5TWx+709E8axMAbN5e/488bJuOMtjXtHxTA8Geqx5LJcp4kchG8OF
GDhLDp64wOYbfb1gCUy5fW8yQvtn0CR1njhxm5Zm4U8v8z3XEYVwtDBAfYX1q/1Hww+qx7MlCRgU
ft37bDKAHhcC914fb+R38FREiaVmZnWxg951Re3bDpKsGAu7v278XhrKCgX2tvY1d48HfQNf8zDn
et6xoLeulKMtCAt+itqfHX6Jzkot8CMUTnnqewuFROH22qJvBZxrg1Ik/UNkciEjK2Zegk5JVpqd
M0KxqJeoGeIRlQLG7kHqNGEiLbOrUXAMSS9bWGxYpffP5PKcYLEuOQFFou4n7/jag7etWGBm6cdx
/96N6MxXjK7xhVXd0vXSAhfOcfqtR3hBnIvD3MFFkKvzDp0KX/dkSL0sqaoy1rZ6HUlRVzfkwWoC
OERvZN29NR53zWvpwLMLnVhG06WX4U9K3M4pmXSeE+aDu3YepjyOVV8Pxz62Euv49Cy1Mlg3dlvj
Cqf/XgaJn8m5IHSkC9GpiSCPBw3XwdkKr9TPOz1Cf9cIHKGcNBFrWL33AEizFHorFeKUy0I0t4Zc
JScc3tvCt78vIU1b6l5a6grlexs1gM4H+EsEVPupQfZ5SotldAJiSk7hcgCGl2y7oOffxLBd8oHz
wQgXqmHyQyAR6QB/ZYfH3e6vOae2TfZkcwBQ9g2a0hgoCTI0Y3D8n3f3F23hIQ784LfHWCmh8nxE
kfDuYic8pVyvFdqqQo/rKzLHuP95CxOjNRNKPAj8kjima1Gbj3J51ZZybFVOGLZN0OWHK7i9WRsb
PTQupXsNmyBRMSyoLN36czjbyJYSeb/D0JaEHGBt94rj0lZ0DnHNPtaJJdsaVc9uNxFs/BhqWHLf
j5AZSEKAMbrG6tw1GYExNhj7onJHn/jAC0BLgOaEeIrKLRdN/By5k15wppYw9t4JfXonpQaQHNVR
0XLlAHMdquvfMLxHpz0lQM+/88QbD8m2QN2lHEm2fR0mPkyfLInmQPfduSeAXhu4eR/934estux0
q2JMxnjanHwrdy7z7Uhe5dRTTek+HweT339kcynboJEDLfSVLXFv9erH7l/FiwijpthKAbNSPUhN
19TOymwLNt2Oqu16lTrHsKVSa5m/QHBD82sPM6Hymp6A/jJZa5vIPSLCzygLkIWA0/D/r4mopOv+
4yvUgJzb3jWdzVZRTALNGojKcT5kNF9zhVnx0NE5lyHFaNPUjQ8velO8E/I22/LLo1txzHKyskA8
IggZcqk2QBZ3sdjflqX/1tA1KQqmtEi8NGR650QAE2hc4oZzO+maHXZxlidK5EUgEtiuPYp9Wz8X
fBRnMwmb3B0Jf/l69jBn/NlehiM3VGGdTLps6sdPLAJf8jDImTX5bO/+MhJtyUka70b7AeNOygkQ
buS+SCB3SoYEgEyvswxj66XzUZU1o/Gc6dRr9krIV2NtS1nM+ArzMuNd02QnP2ZX/acmmYI8Wezm
1w1Mi5FBkw5CKUJBZqT+kyB68VX13vJ1g08lrxa+BOrLToneGMefI89vsEloJBZmiWMc9R7Ihj/h
QZ57U/tuU+oKQpSgk0kTtJb8DslmmUURjfa2MtWOGmykMCcj4inCpXl0U+dmTm8eb2+s6fWVIO4W
o1x9p8lzoz7e0rmRxwlB9Txiv4Ykfu25rLtKq06+0EshecSE7FK/24z9jkoKaXmRpaWuGTlPwjQK
sP98LzLB+MHdjumn8edUD4d46OR6jOhk+nxIH8A9vOUBhJYRgDjXxjOj8fiTza1TQEO4e0tL9yjH
60iwbSHWWLoWwHk5T5CYKF+ZSDUczspVnXpcljCyMRm7b8G9mMWD5GtkQ4W6zpC5XQGkteZGQ/wI
C/ZBa7DmNDBjVOUQxpTFPBmVZp8wfe1Xrne8grkVXMOsYwf8R0wQTQzPLk78KI7Um2BP0rTvd7qf
luKMdvaYByEJCDzZR8Cym0b8IRE2hbqt4m/Y5ivHV45M1incdOvPQcBsSS4cW8IY1MXLmzjsJdtE
k3X1pnRogI6gv8mpRbMA17cczenRuSd+Ulr19Nj/USSHEw40kWhNFfUkZNe2nLRDSw2j8TpJA4Qr
h2AymkA6XuvXOJhyZlS8SllWMCKPxZDiipKgnmMxMqHHFOT3J7eBBBjI39AUHSyWGQYtv/PFGbCx
sl4kFRN/CTb2lwH9mxogDMO1sluMFnrK9Rz3IMN5TRm9sZR6qRRa2Y7Ajlwy+HKpsndsf8trku5E
VZE0NL88hjriSitMTDTWVsI0tRhgSu+T/RC/LOo87RohJt5T4Bs8IN2kFwUbteLBf20ya6JWPlwI
HLYKHshtCICE6y2JfpF9/LDY5W3VEE6F0rAYu1jvSstn4aO7qeG3TfD2UJl9IPXO217dsg/iMg7X
J5BTB8PRS1O/uag1cmAZ1yr/xxS7V0y3vTG3FZCS05lBctB5cTBNUmv23Nfa+1gQ9MqXrEM0sVoZ
N1zwArT05MIUiTBulFNc3nR6XKbRISTCdds2fAK2z2SfKL7GUS3YO00pQ8spqujQAFYxivKfAb6p
w7huvIMeNMpZbZZicX9hjZJk/uaqFG6H9/57SxH4P3F2SZF9lUSkZNlbAueKyQT/wLu8YstU+/qK
kK11ro6bGOeZvPON9gh+IAtXhofQfVIFfzlehMBJOfMPAWbqNPuk4/x7y9voJadzJ2A317WLWYBl
SqQbixfFHSdyXx+7Ggs9zkFRRrrirv3p7tJGthcrAVp+NVLJqdedXLaH4xZiIR3rmG1cGA2sP9Zq
mly/va5TsnZwocAyQ+1P6bVKbW11+yJ+hR78McyB6XiBOsgUWiiD9lk5SXD2fD0812ey4HTWUs9Y
y5DEESCaS6yPceZO4Jv1qNE7UJfB4S6HNC0Kp5EOKHvi/nyPbzRQ5Mz7eF4LyDDyQHCrXJRjLirh
7U/eiAQXOJStc0aaMttk+jK5Z+O0g+xhhgWFJ0vPXapI1vQ3OeoihfdsHnQxe+L6kh3aVNih+oEk
3O/f9EsoMaAkNzxuXGciQlQIhTvF+2gYzMOLVgnZ46VXjJ6k7gAFvKouVp5vPXGmElN+PW5gpWAM
rLyF+tAPfXdxizsEd43CTQvFWLLtxbQCLfUTh0VNQda0JZLxpZ/dPEmAgfyNmBlEfFkNBdbrJf/E
FpYc8nCXHEVcXyWdUtBsRT+eiC15vtgZK39dT+v3ib/F5K82Zxzk+xVOVkk7AleIT0c8mcsXndDk
Fe/EWENfvHKzp2NTFRR700itnBtgAREzJ10KtqHjZkG4i3HBw51lp9oRaf8OygTn/M2BlqAYhnBf
/EhVuhXin3F39R2RwlYqgFhmJ34b539nSCmZ/e6aq1cjYuM0/GkE1QKku/D6zYwuorw+QauHCjS0
YpodYad0B/xKF+QfvmuwpoWv8R7Vw2UH01url0BF02hhn9knSsx/X0zh+LvB31aby0mgT6CWW3gy
BKSU3PKKIzyk6lgk2OukLfwc2GgyH4ChvZzLuw4fgX8iWmUi+R1ZPFI6WEoY4sRYxLdapSLLCZFi
82pyYPl4lf9WTyp70jc0B6zxmQ2ewa4/q1a2vmu6Rv+4YJu3yGyhY5fnfxkmJi6hsWc3kRHUekFe
SuR5KP9PZ+fDJZul6TWMmjH0cuaGoW41E1LqYNPNbLH/b8jYPJk0HM/4GarhtxPG9UxWu4K2pFln
m6O/KJz5NnXFDPdp7TzNlqySwfrjjTV0iupfgvu+izpGFjo4/WpgRTRsdDO9KLsXDrO8VTpuewif
WEuroTKrVMDiMEug+rNUW4Qv9EJqeYNrtnjcrxutEKcX6n+BC/qoCsJEzwjArd/k/kSo7lnJdIhf
NsWMdzl2eX9KeNs8c47hygmTb3qUWnUkDDUlDWBR7Z9WFX6Yh6wx4BTRYRAOwY1FffiS3qJjCSJO
Te7NOPo03K6up6+ulipehddSHDnginI+GhHuuz4SEhNBmcVuqzVeM2MtzlOEgHotKPSTBDXnq4gf
3Fg8mhmRjkTqOE/UVumWSbpduecOhOD2Ii7N+rm5EKbZg9Uiwxfet1ZB6dFzNmJQ2kojvmVhOx4k
AQxpJgSpxmVOF+ZzR7i8/pIQimK8MXcdBg4REYJc7va962dUD3gQ1S2MQbc9VulSW0nOSyzkw4D5
1+E5GXmOKGH8GBgRjLpamtKIgEkUy230HZV1/C2jR3OCf+daAZuduTdeFsbr+MlPrV/wlVxDphq2
gZfy8fq72TR484hhzO5IyF8znOrwm3ArsGnomY93Qiz5THOfXuncUnF86i5EmYegHD7xtnRSiVuJ
Ki85SB37FmGRbzqvzTxD+CAV8BTSvYq7BotnOHMAE2RX5epzPxc3l3AWiQL8b2ZOkx+NW2dbyAYG
BAzVYl87JFXgPNT6R5VmxFL481v9BjcoeEJitwUIgsJPOQVcM/9pHPlTYZPw2BbcGYGfGLQVjzEU
9q6UTEpSvvY+ZuIYKsnDKLfR1B7ISdWOT3ltj2/Co4mzUCGZcWfydQ+8x3L1gTGs3hKhA6UMcmKI
9tMmL5uD/VbJpeQykaR8nscPBfppiwpHZRviQu3qepG8atkSGRZM40iPHAIJQXRGasqtoAz4Xx8e
X3SGCfHJbvCmQt17JXWh2bBuADdARebLyhC5T3KmZcukK1F0NJirwhC6h22HWhidwNnQNrWKaNqr
TgsqwMLu00LaFMcy/KXprVF+AGZa700aZPYnc7mK13soWHUXTusKvlFtAAGjAWa5L8D1EMpSHNn3
2LuIun+T8x7PRlIDT6q5TOOxbtYRMtPMSUlZb5L9kbgrZDWPia73nIFLHqsUIM6SRgFH9LjCOnk+
LhlpcOd9cNgxCQ07xp9hDo5MybW3HD18DwhaSLrTk9U/DHdsQsewua4QsyjBP74bA7clMviIf2tG
Q42z7cAbqLKKzqTOXobVsNmhmsfIBuDivRHtDeRyFaHpNOr2paLCnrlvhHgcFP7/qY76F+wpoMX7
dj7VY/iH93EGASCZHIfjqdo5PbSX2IpEihPQFKACW8GmWKELmMBT1HjnNcj2/vYsg0XnCfdDLNpk
HR0CyMLUW/CNLENJVVdK6Or+amhRtQ21xhc7x2YjzVjLBqBlG/xr6c2zynMAWTGTI/FcUZZRQ0Qd
CPQyYDuOYlbTQwGdE1kMgo7MPZ4p85D2fuPISp5zfQpFCsLPLINnSRQdAkAL1B/4VNrGDi7bdpb1
Hq0VRDDzEXiN7UVLcH+sWrU0fDDv1kPxsSMMxAZsYsNb3fSKEj2lysq9YE5xY8jQfB2Ea3GyQhdj
Ii/AsygU2PNAN80Jh4ZL2cDGMeLqtsW3mnAOXFO44phlugo9Ir2XG5reQmr73sn+Mdsu2iYANLjR
jt+1ZaoMCj7XcbXeSEb1Q9Al2QxXP6hjFlwAxNoLqHvSLuZ/58TQAkdmMJSGvh2x3d8gwML1xDrT
DS4Y+GhwtVE3/snaM6hWAmoc5gySpWFyehYMKo+v9F6zbeLy3InmtqK88yQJXkU5SHo7Jeg9R8sc
bQEQ2H2OsMpFz2svtqe1C/TowZC9yBeu1My6Z9c4GBYXNe9jhBepmsUGpeJEQtqdg+63GJgajgGV
khO85n+mbfbDTZA22aVbv/8etIZV0iOnUVg77h+xEk/36BaPgJ9FXyl3XohmE2gL5SNv17jyJHGo
MRDSfAur0Aur3j73gKdom54zJd8INyR4EPwWz8RKA5wWcNyNZwtounInCEv2NeUJ25Pmaj2t0QMq
cFVODPITF7ZNE0IpcNdKWysMSGLMBfaq/iCbNgQu0m5H00XfxvuKkhanOkosesHeGwHhWcaH1/vJ
mx1RVGGs8Bf4c+Hxvw9/QTFDzhIav3h2nRyRirkkwLuXgMeDD6b1JTvB7lKgRfPJveXoDihUWAF5
YBs986EesUQkv7Wu12cnXW1LZU7wCNj+Gc1xP3bTUboRWW6itmZAqkTjJzpJCOFk3JHcVsHwKnuj
Juj0uNhyIcui02l7d1XTZ7E9eZu8lk2AQAWtVUXS2KsNrW7G8DPWvR0Ob41+C6MPlguizlXL92zd
CRUwW0bIwE+CCVqx5tPVIzzUQu0hAZ1CwwVUSdTGoTw+JjG5gXeggroz4aFDgdb20egt+edPnZNl
NiTCQ065evpEe3M9BdM6ndH61sI5peUpYygLUx3Vu6no3SgmtrMpk1o9va7g8RGvVZETG+7y8wQj
PqRhWNi8MqBsAjWz+4BYXIY1S0CMiUuC2msVSPG/nAwskujCnOBhoTjZiEX/A3eQSSfGhYM5jWnM
qHhK/e4JqdVW9DDgqSDh5Dij1SkDvexJnQLKqJ4bqwLfd9yDxVslxkbVhAyGNiGmRaLm70GOBzV4
e2Yc52GyzIAMgVJ44Opbow57N7TGPJFapqgkcOBIJvWKtTViTnK5CPxw4oJDCbiY/K25oNMoqQMD
n6BRFt4a4/MJae2mplJUWlyJ7Hp7rCxs6Tg7N2ZY50CTfzou7vod9vnLoPH6dhVyuvL8bzCP8jK/
uhdJ6p7GExN92OEb5DRMukO7oFz/bxsFNefLfTwuaOxtkdCilrIEln7j/Wv++5l3dnMVNV68mzNj
1QgDZ/RWWes+FaBGVnUoWSnnNfcGduATrwD/RxX2Pd+dCOfHDtFrwH6l1vG3pRuZMXpLZfteumFg
lqp4ZKGsxGJxW1z8VBd3C5uN8Cdo2KXpcqcT9NsAXgZldZ4aFlcx6E4Lz/ddvfp0UZG+Dz/Tl+oy
HBMlZPEWraKOag/vluwTEVKyrBPN3uMgiYX61itamPFqDDb9Ukombm/mEP0B7G81xGexhRe285Lc
iD0B4qT+y1DE5U+Q+7W5tjzqx2FkF//RczS5RZDlC+NCpd4P/IfW1DTuP6/0X8qx+rn29LkEvC8O
FgBXUH9r5ypMnHwWJ3fvef88OCbgShQZHmdBNkKmlCG9pXQW+0F4pARsz0gK2y5sFlp3Yco4m/nO
Yv7rk2ZuZcvU4JiaxoddyuyweZyaphlE2TCaYX16GRcQuZp4/h90xVf+5MgYY73JYGNV7qk2Vhpr
3zJEIIlvbc7AGsa0G7Op2dlD0vMiL/l1Z+8wH72LZpWz+MxoZh9ZiQZCvoXtp7XlcpSacohPCpBr
pdFFEYC+4iDrHb8Uy0vmewxn0CqEKQUUN6i+oZs/Mpcwv6ilXiXCst9plgIA3RJqUjtcuolhicqM
6wJOTprHg1j6z6DtSgx95HaHhzzTQHSgOG94MjhdP0Jui7yCZLIIyfH3Rm/4cVnK3ef2Fyi5e9b5
kwVDACkdFw9Y1OuPJU3tUIvCHrWQtYLUfAm/dxWcQWzJYCaT0GaxmOy/4rWcONj95sN/LHK4omYA
6Byv+L7XTFeJMGVQENNqBxfAynzEPItNqACXxpFbqS8CYOBzQAMoWaBVSdqJ4lMkcWEk0wpeVcX5
C0KzKrAsC/xmQUClwtd8ENZ5pt2HjMI/Iq+Yq71H72mfNssEFIJfPTMnvyJSR+ZXL29pCzvTc9rj
ErLQO8hHEk3tO682njb9nXHhMVvfo05jkJ50zDnLT7A7CNue19V6Gzc3BziJywsIprSPisFpBznD
Cd4HrMr/CW0qWkglW5X8D82oV7hF7oDqji79SKc+LmU2cN3lcPDYLXS3kF6orqB65hd/3b8GIJ91
i1a9+7VRuo2aYUmMqQLShk/OjfQTwlizcWyQU33MV3roykCygWmlQ0s4WEM5gahJvhvASGiwKR2p
8cn3hReL+8boTrrsaC92OiJtwJnG1oX+1y6X4MBwcA04n9Vfz8TkGWA+qGBGSTR+VWRRWpyivgEl
K7MCUony31C9P8Cg4qVvTQB6Sp3zrniUUExPqzBkQRBA15ffAgJ2sv8QxWIewWsaRmi1CGMr0aF/
T4uXJQY0Qg0Gx6OZjyFZhCG6Bq6uXXoujmthCCCFu/Z91le2G6LWH2syXu5igfVi9Wha7alu5RVK
8JTvVqRoIaLsrwwIkKUuxnaW9XsCo0ORReBuRLxuzvmU5Bpa+OhFnW01fsGUDnIm3TRmgdEzOTDr
9VzwyE6vrpwwzSyS5Vn3bVpPkM3oiT1iADbdgGKM1etBJJv3NN9rVv0yGkmoF3y+dkU8EV/X4GFo
LryymP0iKSaXY+/J7HboHG/MRsK2mIxVcbA7ZYSontPNVUP0WwCu+tscc+RqzD5JPurmn2YZ24ay
IGnDznszAwziG4QFlJ+QmNo/q8zGgTnBiw5nelKJxyi9McB9/S14Uz14TODhGVW9hM7XlFdyMRSS
1xv7Z+PqslwP9XNkA6HBBhnthMRC3gsIx9NV+pJI7TcX4rqcnUXfvkzo9kTUe4leRZsiSh5ZP29N
mLrT7yQW8Apb1Hc5xbLmq+Y8z3O2KUt4ieA1HIsazks1Wb0yfdxXjgdEjc5d64+qKDbcyu3APn3+
xuh3WCuJ+8VfVoMEE0Qe8AgEYRiPhepXgkvV55J1K1b4iOY8ScSqJBQjnZZzW2KuaOzCmsi7/CAg
ZLyz5WZstvroS2m4v3RPBNU9xbFlHACAnqjysOs3CIWEcMX3HWUKY9E+w2RM2D3N1Tpkrp3wanyt
8FzpFbIhGhnRvQTnUFyoE1B0wwtQNk9E4wYUR+JzLJ2A10fz22e1w35FkHqne8GPVaV/C3MhPKNc
9Mtu2g9nN7BLuPwRz0srpdibsONynl69IDdkGRb2wOb4FaG/BYhp9tjQ75M2d5TYdM3eT4TtDCJW
X+7th2gNQeOR5IfQL4sPdngRpZoG1Z/VcLwJfCItwSNV8sF7nOIHaZColYt6tD8S+4ZtY/bSCcE8
/vq7BjATgF7Z5bPWp68rWWMhlhLE8nCqdNm3hIY0zSHy0a4OQGG0cM+4yOfMm4LndR60mityXTC9
gdsjhe8Eh3F3nC2PzG+GiT5P7WDGOVv0vTczxyv/3zYB1nnf9XJCY6HCy4ng1D8Bp3l2mlMz0Q/T
/jJoRVnM9M4eALNKhmuRTTXWUUU5OwZyP9AdjrfYmZy9oMFUBAAbMIFwvg+qgUhlsvPWlxt+bj4v
rWIao1KKbwsq/MYgSKZ7HwZHnu4JVxQ2dQlxYmZRlBAmDi9fP0RfKa4/RuqY5SgA9nkOAVTWUoxX
H7cdUHc+2JaIAOgNgInbHxCeMliTE9lQ5VBKzqBWo7UVfIZqlA+ciBMEy60m1+m9DtNjwFPadjML
PHCRl/iMaykgA6aDrCEz/Yg/10n+v+kidEBpwml2SkTI3R4TrDKtjiFquiJMAdhorbyc1CSfbg8W
lEOu2RstL0H20rPYD4Nn1TXj2QtcD7jKvRwkMgnvgCLGXwGLCgF9V+ygI7jyHT5x4IJDKGrgtfkB
oVKRzU6LC9FNJQfHKvSO54IGa1l5t1kdatClmFBcDTJqy95L1h+YWMS+/1xIhE+kvQStVr7tB6lZ
7Vo0Jvn9e8Ag/FoxZDso3GQHEvwDoBMUahTOnGMExr0W65E8ifyXzkmy/J8sy+epszArEqZOTTW9
YGa2LY08EQjWOK2INSqGwyTQlsntVWCDi+FebXCiIGYibQ8D8qPTb4Z0ESLh/hPwfOjkh/ZdGPtG
OpOYXmCYVWglPBl/GxiTwcZR/MAAVX6XqQrj8weSkJY3Hk1g2JNTqoXfiYmWaRPLExwcgvKQm8vr
R1omONEzaqVoWkTXW8HsAKKcCjmnbzr2WRxerPxaMNq/9NBEbZtqoe6qCmUfFfdNGb6Lutv/VOH3
FB2gIAPiM2cwdD6ji0sIhcCzh9B0i8/fnURC6UdRSPwZoLivO5Rnxe+Bcu17vug/kXbvEx/IaP94
Hb9EknSZ9nw2+0J9XEiK5pWuFYGnwX9FNyY3/N4KJ5OV7Vk34F66D9TBA5HEWq1WCN2J63v1cFMN
Wf9OZgz5p9eR/2aRSXef6F89TOIdQuPtzewN7NaTEdRHMYbPKgcotadmcP6JH//AhkzS3B/vR4Jd
U2+PRsCiB3Q0YH18MzOyzuvbaruSfKhww6aCCzqwDwwjzCVvy8s0Hqd5lWN1FwxC+yE/t30DnzdO
7SS+hc5bgdj7n5Ia0BQGgdLgI/ihdxihtszT0XxmL7e2b5iNhGTlgbki90GmgQIyD7YLf87v4IvW
Yp/1YHMP9Wldrvq5VLBzvayrfrR7fJFZJcjkUXDx7FGqHTND0ir+sTpTyfaNvNRMe2C+ixeFc30q
C7czICbW7YfjpXUofna2UShMP2/HS8Qf5OcgXS4IJsVaT4YG/iB2k3UweLoLfhqzDdCT6yDKxzib
UN79GAdsmCC9f270irsw9WfE6YwGIEvSIiJUHOS+CJfioQaqiaOpzojnLOuN1vtiUwbUeGeWKRhF
WH71jZ30yw0buv2DPieFYoxjEuLpowOtfyc357mK0/LUaPBsA81INxiaweHyHqyvjeMN/586un/v
s9/Q02g828nGTQhKttm91uFwRjIGgR2T530LDcaUQrTGP8deud5WsbqP19KiNbdlj6RZJBszTdT9
x2Ie+y2xKgTWaP+LIJHGZOx0/fn3QU1XC+vG0NHMUWF5863SFekXhOnmo53cbq5BRCEvSZ7JcHj3
/o7+ACode7aOldaUbfENcy4eeXPQlggRYnwxgSy7jYOc1N7+UPGCxAKNX3ZVPDVgZgfdbKAh3JUS
K3XBnsl8ainMj2HgxrbD1UuuYNO4bb/m7bMRuLf23v+ImkYscjmbgbQ1cuJT5lyLg4IMkEh//GKw
+X1zfJCLv1Y+M7WD0GEGgEsp5+JWPTRfGOo8zn1ujv3+5VGj2xzChOPPeQV2waZNrGY3KXzrJ/Wt
YurAAClRBc+LtJMo5FLvgiPxaszn7v89wdB1y9LrW6SyZeTnoPbxOyX/ix+nvXJcErYNFyflf/yO
iF4+xNtzB1+Hdk7nLET7mIQRBpez7vlalzi4DZuROka4umRmXTtmVdM5TLF4XdgVDcnmZa/DcFCN
x0HTWoI8p9QtIdYdKsyYyOfsFVivGHPbRgzKHkMU81OuT5BARGzLlgAwliSnZenLQQwA5Z7KwrXz
yT6hQbuDx+7i6vmFGLisJqakQrDhav6OzrZfBywBvjWtv3SAdwF5IGEystVpFAgq7/dRXRIfel5Q
NDwZu6SanzdVBOn4E+Sp1MkYV00WRJuw/jfrFx73i0CspgkJkNWzpYGhdK3gAwX6mHWTJ8eExdrC
v6MLVBjR1gtwivGt7+QHSdwjyM1RBx0QgGuBd213xEZ0Tx3c9lkZNJXFeXhC+dxRIyfk18wa8WbD
l9oPQAy7vtCk+Oa21Ng0RIHU/z1y6V3X3YLcYafcJVEEAeJOpfzhZq8A8bO8XnBuZFHnahxFmOo4
ryNA0+PxfX6lxiSs8F8EDeT9Ev57MCULPGyQt3S/EawMLQHib/juQyE5MbjEihkMX1sXzWCJ1mXl
7vWTduK1XBYnsqEJBHJA4u5EWnch1ehFR80DrmOcdzv1N/5v2Wy30bFFavXuuEpbskAezhYB3EJX
NVXw+GFf7gub0WzAlP4aXQcgo9UQnmlu0G34eMEFwZW8zIgDFW3XRLp4bAmQr01ACK33/z7Yi3f3
1DIsDhons/cvU/ei94aw8cjhmKFR6BB8B0+0uyrpbDQJOUNJqBgULbo1Zxef3eUZPveyKqNxVgzM
YPV/f2SE3db8tBWJLIHFW+ew9TpCSJkqCCrcQsSexKCobaWk00nXe/vE5h+SDTCA+C/EkQ4svULR
BpdKUyxAYsXNr47l4NiALOZp6s/MjDggtXezMKLn6XBGNrdDqp2i58C5WZxA1H5C+S5m+ftnZI3n
UfLl/1dn7QfmjCIAUFuaGOxMLgwsWjISZns4uvGeqExocAqRV9A0dbX2FJYCPlyDlPoEnBLSezrE
M4Xtt9cDfGLeN5wXFQ6aCYqRTZQ/wqzyCAgFGH0RkaTy7flzRLBiSsHWIcXYKoxIyz8/5dl2tfMG
4JYGBR+ochgklQbY/Ud6nK1WuOA55eh2c/5hz1uC9X2H2DST6xxcSdpYs5X+HpXITh0h7o4TCYkP
sZncFXjSvlIG+QuHycGp9efWj+xiFCr+1IAGVobX/lz64hmz7Wr5mnQsalfOmGBzlTTH5DwqmhYe
vMBOVFURaV3FYAbhRTZz1LRyiSOaKazJJ6siE6Qzs6U52sCMhkQ9SPuxZsBuHMAIH5zi9SKYedjR
b+l7XsKwKZENT3o84gkRm7BDBYPy2BcMcOEtKTimP8OqXxVn6XmO7RDqAB12RcHfXFxT+0+3TFbc
3JGG7lcGxQFMQBG4P52CJeTIXnnJ2aelgg9+n8F8qK+PTXLj6yeMvhsFBnHXmUsE8z2AdXTUk+bt
4TT+TF/uYe3Ppgn/6wAZPthMwcDTXAefT/6PWK7MU9YwhWXwyp0gD0ri6xhwv7+YUEk/u6wEJCrt
4AYr4tzTbHKCEosVGlbagsRSHNjuSwg522BdSQBQ0vW418nzOn+YZcGqQiNO9zZTAKi0CpmAiExF
exrVLa37vB4W4Bayzk/QRNQHbT+x5pdOW4pw6FrMTPOAB0ztcA0BY/S82SAUsJBiFVVBNYUIqNPz
c1rL/7NG/2Cjpy0dHzkGqea1dZmqO23ZV3z2YoOueHXbuFddHY6fHSB8hESLNwQ1XMuNz6Ktq0aq
Y0pMd7NfR6Gi6gbxb0iGUCYdM9yFjJ5kvn20Q6BpDEINdBQZEKg+ohyh3bmxQwqlEtWOPh5HHReX
cgeN3xgW+pZRwFbjQ+hd2FKXW6P+wHKS5wN57AJ4T86IkJYK+g9LPS5Tj34BViQ8USjfugWYzYvm
ZJhJbzw8gAQZjDtXfeW2lu9yW8dyj0rLEAbYqCeshKjKzZCtO5NJWQfskrYVfcPZdlvPPdyGk3xu
KXgXB+Gh3iyyGmeOM41NU0qoHnIB5hh2ce59AbifTZ/Ex52cytvzQZyGr6/9/lJ6RNhSiZq074l7
1jCR9jG7RPgC4rBLEvk4zeE8BDme9/9Qn2TBKeb/wOiMVRrIlH8uKNVCzMkCFlLuxhgf/1ULWGwQ
VQK8o+CAVrvHtrmJUJ7KyF99z0fGxsTN58oMUZCfqSpo9Ay7rmxoypjcN9z0Zuigs+jx8Or9jRl8
zy38ws0FjhCQf+MezolEAaesiMGisufSDPOW2AzQ//jcc8lB1iio5PxBKw2xeSZywkt/OYbuKbY6
1e3R1gDVvK4FBCW++kokj1jV3CDt0z9PNF+MRNNNDBSdJNs9BMB3xL++/+Quk23N0RLMBt/oUB0x
FMVX7SeCKQy2Q6da2H7nApt1veaEK4tKaLwfXkZmZpXvSPG/l8WT2QRLpRepIT+EfUzDmy8IPEyo
pkyQ6ZGB+lNS9ZZ+QmAQkXlsZ12gq+pJBFe7qcJB6m8gJTJT2HKLKWp7uWe0yv7CpyCPz8qPEA3Y
LZFh+tzAqasslLTR8x9hwRI11aB3VwlK6wTFH1snYtN+cvMX85uweaJ24zSwtfXXviXqJDJT7VSq
JhEgmjD/ohRLJQH42K0Nhnd7QN5nL+47NOOfkiD96Inypdith1BZET8NXI+olQTLGtJl0y8NT57s
rHNHQXmLv1tlY3y8o78iM4NY3PLHEzSkXI3+b+q8du2q1CT8Wp8OvOGi/3mmgQ37UzC7dG01RyFv
I0BX4GM2kBs0LJSKpB0VrCFlVhckolV2uTaaJtRbIKdC4c8xRyarDzfNGzxoRvf/SnCIIj6xX7c5
W1AOLN1QHjrvq2AnbnvA6hKoZDl+xmLXVF1GVh4b4YFWI10t0hXiIm5AGcdVfE6RlpvBdiCoRbZ+
lGRtQwkj96muOqd9qwTqUIitTAYE3zwzMBnNbzHEPewz++dhN614ICvDyCVPL9Nqj7jOKWbW3Uos
M376Cf0mJpskITEg1YVETtc9vOXVKT1sfdrhTpbTgc8GcwsxP05gpyhS4JgaAyO3D9qUuU3Zngxb
VGgC5VyLHiFE1KEQo55CkTUdgUBTrCv8ccDhnTisMih9crD6W1acG4KtGB/Owf7SRdIx6Uz0gFxr
eug1uVTlLQEWTd0+CJF2He7aapANxz7ZeeesBDNXheWFSNBC1nchye+mhmagoPhEwVDbXqvR3h4c
kC3gfnt5eb21Hzrjon4imVOjV9MKkMYHmtUQd42WcvG+zIkEhtLXiEO1ZdYJcQh4alVyXU18ET9k
4EMASSLQk7rhsTwmYFIvAQMUuYggDHJvfW5+R2uw6X5RKgqTaZk8s2EuTulJAH5b3kQwwoVqzsat
rukSsrXTK48D0p2V5XnuUVO6ko4hE5ByWNHyW2yjZ9nvKo4KhqFJit8gT0nxGXc+UmVUCDC1H+Lc
2uL18q/941tyZsIjJZoPtGZWht2wKHIdbtsQBBTUhSjfW65Vbd0vkTJAJUj5kXoQf9e5AJlWpRFH
7y6C/XThlbhgeNmo4e7dAd53kGPJRKs+iiMY3IjaRgZKlmAke7PsSA8wMiCtMKwrxemktRNBRjBZ
Ye8n/1/iUrJrBQER4gNQWqTrBRtrMycOsmL/YKfNzJ+1HpxjNjsU9iaR+v6Ch/C2+9C6WC9003gY
OmRSIOJ4OujZuXuJSKwRY/T3pAljW40LDtyRsqKVgRcfPFk79GUFuMhZUedgVc8J0I/k75YejDcv
rlipr3NPDN3jJXQpahpznaqPDmlNxgbItfkNAnrW+GwAz5noHzBF227kmrznZPx/lT9XMp0VbMjD
meKXUWxIXgD9yQYW7A0sFr224++AboMmyKMJjUm+7iJayfnW834NYXycc03dRWoVvZqjc6bPc1zI
kq/X+Ao+PiuTsfmIrOURjl5ypEgctTq7x7Nl84Ju/ucyrR/KYU96FPes4ZrlkokPsAPRokGmECRk
CUVKADRdG+eGvY11YpKYCd9PwjwWBqva7Ws9XI96qVEeKmA4/Qc/+tSQekfG2yRFt7/+GgTbccAq
HB9/u1ldb7lJaaLQiXmHIkXDpKLrOHDb6OHg4HdUTef/RL3jJqPv9HiI0sp5FCV98gEGgc4HhEzV
Jt8v0fNN7f4X14Q2lu9BfbNurmHZSrH1NS4kqdx6zAXxOQI2MqeXV1LUBzVKIf9edgOi2N+iUAsx
osL3CLL2UFwkMDPxK+1A5mWU6hueKPmTXaJFj4iGBQV3laVNaCQwTjoSMAE81xENcptkekH2PNu+
0w18Hw9HuL2zasmVeIyZb3NOmzzjdtPAuwbYO1gf6sBl+mF8Yk1Cg6jzHdkLoPvMCWg6ZhBgtbpX
+cXtQ4aBNyuAr9Iqnk1QV8AErIiP+IJOxwG9MVdDewXtqCdxx9PTa+2XOr3A3+e5S1eMqqKkGO5Z
E/bGR3CTXs5TuYy6S/iItE9ju/0h9uwPUNJhkpqTCwqaqrPFYea/+6dcZdUh8gAKjqpvXb5QKZnU
VUcXs2VOj0exAf247+Vpdkyau4pWL/T+HwbgccgJ9flQebjvUPDUngnPcs0QmZNNNfgn5F/iuzAy
E7hrDnLLJ5wGV3zAe551a2KjO3R0gmz5aU1rSTGDCBvuYwdQEC55hKht9amb2i+TWVOj6RD4xZyB
FJ5iZPmdlI0umauFH60s1hzdGR4InobnNZkt12+cusGFgsypaXcatFjdWQyND83oHCF1omifrjra
LWpZXp1/3i57sZNcWeMTlklBbppWXAt5Uo4ql2w8DZgS69UP2qF/ase+b8VFnrr8IPS7WWR05Pfa
Vz/kGsnP5N9Cc2wbG8ZNB8UdKmOU42v7bz8jGP7b4gzhQZX/qqp0yDsx2B5ozV0RSCpEqLzmzdi+
3RoUFCe6joKRKkAaXOe8zuh4vITDtyp2dymsdQs175y/o7+wsWyEct4VD5CCPBYIxQFrGdRugJMA
NH/xAkH3a7QTcXZtKtVrIPfS0u6jV/7LU/nSdSeGP7KnCK7LLjPlNHuCQekf9XDfUZX4Pc0rgsG1
DIhmQ4QfSx5KeozupsUwcQfoyqny4HC7mYub8+VKx2la8WRaF+vBG/ZDkhDGyncMUBBVMgbj90cW
7FiKWQnrs3Lg/C+dkEZjH5UQOlD/Z5lU0wHuBehWpQ5GCMKJgJoWr32P5nC25Z/b/xSMqD8C4GEh
0/4bFRcGb1DAes5oCNz0I2C1POWPszYHWjqXoAuLuYhceh+7egjGdV+5PrgMhKd6zIArbdJpEkhZ
yokqRjHImX9C9ynLGcxub2rSQze0JQ5e5ebf4NzlVZP0vjps18g+Z8CyKbj3fs4dF9NWKqfUIpBf
xL/V8VK/nWE1jQgnVqWL3zd+M8YuMuzocdPA3rG5M4dd+VAn4zUkb8Kk98WZyJKKTqDb8u+8uBZV
RWwOuIZ4aYe+fF8UERn7l2GsXKwxgD2uUDrs5Sm0pdSQNFPogqGlrpNddwmLPcnPURI4fQZvBXmM
RmbGJG+v1SOyWyDp2GFg399L2WKr/awnH7NWhusYMdE2E74LzcCA1jf28P4qaDK8QKMtQo/XTvLp
Deuk2T67DsVvNM1Gd4wTlBPA//wYAfLWRBsz/CN98LAxPd9DXZMqGsuSlIdN2gqnIf5BcAW2lJsE
300dqNN4UIIUYulOzOuJYHz12jhzCXp/4F8nXljsOKrYKWOvpENXgVRank5VGnIAfqVLon7IW/mb
Ro79bmL91DnRWnZgbDcg8O9oMQ9REjvj5QGqQM9zNKOVpmW5UxYkQWmynNyM6O5v8QDexo6RByGV
8qMbBWB/bTy35TwHDKPbqxOPLDKTcxS/IWYYPy3Gz73g8oZ8naJsnoq73rBOTiCkHseP0uhbwubd
JeKOC0pnqKp3YUMCRbB3MhVEo4+pR5Ta8NlgoIguPgNAYGSuWgs2X8oRw1tYMXjCgaFnDUN8LpWX
2lf6vb1Oy4q3yGKGj04acp13N/yw9PcdWDw3EOhISw/HQyC38OUkai3fl5c2GdUTm7igMazlHwai
QF4ismvej90OV0MgvoNLluaDUwvRe0f0c3Guby0BazgQsCA6YatF1yG+1sxkmLH4RrmwgXWYZ+XE
NaVzQ6pyfFc3RkUULlrxKwXM5bvQkAxwA35ZV9aU5Xw47THBLQ2Ur0GIF5TKjcdOZlFA9dbqDIa8
TMLztfCDwM/iiNkqYZXMh1WtP2byCTaRLSHTMVGUoFuj+ZIOtl7edZ6OPip4NcM0yl+g9tJ6aZDi
pNRp3//Ti1Cy6RA2/+d9d1SB2N+6FpEeji/pk0L63i3hZCyNHeTRvFQNpgDgCVvAVbgQlDRhr7Pl
F9++0PxqAQYxemznMXVJPPTnlpWBgcyu3Q+ZpcJ2aOuCQVLi+lqwDfIYoqLkXzlfliu1VPmH6Kw1
ivJJFewZQzO4J+tw66BJe+krO1E9EM/Wna+HxLn2ZYV9qmZoAQDeaIQfJukr3MHdFrNwTvYcyX7p
BUQuemw7V3zjqdYuQMG/YcRVYqaly1EruNnvTeYY1acf/U5tdxBLaCJvJ0MMqjA4xffVG6BZB2ph
AYB6Qwr0NpR5H8pC8Nyan/mAazBp1mNpACcVR4HeQ/IviO89i8Z4UScMjN8CA4FlwCAwQRSvUq6k
KDTH34B+9LIAuFAjcoqBIbeiAQcKRsxuYb8euRtIou9IaKUn80Z9EdbxvXp+6B78y5KXnJBfrPeD
uovZQ07cC/6ws76e+VBem1e0kaK/XQTo6rl++sE2hoPhBW9bpCTNPkr9ZCErz5Yfa/UET8nXYegt
WKQoqQIOrGsJ1xqdbzW5ltg3pBwql69Xadv0MWtaNQkmQCmloVS6e4fZwNXrNsD51sER4zo6nBly
/6gVV9ZNh3B6C1rS5lgAOW186UGGTp+kZSmEBfINcINbNBj97CUZceXV7qNWrhVzb6TOzZswHpR2
2WKiqzk6D4dSx5KHI2b7SMne3WuSV2YPbt9jQEg5VEfyCoZIeRiFJuo5/0fAt2K13nkm3ppguJxK
1FX6fOaGLHqnBKLv/4nl8mDaNKREwiQWPTfGb4ujDCNm4ku3EWzSGwGNWc6BRlBD7gYSHxS0Ju5p
n/QkU/hHZX22NYSbB5oHRRAwBL0RJHTPSM8ZxULPGjEXuKt22urACrHyNRWGTUqIZlsbHUFPGKzY
adn/oBhjgMErFbKasoekbxHpE6k55y5+jCp3xicQvK170ZU7wFIoZMZ2X6Z6aHbkMYYHQ6b4yjmx
V25cMkPzka6L2wIp5t8HWUaFM1vURIyX+IPqC7oqhr9xkdMkMfOO5D5y1FwQr+OFiWFnAkpCukmn
ePh6nSQXCDNhUprqgGrBe0II0ox4J7CYaigy8kk0IgKIaErwsUeSvkF7s/fr8SHXrZrk9uDWCJji
ERAhMQNRgRAF7DB4hqKRJaCDpOkFlzV0QWxsl3z5aX08CpFWcy2wAr/F2t/9X4ahQOF87DJQUSLe
FunJsi3glfQGp7pVcBH3RxSAbxD6dgVd+5eMWo6oVBxl4s07PgrbSHNujnBTLv/GY09ZTO3psysv
Q9/I+DOwyuxuSxSqDtMGs6hhmw/goCUW36Fce+G7fZSwvl56WeTC4DVHVhylJCnPRsgeEz5ajWwt
IbVS2wxgbuIKyHRaaS6sV2z1rf1L9n0mgO2mKDDXVSyyDsMSj4lKHCNMJ83zOLcl3l6lLl1xb+s/
TBp3AekrqTWaAhNOnw5eoELBErdOVbE0EU7eEdcW+sMmbs8hKAszrkDE6qOPQOSdgVTXoBl8OJtf
X5JQgSNum2qlw+OIR+pXfI2YizcLsXCrWDXU+aF8UrO1rKVgZGLouXy6A28nD4RGHF6HqJwvRiw+
hfDrGzs21qczlsct3xdp4LHY6d7aER9YP1LytloIGo84pUgcuXZCb/Q1MbBskmgYmrtfXBauL4z6
fIN3cnNaGilJQunFJ4nq5O65KKrrHe8mS6VS0Cscl5XQRVgAOCeG/zFH2NI/GzFxpUlsB75v26pZ
XSoF5nzAQjeTMqH6jZZ3ITgEvX3FiZ85/PYwN4FI7utULRjRRSN+L5eZ+2OEh+D1Z54EplTwvHqC
ItsOk5E+UvizIWcUCXBn8IH6SCMMojkYQDzXk+hU4h1Z9xdJm8auXPKlJdEy67lYHZ7dXBMGNpQu
iJ2xHcYkDEmnGFu1OxWD7Kxgb5l0R4jfoRKdr9RqKmbx9DRd841VJJEBHwviN5+T/8MgvlLANghk
ymt/ZzJK295Ucb0fP/SULvbtPIH/6yvSUnqS+DIJFBSNBFDdhZJLs1TbwYO4E151bHfTIafTJhDr
lvivAFfjIBIsTAmctRYNhDkzpFaR0NVCshNK4EAW22T1+fa6b1lAwsAHPmBJ5fyRv4HwB/g60J9d
YyaQvEB/gSuJ7coaMmfC5HlwiFoDh5Lcma6rQyNAGXtykCpgy3QZUyFEfyrasVTXqtOX/Hjht3dG
H0zD7wn6Fl5zRr+IJh7MG3Ow+mw3E+EU6YC0it8tP6hwkFHQhWsM1K2PtnvaBdbFITUDCAve7TH4
8QlxH1gO7h31up8ImneepOH7kpr3N1XU/vy2x+3CbQzgoGhVZPSDD+IRl4HomDS9BI2g+c3Pujmf
iTtApw64cgLtnX/kdE23K5qXXTjQO4QbMgfDEtmktkLcTBttc2uyTdlTzSaVpTw4L5y1leVDhhzK
lkhtiAXCEqm4UvXGxmBUF1+8IuPbrcggxpjeCqBxF28OikqEIBwuWQ3aCwbjzoq2ASPJBpJtpJn0
dgaBB28pWRs6d7sH+softuCiQJPFflUIGnr8Z8GG3r6WZz6zzWkT//r3uM85Wa8C5gqj9dBgzV1/
fvzdLRAqU1+DCD72rY9SnMDtZ0CB1DCuCU+baqKJpa6qvNP1EeDpgbkKCZ88lTOAnzfSCgo/jfGD
Qyduz3H/rs6RV+S3V5kq5UxkmS16hFXS2E85eZSvRTMLaUhMYLRtG+6Yx36DkBoSSPCxGc5xdIck
6r1E61k1M3xNpqOdU3HDKGGdrOoKVUuf7DAePVUiKBmF5TJWG0ujuWpVGjoq48MZNUv/ubjvc+ST
F0Qtl4fZO/wS8gF2UeVBYQV+hd+Uu8Tm8DWAd4ZpT8wu/9rjYfYT1/oG3Xj1HkJ18CW5Grin47xx
gSZmpKQokp0bOChZNNjCd5VMpoq5cmcUywZgZNMJ7h/8XOyG6qGXHssUSiT2v5I6Jng77Va7/e2v
JYhOLfPl2/oXk4yewXPMx548vMnIJblyDuhcVRsC/VC0Ld+dgBues2P6m2QGMD6X6e2YWwLsvmYf
K8ne80cEOgoEEqJhiMwzMnl7TybvV0by5RYFVccBfzP+SNmmX4YqXCDc44UStVVw0zz8V46qUuMR
2qfxaUSyMO1mEbZo/sq3tVo3GqJwoKJFAakSeK5CCxe72cqcIyozrNbhLa73kCdwB5aKD1ERP7VZ
iTHriHKXwDV8g27BHtGvwkegLvN0+vunBW4RhUZ+YrE2cnr8y86N1ZLFM4xGHjJm0s5XFkmMNKq6
GhwPnGYtGWbftf9vSSW2aaOW+bpDWzxZfg+3DfvepkIcFX41a9rJGrXTRtUt0BU8Ar3s/y3ZI/9Q
/3e360LnsiQpAxuH2KWRluzbAF1EoNY8G3xTGdpaya23CLlvqmRiSPsR4KIWNPZUdH6n/Ob4HGU1
1J91GukU4ZoRr0RbszmtTgx00llj+b9B1FhXQ5qFcVNC5jXfdqAj3yBi0bagy81PQTANHFK6XIEb
yCvWkLa2yBpb4TYP+ipZB0Kd/uR7QfDZwCteDtGE0chTUrue0YiW0W4I08+HY/nGrdOeQPplUKfb
WNmJvQPSB+PMyX74PHWeU85+AkZUTj8jGZ9hNsUvI+kg4SroMBTW2UTQL26CNh/Tm4uf/M3Evpud
hI35OhKOkmKFgIgq8SwKtwD2HZ6pAsSep24FnuomOAP/pqi1861bTmGAcgjiFCTWQVymQKvQ2pTF
m07Q0mLcBOVoX0zaoB0IgyUsZ4hmLnRYjPddgUcHrnwMyFs42we0uniCANmaROci+ELBeQ1VGeXI
96x7J5EySIHPrqQhOjNIcASXxxM+Plb2pS+N+qXlu9uIuiGuaj9BuwQl6kVpWFYRGjGgfDOCTYZT
MH09ai8WmdLsDsT53ld5jS2URoL47YLBD0wFcoKDqxxpy/XIKF8b3UokGok7rCCJm9IdaLTuDp7P
s1G60bf7KF+SYgDg543infcL6jYbIK0o9PRQUfOWm6nqAoEt7la22CkTbJdPgqit+uEsJX+RhObO
hg+aCsqJ49FGG2F3Yc0/0Pt4R7bEbQR/7beDNCB/6jKZKiARjLEDb5BAutAEjN7W81y0jszOo1WP
ngCBNMZwNEl+7nPAgD+3xiyvVQsFmaqtcKaFnC7qlv3wSzrJayI0XA00gx3HXdTYtCNVRM18l7xv
JFVUjvEFVaWO9t2ZzBVPxyl5p4TEZ0h/xaa1DcvlHx3TIGRR0kgGJFIs8PDe+GljbWIyDZ0x5EXJ
OpabWsjIsJNiLsZB6C/ws1vUQ478Bo96Z8BmVttXe1xgo9ifbVjRIRSCZMYr4aECqTNPyYh7dQwB
g/A7/4wSWs5ya52KPcol7L6QlcUXv/yp+P5oDTrw2hLseMki0Rkfp1hGQk8aMZZVom8QlbWzEg/x
iYOD8hwuPVUwlt47CB1wKqNHe6WFq2mJ7wTvUMCAFIOO62cetdOGPA8fpsGO7vqdEJu2xThgU2cI
ZquFXdLJ1kzLNLW2D32G16G5vNe+i1h1LIO0t0u06t4WSLChoMzz80W9qANsoe4A1OcR3CK8NEvN
ecQvGOE9JDsugOKxNyYnEJueiULh/XjJK/9tD2P797cS1VEBF/rs65ERuD00Dexo/mSeQe0t/VQo
Mf7VSRs3VypRe6iE3KNmqqqdLn5gDemx7U6qR7Q7zLY8/7LpaWsprCyMvLKfh2AelhA0A/ZE6MGu
fe25kABnQG8wIkmgEqkpCEhnFr5HlBGXrYhH4UvpAh8ZwPZSS173GfiQ77Xi0VpxUszLvZlIRUPG
4+dbwqmoAhDQiCjiTE5KTO7RwVQyky5DwcVyNhFXzgKBAi/k/AMla/vBK5skYWeCTS5hjnhA1uU9
IUmtc2aMayKAbAR5TrY4ns99klgVU/JlP/YqxbNzePvgtdX5mgPjLjRocOzAjIKI/n2vYEN1TH0X
+OXS1t4hkxHtqxI9om8Qvh/EHxnQUWkpZ8q3/6nny2mGBXyATWKWk4XSm8559/5VvbiHc4lUYZvI
6arg6wmP65j5wzpCH1yTYxVnsG2GCXqdzNVRk6fe+cajOZg0PbKdgjootZmvGzG8ZIELuJyIBJIs
iKeec+/T9C8U3hJSvvHQD81svqi9D41EKWVnmmqlpynWz8s6ZKBAsaL3U7ZHHXdX6oYFh8I1Lj2c
zPxEDVDl27FQ4JjYspxCIpofrsiTP1/SPS9wUDGa433PRV/qmRLrMHLypENzJ1OLj9ltVT7xgrSS
vx1rbNP5xqOtMVJWNDXhSPf2RsfrzQCnfD35XcF/iJpjZfXXZg9JFjlXO7ZVykHtpkmcTi/1ZLEm
y4GfjkLtRmKBUPJK3rgoyjLqZOl+/LQtM9CAg536eBkr/y73XvGei8TRGSUsfMT7UzGm3E9NmJxz
8BqRyOvswQbT+IU50en6TPwx6oYVTkPwRhjIDjXDYdMwA2tLNN4UQy6ZW8PtuKUcLmmZXe7O/IWE
9FmyoNJ3n+B2MY43sx5T09kP+e7ZHc/AP11x/uBhf2NFJgvLCfQ7w0yT8SE36kHD5OCS1ZL4v2cz
8gwy1b3Pt4Y5QuyruyB04rpk7iHTsy3Ys81O63UhLEWOF2TLxePrmf4HO12l3oNZnUiz57mQd76Y
vK8y0xLWd/IbuHSPB8yvTUOJ5g7javR5bR6UUiOdMlaqWs8GYK+yQFyQW827qiGxFhHx9d9gA4uL
/CorQnsTf6S3ZMDQA9p850LAT3lGEPBjWaJqHvu1xeWeUqoFrjrUd5FKK0ch67K3hsgzzEoC624s
0C8DSR35S3Y4tSQSQeRbPYlkcDyofVIAq3vDjE5CFqnP0MyTSmz7z3DvMrF+3jdUUGL6QvW4P+om
Msv80ptQHcw+BsSVJU1msAlsFtTrxY5bOm5N4DKcA0mVf9qbw3itbs4Snfg6yI7edq9g0oYQjD6I
JkdyRnKMLTw7ivk/DAoTQzYLZ/bQAbYFfn7Gux9Qc/YAcoBGxnqIQqQufDXYAbgsksLEug4ZvQ8d
ZWGj3+E40JgvsnnEvTxSbfEdcUbOrIFIrtBU9mMfu1e5J2dhUulAYuzwjcl/c7E96j6piS7zMfyB
6yK9x+eIgdtbWlXSR//XXeg1/P7nYshk5Kee0G0PJOi6nx2dJypbw/QaICMnPGB66iwUpC/qJUp4
cPhabMAkhlmCOFYvE+ukJlcyuJwAGhfEuSb5ASy41auzPT+n5iTJKvGelaCnM7oR3CZToStyd5Vo
nK/gHpC/wR+PHORxQdPPyUgh6+jaslD8uUCBl5E03Myjek9DJmcnrXZeGBUP5NyaWXmmFO0CuoDe
ACOyNCaa6o+1Tadeitut9sPlWIvwzcPYlo5emPAEyTqEroQy6/uRnwibs3YuRJuOkMphbx79N+Sr
X/zUb6uYbGWqXcgx6dtzto2qCb+ONZ6kw4NNezI4fVax+noIVm6+6bSsdtfRQVl7fi0nJ1I+jgF8
2yhsB8kPC3yJ75AdA6YeKkOXrEcNOUjXhd0s5OqiuKABBPQdckZP0cBx/dPRKKZHoPmWWK5Q3uDB
aQJGeVfv5YKPBGYCGnEdbQ7avL2rdwgvpWw67+RHvztCYbaeWU9MKBRFhQUEOE28N1HCGPsf8fzX
n+zr/alkv4Gyd4q/zTBCrWnxFWV5lVq8cdK9QSsyHOLzVoDEonbO8m1TjOgdZWWbBMd4nY2EcnWc
Qv63eW6AR35kPFd9DEZ7zixJahvu79ko97hUDQ9WppynDiG7lpY3YGlzIRvXHiuvPplMvduf/P/y
Q3ajB2mdA0CC8M6iE3yGgmV2Caaw7F1teQfoBRwrUEwKdYJDXNhH1t/j8bi/56y3W+OsZ4nxAh7a
zBJX031Gcsa4DocZssSASLpelXIoiYgacuMAyK/Fm8Ynjp4bk4B70xoTziwq9DJriNJI5eAgkwqY
jex967MBVXGGll7WV8qw5CRI87BTTuZO9HTppKvSCwFOotuMv/hzTZZH7khqq4CXdMznmkBdnNVX
ehDW20jNMwjyJ0xyiCxbLQhwR569kuv8h/ewSCF+KuULOum2dzvL08uZtTUdAQ5MX2TkMwDN58UD
dUfjd4LlNkT6ue8YLYchDMGwlUv86tP+6LFMa4zbxrFnhWkRBzjEmmGjSxeoat/8UZLQ0MIKkiQo
WMO0O75Ws6WOp0hQRl6a8K5oaz3ZuUBfI/XIPkeikCyVlYPSHePfbmRRTayvpj7Y1IUGnT9q/1TK
aEc6JYqvvzlTHNyLVC0T8s4FQTEeKtRLfpALghSx56lRPP9QLJKu5TPXeWkRgMyYAXu4xYJVuv1f
FMv6nPbdEpkyjOAxroorna57KXL2hhzsFQWLUJPoXMKQsXDhBcMk7oyc/egvwkAL3oBZrjte5Rvz
r/yS9EHyqymvkRYXdzzyZuMSBY0vXwyEvFNl7XfyweitWbIKPoeyZsKvnfYSdru/h1R41qaz1pNT
uWgHE3F/42aajUWyFTNilr+WRWQVn0Nh98F4hOCb+cf5TDJYmYczsqCgm47Sp5SwojcE9x1qLmps
Gi/DAS8TR37cfzk2vqWZtVAJKphFWuAbKo5iyGuRuby3ljMJyTHKWJf4el2AX9y7vmf0L9NLAqZf
otwgdpLxoYUQvQvDHLH/edfKWNvIAI6ezPiu4OMn5ddcIQCZpQV9ZZoYQFrhv/RhpT4zeEGIsQuX
AnOBAhh56Ey2W5EPcwY9xPvwHKOCyFIDKdC1G8/E4l5AvD9Q8N8qPm7U6ESICBXY1+/3Qjnjwcr0
6Rj3L+L3Y8Jr2fwH9e8KoBWC4vlIb2tacZfdxYKZs3XQTRtQAkRrm/15KOpM6QJ3tgdzLc0iqg2m
glDoAuFxhuOrZ7o4uihagpwH/W4BYrKs1QgF96ZPdh+oam7UM00+FpBMLzBQzAAEcpFmYxqoNhKs
PGyb5MqXvnANuLHrnfWoLX1ziBdgU73NvudH3HlllBtYApzDEmFGnQc1AWl5hm4SH9o/0GGqIYTG
uDAdRTZfW3fZZ4tNqo2w9bLULUhnyJM0ZlaLnChi6tJdZ9M4WbU2Yv477m9z8Q9zZRXTIIzfvaPT
y9WdPhaneey4DyeZFiiCSerjOEpbpuk8fIbx3AqYqPDg3Ej+mWAF712vQ+qGjimREHGn5jngJtSg
CQjLpB9FtAeqkZwurwM7qJ43tJp5wAL17tMtD93c/jaQSv0Ok0tTXqemwwSgIejT+RIiGYXP0G0H
lJDcHruehc1rvJqAkvxKiwAbI1WEMSVlMfz5zoQoUKZ8tGqqf9JXaTnxDJfOHtRrO33uy0zJgmYP
JKg85mF6RkPJPOpvRFwnwrXnil7Do/16i4o255E/966bA5SD+atejhnWMBigWTDAS2am0frAb5MN
5/upZeIF5mJL+83MO20A8xDAKEQzkp3eyLmPRzo+kOeKPoUxG12QtRm80+Nrt66lOJM66joB9j1q
lvY/peFQrrG94cNLwYW3UA0IdpvL9J9Rx84USnQPd696TS5XWj43YH+1GGK9dFykJtpAFcng43Z7
OtcdWIQESmtWFVogQLIwChUeLZbl94RR0w6P0TTnQfTFR8+GwmHN8CivKNgmbvyyjciYyDNhgAhB
HAHuLgFCsEauX04ZDULKMnQt6CbmATMgeFGia+fpb7dKo7Ax2BSA44dKcx744UkMMHjYkQEHR74a
Sm4p7xnwMYXWHipFQOUPcUjsqi7g0sTC00dp3DeeQtM82xVhRvvYJOBZjnWK5EiyNDfpCpj7DaOM
Rc3qGXNuxFFGCPpWMeWpJ0nlh2ktCUL4EGQvA1uFZGth4a+6fEeNqbZ4Qxz4T32P1fy/gcphE95l
FllH3VknfrpTw+mTpcQHs1HGLmjP1lcCxMkKqWr8I7/cMDj/vlLhwvCrfV37M63ueRFTWoH7EU0C
q+FE4qq1yBHOmuPNPjN3M/CTysH1c5rQz8h6E6VdV1V8741OL5TzAYw5LZy8uvzd23D5oecBxfvD
MRyt7lQ7JjBPKEvfNORQw5U9FnhR7tCAx8vehOXYKZSh+2skcdOzZdMw7hvcH8ya4KpXJBz4SbQb
Mll696igQxZEhNcLbDHrkWH5TzHwffRb5De90EVMPEvQHw54GIW/ZPyb1Yx/wn1GuminP/PowUKS
h5Xx5dL7+CyEsdeFASxV0Sv+QuChU68Gsn+eNxglYotu2mfrTMVt+aICkCvG2rUS0tbgH4G48uue
elxtjVvx+iChiLT0dw7D2I89/pHHCnJPB4z03wgKjqhd9me3/7iN9spdDG8tqbBoG90wL3jgMlYl
cMTuPjUeSB/LVoZV+adKtL2mKkhbTnsyAl/ub8TnJpO8Xu/34VPlyytt4YJpbT+uQXNgoV5COb54
qcdIe7ifv2/Px7/9+ZkNjzqofvni6XjUD4c0aR1d77VHt0SDmOgvVl+R1A3jsRsR5cdDbNNgP699
w/4E3/xlfZ/o7blQQbSh8FBYwjxKQaXZSW+LmdPt/uMiGnhcY79m8D5GZwwvZ5mopJscK3Yi3FBJ
VnMjBEwg8Gzz8rhznB+Kc10XI08D0NI9cusf4ueZ0QrbMtpxKneEnbG90KVspypS9Dd5+RTXjDw9
4WQMcCJ/4hcMkPAN1aJdzwSI4qNSLV/4yIiuqUHJuhChN2cgj1RTqmo8GMsHk3t1IPHTN5K3BHkK
eSju3dkPmYH2nuBitrjPfbz7QPwK1rFPlzNbdFWJnoReEp3gfb0k5ruwZ90yvwgTMNHwT8Wcmhm+
s6DO5W8Wx782aACQqXRCutuZ8KN9Mtq+0TX6ROnbKvYTtlfyghC9y1TzOhkm6zk3LZ6vswCswu68
kl9T9APFqMpAZvxo0bqSrkeR+PLFpyOQo9cKGUbPcxobVjwB5Z5sdpGKWFMzNBeDeYDkuE3KYaC6
Gtn3f2dQEdcskzu0iP//lHgwBLs0W4ot7tSMYqYpNaTVyN/ng/BNiG69FdGqbddMfLjz7j9+XJZX
5bkyAqDqZb+A5fZ/5HR8PPBUW6M6dyg7lxo7M2auo1Hd5AzQU62uML2amx+NLndZPseRkLWxjBZ1
dRkKtCo4LYWHCb/ZfCGi1dDyGp4F4b7LhLuIlOVhJvPajSxntsPY7elq2IA2xB4H4RFv8i5HAAKv
uaKWXmHDFIVZvRFET214RImJpl5rgohEiP9O2gQ1M0hNtC3wr9hlts0M5kTe4kSZezMzsw8F23vK
SGjPeTq5Rs748+aqbWU+5RgmxxCajtMLR/qf5VLOROcxrUWdHEBbppaNOWH2AZHFKR8Y5v+OER9h
YytJgkOWZyEavHE4iFX+oOBI5dpgdMZ4AA8Ku+1pwWDHI9z3hVX5FVxggSXL5Pe9h4ZpTk4Qfzvy
IWtjcqI802IzRSgr8HIxnW0+nOvN7mV/nHUxLwxNiXJvDFfW8wZxAnDmF9mj8SVX+1hAU/ANz9Z6
BpUfhfopbmlWIik0jhBFYea+hjZNyGHQ4Gh9wBs2DeUxqDlp0gla5PhgdeOjoa6VR1Mb0XZXlu+l
rFGoljjRmDk4+9w7tt45fISMGZP3aNPT783bFL1X15DDoFQc4opRTRsGB7aDbQU750d8nSwmMtyz
UOixgqTz4Ce6GBheEnNAHKSCbCtm//ES4kaqS+LFadbOAFUwjGZFc65LfyKuahkr3fQnBBBwGhnF
X1YPU6trPPrfZiTdL03O2U4BY+/bRkPQ9rixMeMYPbQQJpvBinlGMWcp8Bl58hfveiKSTDydrgv6
AZLZQ/6fmMhfP1vKNOtsILuG9Xy/pHepII4wqYYqG14RMEbAeBF2okv0VS5mUbK6D8HetE/rb5bP
g7mpH72tsVOOPBCrzN59sEkzmRqTRPW0yTOpdXgpDrSdMAANIvk/5c82k2pTFIo70Gdo76Z+usjT
0cJDwS+SHaQXorVwLfSM0779VLW1OknwfYamOkRnJ5sI/oRgoFq+6h6puiDxQNYXx11wlbdFyocK
1RSE5KWYXYneWjBfz4Udr07AMlRd0eEoIbCv5i84KB7GyzQi+X9/1v6dL7Bkc9hXn/AYHKJ1X3ls
9LBwdj9eZvt1LvWuSlMyAQucFBqDVRPnKWo1E9uJRVI5phxGCUVoKZuijH2N4KGUNWEnHR++JLRU
EkSCcyNVQ00yZtGWY9UXDfKUschSLmaodlRg/79mrWZx77TYd7hSRgPCufLy1QHGJnCQH/SmLO5r
HQTmFBRngvMT4+WIKNJMDqahDsQbBR58OWhswIfIxiJbF6rDa7B5yxIAxnZCbnUTa2n6gJQ4nVZI
GY6wKnUiYivXJetq8GYtIZ7mNq/4sJNILOuEGCuvW2q7lasw+ohocui3ufOr9P+HdDBBmpdlhsJM
a15syM64En/OcaazuuZh0JR6vJC191P/irFp3+iG1QO8280nANoSnlcM3wp1B/PCbq5DR+QwdPPc
TvPT2urV/HnbLa2Un6Y2ItR2zTYG4b+o4llSzlOobpmJeezkC9ROJlar1OfsP4Kxz+imlTIuufHa
YakIaCeULFru2DhCgXQjUjc0QfInAz1+KSwU93Ox4MpbNCd4UbUBMdQNNznAvalhZku4W72HotDn
VS4YrWcrxEL4vyRa273jkJOAHdlZF3N7UeKL6zGF8jthIKFkbCKflBSVSF9lZvaut6fRzLfAswRi
lsAHOD8Sbkxx73/hBMaS53BbC0nCWLtNFNjup0Z9n23+zoq/1TsWvGeKZDMCwSBvU9M+lVfE/YOt
xghjsOdXFyLYY9FqSJRaUQv8Pz68Yi9PLZjlrWWiDPFOH5gIDzeWKIe5j7BDN2di+q3a7meS3xKZ
YwVx/QQZaerUo8/SeE8FGRzGscXfVr88W2kafaQ281dlLUgu4MiobNk/srsi0j/HUKbvV7zdDl5n
QsCcs7a7kg6Dy/tsWZnEp6/w/z0uIGAdfJA+zt/XNsc/7ueHIcelDO21PopYG5QFlEqJGsyK7hRZ
HBRHkAR3becSK2V0bAEgcQLrnAOgC5oB5c9UtJWuX2/PuJI/RhBKLRzyjj/boV7u/86T6NWsUlHz
p4YnfClYOrnZn3Zab7zfklD+DmMe1/tm9DUb7niXjDSLrkgT/iualEuwFHSNrIUdZYpSmuQSKepo
E60jLDYGo1gVdqMWa1zKQcAY+4I5d5hQMgo7Ne1+vZic/65Bp3O0a562b7lIpSzoyVy+IRSV6ppb
nZoMY9LPNcUeOkoZyADiAbMD16iOR5mDzgPFzrMyiwRDuZFu4FFRnwo38LqPXDivvyet1NCexpa3
YazdxjSULP++U8Atvnuoe5uqC/C/A8Ei6+YjNGGfUdpzdrt0Iz3mS3CQMp+lBCUJDnGTewGIZhr5
rWyIcdLPInXwmicZdhqi4qAvTmFrERfBHTVp3zWjITSIYuUxGIdSGqXLfWYNeExV8JuiIE5MK6qT
V3qsvIk5m2tQ11RvjPz9SZsnjstEFewGqgFewsYXk8UcBDEqoG/fuUkP3TCH2Eq5V41MKgpQSpwd
hcF4pBf+LxBolnU5r56SrSz8mEGzK/o5Lvhn28FyPCKur3NOYxyAAFs4YFU+UDrd2AHjGf5NE3VP
ntkPAZYbTCrfXRsOtPHsU4TBWVtsRmvuthEW3nMecriZFidSM28fvea3rKwBlDMUbGhb4oIzJp2C
CqOFm14YSQ3gjZilHm38tl0bbdhvbl0FJ/ZzWtrFrdtBTNp84XBrbH9vn/cXPR6jnqm0Xs0pXtdn
GGxOnHYYiCZACpijU0VHHZ1nu0Cxk5gGPs3kmK0MY/uCHuqOCgkkNsRnk0DIaFFOlqlpLS24nf9X
Sp263Dh8Umai4wT5UrrFRXf+omQd5Dd21Rc6WL6+YJ5DxusjpzFDKNGNB90UjgsgPnxTPzBqowHg
7BoPMoeFE7MXEdP9Rm7Awx/cbR0oylXmWSYTlYGv7d+DhpTZTs6riQi1+YtzRdJafEPvnRBu9wDd
ahfdUfagT38hoxpf70Pr50pmlqu5kG1E3CeX+wsHZLafCHLz084jvDHfqnqA7od2jSGTbzJtDrtM
3Ot8VhygNCFII/LVZTCPYBvdI+o35wDH4OmMZ8LL918OiPYdEV8CkxQdrNwOh2n8PsXj+LJQGH1N
3F42ZszJku5Bxu6h4IfEFpJNXLi3PeHLl2DBxbatTwyNILEb/e8g3px0b2H6LqwuU+4DqCEUja+q
fink9YoN6KlWWUNz3nCSH/IqBg1D/WrikhMpAJqwsFgtYStodhEHmMG4GnxlYKhfI5nury3WJtIk
E0WwUupV4SYFEHvNZIX14b+SdvdNNdDFzcxB4zFbh9EdG1PhL2/hNy5ZG1q/zwiZEoaTDSQekA9t
uIVJi3lYnc4wHtydVng9yf6xkeaQAbiym3v1huFSQIbAGrXCMX+NwFdWjJxXzVwGlRz9cMQTfVrg
uaJObPkZ/Da4V5Tf+fpP5TGt0INd6IAJsTBMWQroBQiH4rhw7FuQin35TIYbOgSb3R7xEIc9qwBS
Vc3DpR2Mt/LWmmp0PLKkOZdOPnLJvS8YA/8LVGHI06Y8OV6OehGkFIUIhEdQOAj3LFiVorlWr4Gi
NJjePlFztn1jposb8y5wWB1wgYee5+/qVuQnzYIyq9bF6V2G4FkmWs6VE5MCtuSf4xVqYqwcEGDA
4kZugi4ZWpfRtmg0dQCfQ7L0Eb7dBq2eteWJDR3Ct713CmKwG1i8zc8O8BhoNDm3wlGTzfRdhcbx
q3Pg8NGzI7N584YroxrW5hyTOdepIe+kEPjIky0nIzNiQI8y7RYYXgbITDRiX8rb4/ixsEveH8di
6NXGZQbtdfmsRUN2UMmZt23rfulUhd05/Gtz9+Mu4K/ACMEjR9/9tqDQlbWpecrvcbdeGViPZHLb
BvgPCyjHWY3x4UgsyzG/6h9e0KpTyk9lIGlyuKIykCgo1GvkDuqlKmEMAX3VdrzYaVtg481Dlacs
D+yHqDrcvgTWP8U9iF4fbtO7JyzZv/2hPyZNiRvfWRQ7VJ+qeCDp6+ahSnzpLnkfCgGE2nPB//UK
G7Vgv1ODO6OOBNkK7c3yER+HaSGu4g41Ee/TZeD11CokfCVcqz+M1t83R2mYHEV88Qw/OINSNBv1
zCIFwDXcTmduIOAA7fd5KrKwGw2pexRQQctA+NGMoqFzIIsmdLbP01Gzhnlht2FA597pr8HYhAKY
nW/vOfw4X312u2rj9jZtROKBDOk6LLt9ltN6CEKcYsw2/Is5kpUit8Gypzc7zuDmJHTScr/dx2ik
HNBbc/E0m8BwATry/Y2LNn2s1I0ZUU82npOJM4ffbFnLcH2sU16UGIO3r2sAvgOMPG0x0R3Lff0R
igMxq/Ph32gwLRvauAl+WBFE5wT1zyQGqsDmxF5MeaG5RdKXRxmr9ugJ1ILTZGTEEUCqbhYHH0Fc
S96yx79gt+O+ydo7lS9G7a6TXyxJIQq3lDnA9HTF1mKVVNVrEVSTGQcYd51lnuvNQB9Mh5p0IMne
eAPAZBtc3cKJLQFLwL4NDjof1TA5mcDLKicc7BgGQX0fYjsJo6yLzHXLKr4YwEDjhequwZc5TXuy
8J3aPgyCItgnEABSTLRDsd7Nefvht9bSWqZAuGceIMFwKIXU/2OLd99mHWOPjoGvc8GlyfEbRoqY
eIRQbmTeZHVD9OxYs6/epaprK8PNAd2huxsqm31WsP2XspivAnK65PU+v4nKS3szRzN9DDxBXFcK
X283+SYESD1NdVUbvxzuyD+xoSGPrTJopw6vTVW0B0KoLDuO1SjFUjmBKQ9YLXuQZThWwVWPKXqn
Aq2hyZy2fivLiTXmFE2Cio80zkwBgqPzyKdqnyMQzaPpVbsCiWqo6WfhnBxxyW1pK7kZQYwobTsr
hxhNPUkCgn3OG95rgBmGewdL+yeKMEz4UAFs0BfeVF+BhxcEsPyyG9R4a6NElMErV1ZuDJWTM+K8
p+MD2Mf0iS91x3PBfyxtpZdmuFp+0vr/vGf7amqP58Yrpe6T7sFZu0/EMn4vHkyDmsufAsAynhmN
D5+lw3USxYvdXiafzcGXIJxYMWmzlilLcYOJRmqQktFrcFahC1xn/yekjrqtshwMhmpxwa7Wyop8
HRuajiyiFSyasIhcKyCVCycRGcTuNosbU5IlILhWAbdrg5IoyfYylSq2OSV1s4n03lFjDQerWsxB
fdmWtYN2MC71H+Tg+ljh71r8N4GEwQ6mtdyzcn3lUTO9+1KtUEEUt5FLYbEEhwITXEBdP9UvA359
XJJ1trgA9XF60O+F16/3E+mtSmLrq16j/VcZT+KAwt2lVtY3juJQfGopY0PKVyZDdhXUVS5XXs3r
8A7E5yrQPjYobDqUQPRg25XvQdgmBDfYwOchY6kBoRnPu/0eqsB6rNpoweaD84sn4NdpQaphMLkf
MftxkrozWL9e3xQiuSQJJfPw66zwEqkrw8yBeIoHyafW5L46gm1yi500kgFspOuR4AOeDITW4Y/N
02jFHx02/HYJml6kShq26dZ+t43jIyfOAzEkLk6PtltQBcp5HxxMcjvgZO21D0gDj8ZLHRZLvGn4
Sj/v8m9ZZADq65foImtN0Kf1mGKSZ/uWY+qo24NGqb8GM0DbQl/y/DSJK6tm8CGMfR1O9ba748Ex
A0M/dWU1fLSUv6bHPU+tkYoaTAFO3kJjdhd8UtquNmWlp98IAVYMzfavbztP4RAbS36Qzvbkevrw
vRa1iBqiIAv+LD8TmVfFAdpGewbqHOv8Ax0AyWJzMDJppoyNZtBFV5Rq4CF20mu2uyO6rFbbCfJB
oyEuUSmdqUa9LOP5gAehJf37GmnXn/bDMWxgCtlvFEUKTj6Hu3dsAtBouOr3bzOfB/rxvyOGA5jT
35pp+wUZdpDfZ0MQ/+YoAtnxVi7bGqIa1Cw2WZi/nB3fdAn/D/dBZ1zpWy1inF/I749hsIAcr0ZM
be+kTeQmhvVxidb8BEcgtqdAYMCoV3QWiyb9tPXl2df2RC75pcUH0fBO/dJeV0xVNJ6Cz9lv7utH
2i9WjbtDytMlXhK71fDPZSXeoXkmSuh1+UU/j6dvoQQnkwVRJLXXyxq6zx0M66GNoxNvOgPQCujP
St62Y2TSxSu9Lr9MmByQiYYsKBtGW3CwFmjOPe0yxQw3KAHFzMr165yXKgYzpyJbOnbDFAwKTpng
ndzY5HL4K1y8g18cjCU7awWc+LEORzfrGsoouCcRM3wcPwiFbKovW37ip913UchqAcJOCbgc8VgY
EyYTojX54amAwqDoJ8z1iVnRZrS1QFL5tJtgl9MJuIx+O8k1QFSCx79Nb5Btyg1vy7pSqRxMnxoz
cLntxFh4bh8qrtbw8EieGpOpR5JwW4An2QR6HIthG+ByUOEsYoW3iIaGQM9wIGGmo5L5mJy4ptXI
tBV5/vc2Lo1uJzWMW5Sw1TEWgZzv40u2+oCvwHRI8jWYbTmZqMufG0MfIbuoupT7i3AW4e8WgmnA
6plJMl4ThXoet75xXPcy+Qeq3LDIDBTTnNcAMveerc8asptgsl+vVTIPna/p+4fl58+jV905DZLg
ki2quqvdf92oc6D0lphPFA4MnTEtYdBcWp6uiM/CzNYEgH5PsuMMH1q1f37JIhpjn60TWZXdObRu
RzzuRcwIhjaN+wjWB3zZpMCVQxwgErApbD9Dc0fP2/IIGdVA3sWyHQt+gvBxvbFzQQoMnY9JtaOb
PH4FBKaeYWfvrxd3FAmRRf9+mlSALt6Xrd9JpOiz89ma0ya6X6EK0SqNxWXLhy7YpbFvjG6R53RX
kuAMFZ7LkP7F2TDn+cwdKaUzvWLMcGn1EYvTh5k2IhP9E1FYOMaTs5w6Lr5Vikjky8yej4kD6IQc
CabGszBBBOlXLEapajizV79gAUYUM1qj3SyOVvDtpMw92PouKRFyp9+HFGtKnxMnyca3aYquVR4T
eZFXx/VBAT5i8vnvJbKH0I7/tn5/B0Exgf8EgAMz567KSSQVckOxpz119+UmicqBSbUu7COyfsoV
5JiCKR5ohXdx+gjNIAs423LHj9H3M4UdwGN87a9NzzSIIUWEP85GHEkRsoFVYgeJV0bmibj8PpqJ
cVhUdhsBgNyxjiIaYZRT1GHzKKxVzX/JLQwRK39DUIkv+CiaOfWxVkN23KxLVNE2vKMbdpXbCxGH
ULmGJ/YukdvmwruMQRO/PfwPZA/GMGiVO2ofxI1LtACGnS2noa5mbJAhAI9inhNgzfEItUB5YgmI
yg2g/OdBxt7V+YPP28C//jhFtYYceUUU8EYLSsq4l9a/KPuiTzepRn0X/0fAVEeLkFXd97PzxZG6
qw1cGiwd63X7Mr92TZxD5rIkkty8l1Xf4jr1uAuhg0mLVBiENefVg4SJNDEKFusehQar1ZSVQfAu
TBtXdTE3kPmJxROJEtwOUnDC/OA0QDXfOcu1IBqrdmHq1OtjnWc5REDr2Zx+6zNlQyMa7BobBSdU
dTAJDGSXvi8QIb3yHMl+PJ4S7sPdP+eHo6xM+2YP3E5wqXKv9wbPx8KHZtS2g0hTdyDDwTrGaLDL
SIeledmu9WafCA82rkhGroiY6aJ1r4VL4WZEh6mbZmdmqm6WPH/U6r3BoZBKYMxq6iKnbTaQ/VOr
gh/qy2i/XC/u6qNfQDBkWBjWvBBEdfZOrg5P7KtzLYVqEiUdsiWRriQ5pgzhhsbgqeDfajeHhH4L
6y5FuPIuAzXVd0yJtiHedjaOPL9XMkw8QGt4LlRNaG9SY2JRVXjy5dQPA39v/DB4mBxxb1hlf//v
rHd7oaRomn2x2A2Zf9utuJhGCyraXdVwPEkOaq1DI57fq9pBoHnfmQq5PhV88PMufDoBA/oIAYTq
dWCnQs7eTjKufmNaLBYclzBhKHKUdhfThieG/Xm0CXVNaLJxvV9V8L3Igzeo8Oi/jMPYf75Esw8o
/bLWfpTYEzHXubU068vrJ5ak4yb0YL4y44tkNDwe+2eL5KKJAtbqdGC8sndWQQQAi8640U1QbXBA
S3lyZzCxzeo89muVj+4vgxDOXkU7Q6gFhYAEtwWz3xfF43fzHlmGoeKri6cfLN5iZ2OlDtzuIudr
Y/Km/mcZrXyh92pdzdAqp4xpYbWfOuABiTdcJjB9RtIm7VUqVztZ0mq3RpK0ojmLl48nEp4Y/2ui
apd3XpGIjenrIAetuXQwV7x8WoQTUXwPb5wBsJQEPDRooiLdEMx6Cm35SAyQtAZhwxl2NRk/k8Av
FuUMxQK8U9dvKuumdCOmtBeOXiJQM962qbFmVOmUjmhZtfFBFC2+9LYV3UnP+1hhUL5Fp+uVgSbv
5Je2T+L/2ekpRIQR26A1BtGHK8GHsxBer6opWBF9Uc8eqQn4SE6m5hIDJzNssFUU+hq+KfWOhH8m
XqD9oZeOdcHifTuJYz07Tdggdl2j4iu84z480zke3gVfkPXJmo0nttgPvUFyZCsh/DY/VYdQ187M
/tlpxoDMGpsrCfCFUV/HYKBtISRkFoVDgjkooCUCDnH/7Aga/UVLz3tONyCKz+M1fRJghA2wswuc
tjEyFy3ncNG//Cp61SavUkpYCkmjMayYO+v1G3266nBM0Tx4b0I4ThqDSY3YCC3TXdUClf9WSLgT
R8RhQgzaqCKuWsbHYVrufeRGAcZCWi4wjl4MyFzh5mPl2hdlwFVddVb/CZHOQyaT06tVN6bnLDs3
RjYoxzPRosQTlHbitCb4YK5qJ47N0KRzNDAcaowhJmmXK+Nc67TO4XOmE+sIuYmDW9WArtM0CxKM
0RKf+1UvguRAV0gFiJn/IGjHZT027I0cZzkEAOJyGaule1bGUUUl8YgYzz36sCORJI3CdupsTPE6
3mXj87dM+vG9MTrMvRAEslW0Z/DdO9LOw1UlXkTr+knXmJlF5q1SDtyHZiwhGJ3CYRV2rUv4tm2s
X+Lg70qoLE58j4YojY/+xYpGO7suvVC2GaIj23E7WOPTjHlO5/g/plA6lJOEKShqVR0Uoxa6duNu
2bzLnDwaRjRL6PwX+Ap+mnc3U9dvcblf/u/2DVoZ6bRpDjapbiTEAa6QJ+uSAy/l+wQ9t3neeKkZ
kT5GgJnHyQVHKXafHyKtecPE6JiurhvpVMpoNGle50I2PYSpdJ52UAH4OCte7dAvocAXuJhwoKzX
74pb+aVzxMB4ZcQ8W0FRTN6Qy82S+wdHtfjy4/vDphWB6FEAe+d6c9Wd1z60GKTOEFO4nGRh7dKC
JCDM1CkZ7wDNUt1wkAd4NGUzry7Azg++CQ9ZfcVc1osON79EScHE8EFc7IEmNo6/8LC6cONVO/8R
ppp1uvnYVo0lyUbuJiTQVmiNUO/8gn6poFxq6X91VNPPlseRQ6JId8Lm7YqveLJEGq7lbCzMSjBq
MWod7G97o3O1QAxZBY+FzoCBwK+Tqkghrzmy8Lps9J3nwqyjnjziOgMvIBZROWXyAU6iFBxHA6lC
sJswvIzzVrZ7G/J57iXajMrCC1Cy9700Y7tWb0VmR2XZ6IwEoeU3n0CHFiJruvJ+5A/Xi02mQkWU
cB1Nls6X9Y+9L3CkvFl9GIiIxam8pWgm17Y/gI4hkfZHEi7qz0iAE4g54Zom2FDwxkZ2mLZ1MfNt
+Oqwb2M9vTyPaaInxk9Rmhn2awyHMXOukLqJlF4MUM8LOgDY7703BSk9Vp7zRATXRNt0HlSseQsK
Qsd2l/S/EZXpzBF/0pD51Gv2g9P0kUTV6w9evlyDFuLlMIn+cBBdYBhi9pqoQgVBBRhwvTj1dyEJ
dLTx2of4Su+1fJuP6Fsuuuq+SkqnOou1e0Xph9wSm6ERmuGrvC0/YCr0n+5E/a50XqJlNi76SiXW
mR54gBbKscVuKuB1ZBdJxRkCNuFd838C1cphxaqC0A15FPCD/XYw7DntXBGIU2Mgni2jm9oaLqZ6
0e+hHlOJ6FskB/o4AZju397yc2vWYicKzXhO/FMQ2bu1IKEdyPaq/+BDykSjlg2/hI7IdT2cZVU0
ZkMOz2POPVpetMXlZDwVJBlUuviuLrXxxXmRfXhfcrVxcYixAj1qcFXk7XJdIIZhbzOyRDUvwhaY
pH5vF2gpcKrkh9AkvdE/5bFkK2kE1Pt3OQr7hv2gDuDipzY7iv68zMiTymC5bKvsnxnTvZXPeRWX
GT/TTu+IAecF5h0fqCFTozJ6IiQX0dvfANju2KvzbRICGN/dNoYacO7JDJJnHvZgBHMsOYghPviU
VEMqeYTynJdYRJHtxigHkJf9Z1Ey2ZnqJf2iqAhfn7FKrt3g6L6czJnaDk5FYTM8mxB0kYTZlavR
nGjsmXnAgCi1wksLgASyd0K8La21lkD/ZEsCsrh470i7gdlsjE5EgwttvTT/s29GYrDMKWGrXIQS
nePUcxl0n75VJGbIlFsxwm9Kuq+i+hVGmkJPbaOn0pxuXVENFq9xInsWla0SY1ag1O7qjtNs94qY
NIGWQCmx6kKzEkeQu/6NsNkCVABUSz9GdsHHjakHwxiJABzqSWdXDVLfqtGZqXwnYzG8ROaHhS6n
GqSK2r2jemwbZU5MDeLyNITmK38DvM5pR8sOuanJttOAjUSWsHANzyYn+hFzt4McbVIMIvXh+EMy
Ku4wzo4ZNkSFfb3NAXRqkv2VF3V28LhtAWDbUgN9H66/PBdPQo1ZFpnhkX+gZ2gKPIYgFL5DK3Xu
HGTA6w2I8wyRZSpdyZoyQ1ARs6cVP+myoL1M6EDArWlH+D8iMg7Vh9PTQTVqpvEx6OQ0dRRoBv/J
VC03tOLvGdfrCM0wVwytMIwo4YbOA/bjYH6so+i0UQJaheOYj0NHMhtK+20/qheRo5Kh68maQeBo
T2Fo/ak98dwOtgj7MJ0XRZXchEEsMRT9a4WlDosIdzN1+g4aOwFkzP2axqPLqWssm0gWfw8FMXeB
7wk/jbno92a3ITBEmlNXA68ohbQSBm9QlLUg71qbBj/+Zj14w+8DWbESnHIHIanUiZL8HgruZha5
yaIlTptEv4C/Otq4ueu4Uz5Gfz+g/04UURWd0TBo6QM8CnXi0rvONwUHbdUN1igOPbglSRZHgdF3
G9tRvo/1i8ad7UrQ46GuUfE7JYbrcKTUlNDq38qd6g9DcYD5ubpvhZ/5yZ98gMpJCULsyDZHeHIw
u9ehGKQTo8qXEjphRK8UEGbr5ZtdWN8XHY0LZmr7WhjgkbDjQTkyJ2UaMF3rItMwPWiokcfbxaD+
55DaU1W2DHJXo7lulz1RVtMy5dFDIT4bXYJSoW9bXH8GfvXmwRoAnJX5TJjk7feM7Z+qQ33mHX4c
H04dTR42AExIe5OrabeuL+SF0LEy7wn+b+fapCnAaq0q7R7GidVEDAZMhPIxlMCtYdYkaw2vMDRY
oAktjOmjZAz6kxE+pf5GyH79DR9KtEslJ73bhJACGhkXBc9WFw1SfHONx2z2aISVWnZs07yaFwyt
kKBofZ0GhYVxdoSbtvB7MtOmtyHzKbP7D6CUpCU3NZnKx7DVVURK/HACXSBqNLu84Bwl0r6Hv2cL
YplPD0+ksoQJYwtS3/LX8tmMwA9b2XIeLt6vCNd7N7plNjhRZGODJRy0/fk+wFnirjW3hm2UQwCP
oxHSik2vgxno9F3ThCEhnVBwAyfXsumrKV734GW3W5gaY6eDHEFGWYHxImOJ7WNq6cygjdYfP9q5
B5/HluAmXoiXPRPwi8+Oi6PseXHId9lPNXXAEwCnpjKG30pO4Cq2+BKuNkdoLnbRo/s7b69I0an6
RNOgCqAiQZYKlnWFM5G7ItfGBe/SYfLfk2cJjGKE66eRjn0RAqteClxvhCtvQ+YHIobWIRJ5AgKy
SaE76xaRKp3fGIlfhwwfdadOyM72HGunYtdva/rs1dL/ZGHycYMvMu+sBFYeS1PLfsJL/O9NXyIX
PLei8bz2Vc5y1AgFU5yY9oXN7BF8cHWzs5U92PzK5PFPVPIiHgoLgWUtaVU2snQzVgOi1PijkAQw
8NCaloCuJa0tZqDaYjIqlE2f9M0Be5Iiw1kZS0jtgy3hm6CCv0uF/eZ8BuUGdsI/mBta3noVHkfp
dAnFN5cACiAUY6//DSsunhpKJmRdK/fhCsMntCQNe6ZOSKYnP7rNtIN4VNgFkqnGyOOl6n1Js4l/
Yl1L4K+eD1AI2nY5WqUN4SCuFg7VrpNEwA+wdRglzH97r0y5yVE7YwglDXIsyv4RXcXOTnWtxfth
ctashp2dPP3+PKrbU/kLAw1PFBqiloKzqAdBkg0pbhyWko6YASsJFt1zhlE7czin7HSgRGupm8yh
ypOQwBvsw/FPSDkS27ZDvzGg/+pCHg/mCVMzeIbT+EkbW4WyT+nYf7NGBM8kMvowXOJ8HvSi7Zps
w/h2kXN3r4nDkTxSeslMGtf5k+OlB7AGEBW65JlmfXiaZcPYsghyB4VpqwfB1wT5QceENWETI97B
5IcXVdX1wm+dBwxp90TeqPragfhx1JHMiF3GPuE4TPL+6ZgIB8LPYSc2IYR+uiandMzf4Mq6URwh
sKxEpNYoe+SWsZ0D5Wgxk0bngUyfQrraVnGOk9/tjK41qmvkka/kkNeAdPPrKaPrJQPrEFGU23je
hMpwWd6+IHN8D9/hBYDV0TFp5tR1hb5yk8PoXRxEEk/Z5q3qz4sCfn6xfHCAug1Nr0nExe720QoW
g0u2kWHPhEzEEfXRUNuIrM+6562TbQQCNOV/aEyGP+q37m90VeT1LwqueBLajxY1BGmF1gXQgnFO
wz7YPZ0BZAeu2ysA+rv6JPmYEuo+ClI1m+xEiZ9AeX9xjYdVgZO7zhmnfQIyfvlNVRQbwOrZ5evY
f+SDMSFtlAckXeo5JIPEBNfQjL1GgOi+ZTpBvljxA7n39wcmTVwXJRExPjLNSBvxxxDM7blNPBdx
5w+QrC7kGHEHb4tKM7yaA8x58CeKcbCPExXhC62eR+p2FjKKt2oxENUumSm1vFHW0kfzlQvMorkl
XYhUglJCLbDJDzx/ok7RNgAvlEonFrV2Nv3cxpZnVZTbc5r08JGfFa9UfgZMyPWHGyg8D+Bdtz1Y
iknprsIVjTkdORZaXkfjMQ8ZlU4rhVrpNOkJTkx+03IKstGShxsMktfeM80XQwtzAATShZ4Z4w4J
h7Af3dIkh3RJZAkZPDn+qbz7SsKtSp1sd9u5qCdoivZtUlRpPlHVCnkvEqAKtwwnKx5kY3sLsY89
S5HS+jqMSgcdp5c6U+vkg7zJuQpB1Br1xMmvNJcdOZVZewBZyrUqa0v+dQmGnGW256EDX/UwtEBJ
YNr4ZVs2RJ053E+xCHP/KMdQ9ovi+VnTH5DaQhDN7vcZ7ja32HAAMV0Y57FW/SW0fvNpY9lXzyfe
s11bH/7uKjeOMW8ItYgfsW9mWqBb1SN7Dwzx9ab0aUYlnsmlhdd2GjHj3LLmHMyiFf++2Kc2ushz
l5DwWged+drJxwbDE4zJH01LQVFKdoquYuUDcij86p74Y52HsmYgQWaqnvaqx622tmBtC/EQJ4KY
ZGW7rILT8Aand7yuFC8hkp7Ha58AZvI4MqmnBI/jHlTNxu2dbNpadHq7S9XU39N8+Wluyo9VSNK7
j6hp3q8hP/1O65j6bLFIz7nB9uahDA9iXyNgGAzQEd0yxKF/I6TzLS98xPh4ojykC5a0WTepqewb
d4Wkq4ATf/l0pdrJWsXOkOrV1jCtXEh06Y03+t2ocHFm3iRxDaU46XJExpsSLz+Puu6q9LXwqybc
iH4Ehl6N04rysk0HSmsTO/jCqYpW7kzQWNEYpnUJ+hW0P3scQKy3NPbGOBy36HFQhJwpS3KX7Ejo
2WrN7gl/d3KWmCJwCr7vWXwqrXuGSBSvHgDrsuIQh5Iojsbmbe2RUwqwSE+BbuRIRsbJgmeK63BQ
QKir+c3ziO3LvIG4yzvmJOS72hI5d/GbgXcHGdcSz2ibFqymP1ev4etkIbtMakzZ8IjSFej6ETGv
ubVni7zTZBbVknW/ujt9qofQMLliMQ0BNjlU759ZbU5z+7aVUD7LNvd1iSnzvizDoNP6stB4RP1U
YEenBnw248FlKOibrpZDPGNaxfe+HjuBG8ufCbsNoySKhl14zGDQ0DIuk/WGUA7GqHiafy7KQwp0
SDtKBQax53HXrqlx/yTtY/muLr/nLjYxz4G8SRzGqQyfK7fbBE+43pdTCH5aWm4QfeB5v5/bPXjV
tAQ5iPvW+XaY5HuJK+EmnJtfr5qeoCq8fvMSugaWNLLb+2MtSmfjp7PgnQPep35KkDFknfG37ZKY
ZtX7sn/0NLbwuuGYvlNU3VzdYbghr1qLoiPRTzyd1IGa7E8pCulY6P3gz55BPFkHFz17co27NqX8
Zu6JHB1YgXbBuPaPiIULk3B1Jh4ib8K1BwqyF4AVpSaI33mWvvv7G5fmzhSAg4xYR98igiJPNotP
xMUcNir3D4mqbfZIqSvBo5vGYBtoIQWKHU7cVVG1MOcFWH2AvkyJdpgFuTDazjgoVToAQ1i5Imaj
v6M105kjuRJqwgVHkNOK3euE+I3nQ8RjJGKBOlznfFGKWoCh6bFK1fFepeEXW4F6cGkhyHPpzpQz
C2Tm2Ilw5z5DAirED5y1DqZNX+EciKawhGpOXgcMXy3bF9lfZcyfhrF202TDhhFTY/NIMVkbUIUP
mzLcwA+lLZ4TmGuDxQD+WKjukiJ2TGJd3IOgUIZ3/0Umtr5MnQ16cncKfpiDZLV+CfJE+bYYFVDD
bmne0DuWjwbZRBzDb1imEYf0VA3Rzysq96qpyoLGuUUOfS5lyRZAS+9+eEB4BPiJei+OGk5RMvgE
PTMfol07WCaUkniXu6+WeVYm6iwhiI+++ZqTKNq9W2LiqOJOLRnITcMmzgkXJuwfaj8Mt4IB0Lfg
x5vsYuDWqwuyiEb+4M5goi54BpEhJE/GopJ5zIax9IJhxz8eSaakVqiv58VmPr2CqcBFUDCxLT/9
/iWbB8bTUlCa41r6PKs+HjvRbkY8qrKp26hsfkZumBECx8pZTVoziXaYMbviHQ+5gtzUqeEdyors
E5Lqeyqehg8LbshvNlK2Q9adKGnllL6UuYWFu9yrMHIuwQf89pOq30zpDs+2gNrqjgRnPKf7svar
DHPA+bHBhOWwW8rUtjj40ZDvjVrdFDAXd9UOaeE4qXgYarksrM1F3yVsyukmuEOfRnS9P8Io1+Yw
H8piPJ9VnLzQH9scNspr1ffABEByd2BVtmv5ixC1MEiUcALKjnHS3BgLIge2cILWA9QLtgjsPYFT
Pcagv8zgBHX8rxQLF9NtVNDRjbGKpHzZ+Lx7V6O2tFQ7hoWGom/sb8Wf+5vIZE4coFmFIhW+D/T1
8WcHELi7OWWyF/RsKwi4lWm7r5ODdV5kjUZ0i09ARhVEGundDy9nUCjFUF10J9UKVm1mh244Fg/h
Gj77mnd47kDA4dp4ILu6YnEfxlKkfgWafuy1r3ftc2XwN7Tn3lQIMFmlgPZP6J+XVFIrotOta19M
P3gd0gaxrA9wYNPcAZqJcoMtVoxHbPVqAO+cE/yF6y3HLURm5Q2agYamKAGrrggY2TQKTQs2eogu
up5Xuhl0YTLw12YF0Kj1bVqEgOXmOKZkHdprgvS+npBD7yyMeUM0FcRYNsM2NO134Xt+nJ8zDvBg
E2bYrZkC9wgRr5hdmOXgBW9f+C/ysgrcDvErVxOZlZtY41+0OyX75ZzxNngtTD2ALdLc/XefTwAb
qeTB4IlMjqcNNXjlbKECVfu2uIIw0/RNqgOkJ83atdSIy1N1DTSpD0DRlkorugf09qsBtaMWKOUu
y0/cYHim/7H+4WnSDoyfUqhLsKXK348v5/LEWADQVS+RT7AfR9JdZyYACG10cguSjFxQ8CCD8aM4
53jfBYc1fwR1jQbWI6a6Os3E4QpFTdvjTr33RfpEz3fe22hdmnRBy5CO2tNuOfZ0bj516ZBa/PHR
/AZi1crnjEVjVx72FkHkrgUoVlBe3UnVPGqIJVBGvlVI7+KGwJXFmTSL3Fmzkn78GrzUuld2xWB0
4n0/JA65txbRwZFimakiUhun9TI6Ssmf5h6i6LWhlcMTYuc3+eY/XDOKyf0RXNnrrcLJo1j7nyg/
qwmLHGIOVbeVAg8wkrUPVXX6k42T0sn5ezd6GlJTMnJMuiSrugb7ILa74Q4MW1e8QOEPE1czuKma
LqEPcXC6BFQ2In3mCiV5X0duZmsnXMO9CD32xaFBuLvPg9GcO+BwxzDXIfZwM4LeAd5OvR3O315O
a8khII6OpweprKVJcl6lX8orgLiUlqWzVgNz4azpcTxrBplYIgKbf0aoC7Znj/WGztdcLPzxe3x3
4NxBPD556oSDg9MRbtcTEbHba5jxJXE5m9lQczSYhkEKcM4sWedwcggi7ZRLZUI3OzgL8mlBnsuI
9Xfa6Ub+lu7Sv+mTcbShcEWm9797vp+kKGMe82a3zK696mA3gVMYQg7K1jqmp3NUex9wa/AsjMuC
hJHmNCIhh04fIZrbC2rz8kXvK4x1vUfB2EV7hLyN16rcWhB76ZOnF1SxCXtSAwpFTz45QtWCyrC/
miicfTysVsnTflDB41e4RYldk1PB4K/qqBKKktHoT+Gom582CEPjxTYwPaAT/1f3yPsaf8tFOfGy
8a9Sluu98U4A7Ax7fFw/Xhui41mDYFD+6tb4/OlCqQTQaIC4cdhO0+O0ICWLG8NXheP4lXRFgJ5v
bZRwJAqcgqXYJtF3OR1I/itNnzoqnd14sC9G49MMllrFzgRj6Q2M7E5BS4paQTFIk1FQIWnz+kEK
P3mbGeYYSfj1EISMgiZ9A0XKmqz0jU00qOvQYMLWQ++VsaqUqTujJtezkPHOHPQI4JsVIzzUmaaT
TtgNtne+e8Z4qKyahOluuG5wLk2H/WVmYAH/t9xXWp5wPSBhZ7exvrGdgw9iorN++QmTdRNj+dQj
5THr6n95AfVUA8f17Sxa05+3IAoEObzaSxwpaMYee6tJVrbo9x2HmAfmpv8VuShkF8DsRBw9nmd3
FuwJJdaQJFRgTvMy7aPskRoEl9f9Iz8qjb7Joz6s9mmQRZ7+eHCaXYhgJWATVy8lqnNnTHb/E7Ij
MNkSn7YNvuviWlvmh79LDogyKj0U0w7zkihj9lmlKyFdCrhbkpm3z09o1ySI+8zGT1XVbK6slIrM
ZrtiP3OM2tN9w22G3M2+Gqb6eS3JRnNckhTo7LCvtpys8xjx3w+pa02UAtAnpoGvjVHC6UAscNjo
uL2/0iqg8viCSw4A93WupZB0Y4texw0tEJ8er9SLvL7didLxFCkhPILppVoNEdPWKBI0/oef/OoP
+1L75A9LUQ8FTOP5q0PmZOBI0CYf7ELONsDrgLCkDCiiZ3i45smUg42kXyrw73W9P/BfPbeQ5oXh
iJEf5KNlXXtlpY2NjNFz72NBDIDqNmBOOuOwWlVvA6VUp83naonKQmOmE7k+9AW3fAa84Ltxno+k
IAcb1HOAtNXNT4ROD1q4NZPqp8vE/u1BfMWR2wjr3UdfXnKc5gg1D0ZOkfyC4UQ0F4aAuqMgXOwp
nF2/TBTQlxDgiiLOHW7NDUIGwqa9WhS5O6HOwSISF110ssZk0el/HUMHsWFLLEsciMfWoSiR2LZC
cVtkLK6NfUhOOplIudBn8oiWlnO1xcLgewPqiv8/hrEFPDV08PHjj7xV6JTSpkADg3o8MFdECOGh
aiI+1Om3HAgXN3W5J6F7P2/HTyT2u+KnH3XPm+FGic1C1mRsgLNpV53mS6IpLQL/XPSx3YD9TlFX
06XtsF1NeVILKwe3sSkgC/COP+a5F45/7HsSXOWLkhknQr4twyZHtvLtYBXNK3QSt2T1QvYEx/+a
2+2u1zlvJthDEDvLuTmsUst948gVhTul144xrWqPCg0eNrB83Yv/ntdrpslqcJEqgyHqlUQOebMQ
xDKndb/fgXKqIzosi48IlXP4xSuPiE36AmLpgOq/qmVTDQDgE4dPWYROFyAFmDaj04ob2l2a6YVP
g5n8v/jJ/hhChxrE8WWdY/hoADD8upG/nN7ug82SEBMj6zGOrvAFhwb/zTF33gvx0NGlT0n8kc5Y
4jjdCbNTEHD/ulKZGQe/XMKeRARj4uIv6CaWBU6eifuGsXCifKBoyVHepQbojZF2FAGHFsxTSKhE
DHBMeje81Ximq4KpA6iUqe6IXWPAM7NtYTJiE8FzZOhDzwEJtMVJ8zxda0+DhBKaFMh6/OKICMya
Hg4QXHMjxffqp3FWqYi0bzVZ9rMKto9qvICK9PoyWCqby/WmP07q0g5T7gHJ8HVS8vjT56ejGvt4
9RqMnkNwpRW6RZ1uYhq1jltNpKK1xrAqd4M4VBYItWYdYyi69UzXO2NkFwK7YJZORzBmVbUQmmbS
BIloqWeTHFT6O0+mgzN8ij1+EAPzOMxYBneomO6Bq3U6iIJueZefQouK8OCmLGmU/JUESJ0AdhNA
UW/wrNUdu9LDfBlS/4iPVJOWSOh2nW2S4rwQVttLjb5Aq3rZP/N0x3yu9g656orJVqIwaPn06e1d
X1iqRviezXyfNXjYlCkbMD1ALE9qMomFbpo8B5cfPShUJEh8HQAseQNWyBx6K0IVbxVthBibNqH4
tBXKMe2LRZgNDqaTyF9BU5RXorxwGpSorBJZaP3nIIe7WQ9C3XNfRaEUlU0qb0VLanR/6nvzswK5
n9zMZz9Su7Dq8svf/vc3K4Z9cHoeEZ/hREd5hRdAO0EX3ZINAPubLl7vLPa3XiTCJIu+c4e8rnP/
XeIP1InVVtNd7zohNzndEXBbsPZS9Nff/SrwhbXmUKSgIS8JngFs7I57DHMHlUnvcNb4xiCFz37C
TbE3Eg1Ai5+yRK/ks5q2m9W7+hOG/T4F8/0L/u2dKJeLMR57isia9ee4qC7TV1U9k5M7INF2lznQ
Jm/pvCHl8ONZh2viRjPfU3vja/uTic8a/CUrU+HBJ4bm4wJLu9JVBAQaj+M6KlDdmfPj5vkLMlRx
toWOfuOrMj6Q1InSgfW4cHCKDHrQbVPxZt5OZ4XYco6cNQ13nJOr+uWXYm6lz+961kzDvcdK29TL
TuojLhpm0ppBJZxRUmiH0JC64AERgErPOhBr4IftuQlp/b5dnTuyyVmQncoaWmhLCdik+ZX0Cp4J
tq7a01CHQjSm5S7ApYDfrlKDbqCT6K0osUg0WaD8bnXxhpztR2WVI4UF3OzO2Pb9OmJgM87wbzfV
n4rXZpZzUSTwdGk4TtlGNpL4oE2vIG04btqt1gPso8BnkH8gm6dBH+NHgRApo3124hGQhMo1R6qm
8XcKlmHfb73C+FLrrBfEeUlryyZnO29Jiw0eV35Gy50xVO0JLrrwjxMDCYDyvKqRuGjFKkqdstyF
WXt851yYpMcAPFOLDIkQagJXMtgEszlDqOxiBSQpJMJ6nt7qVgn/G2vX05RcDUaRW1ZaoE96H0ZU
w8HzVsbvp37wd+u/VuHSTHzP4HvFyT7iUk/yB+QQiWHGAGfyCaLgUrW5VEZ4jiRP7fCAXO6NlC0L
gbRvisBDzgyZqm5IkcenXSYEW4mI/qbXHxRVOPLQlVZhvC3ytDzIa8ET5gXWeMKCDyhoRceUYueS
6ADHjFPgjaGXXQHJNCW5CAHu1LapMdoGGgMQmx1GE9Invh0FrjRPzcRfKSHAEvj3+1RngOiSlLfF
Dq7/x5E5r9otN1UdinC4izJYmr0zxG4AbDeIjm2QB5FIBzeKIM/J+pTX5EOSYV1weVG5dscR6Uhp
W629d8JVZgdVo2yp5wLk9NdtcQcdqwJyQ9uXXqCVyT1Rh6TTIuAzjs7OsOeXaknp0/nf1p3gz7HO
v7d/l12qmqwh77j6WgLf3wUvwRqvdYCGsxS0BpjuUPU+XPF2xgPDmd44T1Rt8l0lZWsGoafIIWRM
St0aUIE9AIHclh4prCL8FxJ6v6ITCQHH17FHMqeE/XBxNMLtMzQT774RljlOHBYNjF0wJqwMWU28
4Ef0/b5castna8t94wc3xAwxGdbHG+wyly/9Bjbrli4jNEOXSvtdUz1jsbFtThHEKD7yASBhw73i
dhi08CPqg0NWrSrCDgETJSZ8glVJ7gj+qiUUBPpQMcZHoaV9hv6/T/+uDC2gyne2f936ktjcdCzR
QwXmd6TUJqIWYRq7Q3f/yc4/hmy9DRG3sbmShDKnp19eMdCcsxETBD8rMnSbZ6q8V+rr4aGC4J9d
OMIegCs9PbdPeWwDG/zWgbpUlNc//SfpSWcvfx7NmqFUji+u+jVpI0TTtAou05RflAMyfy87hfVL
SnFnlY/FbqW4wfoNZgPHbKQBMuwPbnVLKmamjPID7ftYXr2SR+2QO/DeOurJ3p7nLvN+BqjSruCL
fK0EEM1NThmxCLOMDQ9SSkqkYB0VnCUdBE4gT58vlxBIzVDLiEYhLyNJaEna8PgYMAvxx20WPT5m
wRUs+8kODhRDuYoyItdN1giQLXzaANQEgFoYklnMdokvbG/BL6dmMo3zqRNgj3qdy031HzetMTA1
h6fMkL/uqiVw9H64mgVqpAuK5/CktXULjcBC7Z58e111YgvrJ9VULCM7SXRg2dcymFR0MvKvy7YJ
Esyxc3tO4+YP00wE8B4Ac8DCiWivPfHuhs8mmyOjppZfryxgNuyzY+EgBX8uACRdcRRAK8iMvtGR
aRJ0Ae9d8r5drf49lFXV0K+JPIASP5NgtbS/PRmJaKMruQVTfwUDLtPTe83DHOaKVdElX1G7hwiu
Wkj1kOkVYT5rCVA6UrcpXywMKO4bE22RlPVn7TYO7TIUHOWy0r1dNUFgu0BduVb7OQPuhGxksIpQ
ZOptKTsCvdA8eBogoe6+9q77UIcU5I6MWsTQ/aNvzmuc3yW2NBNckR6BsIdbdrxI30Bp6z0zqbUE
JAUmCMzkjroBqKJYTYvPKLRpFzo+dECiG4MEjopJg1fLNhc0vxsP0T2D2pEZR4uo8NZINji18hYM
Ug7/PLQR+dGh/q3RM3AJrX+Zv6NEQEypGKtTmCsJ08Mm/FJKnchDGIg4vlIJl507nDqJYp9DmRbQ
n9s3Nou7BKlHkskQaaKmm6hrnw2UbpjpP8fhsFY7w+QCo8eXnHokL3eI2A7KI1PErGFfgWJiGrgj
wwHb8U7qByt93+wiQ3yy8U1BvoO9gVbjsX8Qd/cHB/7m2W133f6MajZvQnuCVvZKvzXONHh4WeeX
By1uTWHdH1aiUifWBDjPo/M1XdPVD62YSAnnqbqrqp2OsSVX/0HZvqzTi6QKbH70Xh+UiakAKSa3
uJlCABPxuf3LjOgKY4/nVVccUZCupGgg5CKfm5uoCOk64eYVC8EHvxCvEek7a8BQHPR0KHtRB3TR
bKqfpe7YnvubYcno05jEuAJTBBSQfnAia4LSSB1bjeJAPy3tenSK9NQRDFjwVHU1szGbW+6VPe/D
3A53WCOtSAq4o3VhswqB4dzznhgEQf27gdxZJhwL0pz97hGmKlgHuRpt12hi8PssjSH+e4K7H8cA
V5YnsR3zomTsK0gsud+bVhQsi/yN3mq/SJrnn067Mrn7iGAG/Rr9DZ0nH3CAv/8AL6vDkeUfJOiV
1GC4o7niTRM9Dy36sTSWCivxDardcdK0Ob68Ff0AnaiCu66GzWsSvTneBKxQFjfBGqxMp0OOzW/k
Ijv5CdWfz5HNqr28T6JXbLThtaaAnzlHA+xRz+UGt/JkLfH0aM+lOC5INzHsKiUU4Jgw/IELbJzI
dKQZEh2eHKr5OlObCdPihCIjoy5UCUsPQk9yLBZ8lmI+Bi2Qky3QNrGVQ6XGEweGVn1QEKv7UmEK
c/LJvne3QKnRIaGq0K+vuoOzlFTyTEao85YH3SzuaAsnoPvu9bN2pWmVg6BtZMe8ZlDMO8KaCFLP
0X9xB/7Rq/JXiYW6sQ0Sm27ir1G8RRHDE88cS8Mzc+ql6zmBk6knNYbUJi7sIn8OU1UeHcXx74Av
iRMhztX1mfiqiJsH4I11cpn5MbK68P8/GVlxx1UE37gm2kwlbAxjo1Hzs487xZ8/NDkFUmJh3qoC
AhQ4bz3zUdrTEdD+JkCABz+mp1n1nUhBZvXjSY8NZ40j1M1hzw77m41WHw1FUsXnkFW9H+QuXZw/
X8tTEiMSt7zWA9bdwnaQ3+L2SwDbmMyAwfkVZSpqiGsd78Moeuj504QVj+MYkfRdlr8X9meZObhE
EWhONaFS75PM1+PGxOSjqeZDtZLrqsBk9mRJwkwD9PLabZfnInihWwmPcNoz13o7F9wZNhdD9MtF
ACfIQZiH9CrKSGh9pILdj5fs8yW4lxpILojtTcddIJe7qenet59L7jKox6lnNm7DheJP+83Qf/KQ
o7xXF2LOhlZGuzH4oiDpDYz+LqDvzChjSPsEuOMkx1MOWbNau1N4mpf/cFITJY1hOZaCYmcOq/V5
uOFa1Y7AJ6XcqGn6pWcKJc8GQG0eEP8bzgLUndxpQ70v1k36yaI2W2895ws5MOkNzorBe+xZWaQU
rB0ECZPWyDgPCY7hDeQGE+8XajtL9O0lO3Xk6wBQkfqnTMS1om9lMnpgrWW9b9i+esE29faa0HuO
EHdyFUZ7Ba4mH/Upj0fhikQgNKGA9x+jptBbXX3NGAQlXrcMr/grWJNpHPrtidDfkOCj2fbL4YJ4
usfi6sScZb/Vk46Os9++MGg2CBBXU6HQTSEt0hJJkpDab5Fb2PYqfvFvMopoMmNvaPDcUhHhFJt7
XNI1wucJl3J3/Lmj6sKKN3KNcgbu7AVKood8dUFlL0EdyQzai0Lwr717jAwOQBrNBaoec4i+uuhL
ReWPox9b9UwjysBABkJYiDAVEaKbxIZgpjz4zLvb79R6pcJpWrRXwJ7rCkPigeFK7q1GARxPWZGp
Gn7OhRsAP2Oko58y4nAc1F9Lq81wQy0JdIc5mKa/evmzjZN3dzdQTw5wm9LunM0u4Z1d7nrb8XnM
eBBmQyt9CFeq2OkgjE8fumh949EIU6WoTdJLVWUHNkXwZk0HUxJHev1LT1KmHPtPljepv7hjE4rb
YjJhHeRp63RCXg+xmK96hK8YvDlTqi4fOEuqQfq8PfF6WOQu6sAO8Hu4yAApIStufOdxWaaOz8Mt
82akHoWxzOV2Cb/yst087K3x8l0tnvo7uM6Z+BLvxZPzklLKeFzj+qQnYb3tA1IebgrJgr3j+7S/
EVJjPDNSy4t3phAOqdqqgR24610FX6BDNJ2bv3RAIQ5TLmD+siYzaX2Bq64ED/pbB/BF1pK8tSDW
HQlNIWTBDAXme4X6LC9LYwogkNSgvjLbh+jCrcpKhwq6z+fhX03hKBKYvXTygE0anU4sH42Mc/sJ
YCppcgC+p2IjQn5A6ri7p9XyTAYl9otgrAmCEEjziyeH5bXbPj48O+eL6q40zfmFuuN4gkIbcveM
r7mM6ne0IOjJGXLMcW0dyvMa6UFYp7nQVysTn8LBY4HR8HSl4+or7hLjBKmNSCdKfC6lFHy/8AyZ
EFdufvlthN9p5gzFgKP1ulkW4rAQ0LZT9HEA8k3ZsqHB7YowH9TIF2zUAUx5aFRKJW5/LuG+GLpe
ObMcrgkZNfehYWiIHUCBiXRDluLvbqScvYTYwtDOeGurKWQf7rwq0p4CoLglxLSjIk5elsZ61kQm
4Q8gA7B1pScXcyPN2WQCIhMMXX3MYtlsWgaTDCS9lVVFylWIRdKgTfG8ukCa1sZBeuwhVHrgwzYd
/pSZaZHLkhLc1+D+BpBoYzVanLdSpXUr91OgCq13joLQ+w6E508i4IwofWEEPePs3RUTw6qZ+Idv
X17nPDzGS2HbN4cJmXuUYP8/dFXUw1ACTcMjMy44jEn18FZv2gpQH+6PlfS0WnSmdVPmoLV8hRNY
7/28+owL5zg8LzjlfLMbwy2yyUTmHXjvB0OS7GrNx5zNZCZfNkwQbK/4k+tIsVz8TPNFo4jMtVyb
SCsZqZ7gjoP49tPqsHOdyeLotuoJQxBAXGZMv/wnKfcrKfZcF1f9oEjIsq4e+gHgdU2RG13ZFq+N
CxJP5s0kinnpEtqI/i8snAxBr1fsvQP83lis+S3ZbUElwrgG/oXFVw0m6x+OsVik9PgItghOEBx8
pt2+6K5zcnClcjQXoN4jCKWhymp1zbqZ6jmR7lDqGj5GGFbr0WLjudByxQqcLhhj/TVO52G/h0tU
019GWKdsigMMMJ+GGsWcKPKFikFr1nVvakEol9qbtsPn3+gNQtZzsttVypiqXLs2yXkw5YHgHJuA
kjuI1uB9KZu4AWWtWef81OyuaiairkOTWdc8OiGx8TPY1dHC4OY/js/RO7jtxpWdkFu/7dahQLYz
ebm6Yf+SR0allKZeeuznjNfXH/iXzVhB1B0JK3d3xCzfjDPXB7kRxhLzs/n6QGF22KGjnk7aJ2xN
BZyWjsujUAdt4dCpLPZ5k8QYk7wfktly6j977QUwsQ31j7DJ1lFD1WuF3XZjTPQCH/kOUhTfGj5A
EOAkeNGE/LnRlduee/pASsOwKyfj4Dz+bAlA2ozKfqH0/uYFoS6E5pWkxpo+6KPEhkGqp84tNa+X
6fLYAiR3Y75Rj6t4loqVq8ERa4FhzdI2EPKvDpiV3ikli5babZky9oYf70TWI3iyG6j8I1+GxLto
ALUxLMO+PJT3esp1JkGX+mys7bRIrR2o/qX+/ngFSe48d70vZ4/WizLRNfYx0KUhZ43VORT6Vp0c
WGyLD4IYgMf41CKPq+n8vMpLV/IjeFF7ZU8Vblh40pZS68xm9s3GnLqMkkHK1gfH/Tb8pY10wrRO
j5J4BIraRXlO2JlM87exSjoN270/kBDKuV2u4nufKwAnhYwdHq8L5RKFP/ieQPvkYWE6gs23Q2N3
ymolcXPCamMj3WcxwspetXU+Y5+qppQz+PKH8Wa21GmavAsRPf0k72CzwXR2Y08A3qz0+qQZJxpk
4MLZrYA3L2aCVfXhYhrENjO1r1TkWc3A1k69d1x03u66ZBx3NNUinVb69llS/94dtgmd8vjXHA2P
fXCNjqYp4evmRjW+16n8EavHGYdEjSuhfrsgNOxbdW3+KvInu3RSBbtwEmnIs13bdooCki9aOpoH
WqpCischisyskOzTrP4GCZo6XcVFwwzfIXfy+pUKO10dbQj3qXAperlOQprlLEadXF7SrepIuZMZ
5XTrQAA3/OwTFSLmc3vgSuqTL3dce8m1QaN8/VacGRbheOpeXVTBlsMf/0hqczwWG/1ZZmaDJtOQ
1DCJoAiF3DvmcNhUu/XcaDLceJ2zeu7awV+S3lYK5tNTIkrtfM7r3oe+vnTnvTveypkimaA6XK8p
VUfYD8kQkipUk3WRmpQMwhM2SkWGumN1SvMJRgQfF/0paV5pwg3Ic5PhTLJz/FuKc3UzATRtf4/I
aSbGzVGQPbb6W72t9u52h2K+6Gyzr6/J7TCEJNxG0yLjOwGpzB65E+JDjgsuVTtXCTqU5DcAXXUU
mfgvCr/qBHWmdM+dqwILNC9Vs1bvGJBN1T6oeuyYEW+Vcp74rIPwMv/ORepedwzBsdWnAUDvdGcR
PAgK1LS8rCZ8wt7EmHJzmbsia5+tmoHRJJiwDwl2h7ed6FJerLZyIclt2eH/nZO678/09fdiNI61
uTYhYSlZc/Y9bXbJYYhFsA6hBvvugX10SfdE+KxrNUat0OdFvH2hAHAGqugPNfzcUDNx7P57ayqB
oUmja98OGoTfeYeCQApzb9GE9qBUa57faIUKklIqy2pZho1xhq86J0qo43CyGoIvYJBuycrmCGfz
D2CEftSioAYSkSxexMV9iNVO/DB9pWBXkHtYLZbDntt+yQgr/80WLqNVMe0xgRpZurARwUZZRJ0D
4u6l5zhITm7jHzAAW67IW1qfnK+uM7u6Q6ijluV1oDlLzmUu2fCD9LHFDwLQd8Q7bBQua6SQ1uaJ
PDhxz/l5xQiMkrIhxxAH2LZxi/1C5VqbO9NloYdGtuSnTRyMrGuPtkuJCBnTtyaPkVz8S8ijc3B7
ZBzi3cgEdYd4sVf9vQG0lQFTzFntvvmTdS4NLgGVWw4CVcTOfh1MufEFuoUktrPK/6XgxVRUe2VL
1S6kTggc9SupjhTm90d80slqO7kudpEpQS8CAdzTTlEApoy84C7z9DVaFGrKmUMuzEJyiftxfiVb
/g1QSLnZZzekHoZYc75L6POHw5/wQQ65Ovod6C6Cid4pfLyogn3ucy0wyKMQfJdUUHfkkwNhOU44
xPpBgDLIIvq5QIyA32A64PvdsJTtsluJkQ6WQ1fiJpWNB+pwsuabAlfrc0nu5uqgtXyj7Ik4YLQA
qelXzqXwIpiWd/Rmv2l1rkWNGPigHWOKlKGabWxZdNKbbS9zIq1ZJ4NPb/eUnb2O8BP5SIFNZ9/2
9wvW0b8JClKX5tFXSD2qM5b4xNIvebkmZR48BmvjFWRu3rzlCDfgH+M/nbodXmbrVsX52vk7RWBN
b/+xdhmo7SoS5KSjKg4IMpATTUqtMt5AYHFSuBHD50Bj38zqDZF2GGIZR2a6FcrJvhVNVpSNCX0C
yQPsgjvyneoyvrbZUwdP3ffw2RWSq2H12L1TnN2LpTnsY/5LUzUspbluc/lRET2gAHQtEMEjM9bq
kEmwbac76SNQzLTJQEmfxEUcVVY/dXk1LJKjwETtwX90Bhsn4GplHkw8L9b6E/57A0NW4PLZ+3nw
gEqziLlaYVweT3KHMdKuV7TyvKfrjQ45JrZclD5+ATMvLsN/6XiqJVCKcVxyYZ4TIabudOPWKYac
TbhJ6MdUuBqHpXxxi4ymUWOB+NqxewRcx4jpZK3Vgj6Z/RLnzvwj4Cg50Pp3ZvE6DU2VTODtlRME
OD4qCUG108fEKG5LvAlD/GwsWfEPqomuFfzJXpnINo2IjtO0x5FmpPbVlWLju7e5cRzSEEYXQSgW
+6/ipw4e6sQMANMVs4G/8CFIP5B2nkvT6NOoKfQbxAvEgSWZopjTRMmkE9Uo2xtgiBJ2g9lKQGFd
LlZ5CgqTobuOZDYk3Xwy4xTTj4Jrro7D7sVsXTR7TNH75gRSbGjbfdCgCiuknkajbSVx8X+C1qwz
EBTBEuVmRTM73neqLRte5c1cu9LV0e5HgqYPXO/4KL8dwPv4pXnX9KhW43epSf0Ko8BIY/XsAlWU
zBN6h9BLzh6z1j0/0khJrcxsqqsmtYMWObVrL3kP/6ywpeDCpl6g0Rtpi8AwdS+fvu2hIO98ckVn
q/zGRoZKtWvWJD8Bpk0I8Z/DzQntSOqchBNKdkWKuqo+WMfokrShM6nH2p15DI3aaSgcfqjs9Bm4
2LeodkQAcBI6rTrqmknlWu41PCSUDm24FxNJywqUZXQ5mMA/iAyx1yptw75yiS/Df9tg3rcjKeBa
Vrn8oZeOCHSYUWoRSzjKYNDXuFaoE1y0tdUtsScALvgAFVdUQmuJUKkNDgeA3lP/kU600ugefZju
PXYJt26nkvMRfkuvSwBBw8ZepDOx+upOLkI735sN8puk2pBsNjM96QW4hTJJyQQxPvoUotHK8UJB
4nuqtLQFjHhkWWbVBNaj4f13b8a+1Ph+3B1RUMbLVuKnRvNZ4aTSYS4TaCg5u/5BaicTge33yeIJ
kP/l2Man15F7qodAs3NMamPXVpkXiBGU6eGiLZ/UjFbNKHUkFpvz4Y8GOZgDEQcqjiPdfiMVDyuC
2XruqkjrGDpOAjzX6gejb42OuBvZN7/HwXmzDye/ZEUdD8nfyreo/DvAylAZCJ4M+m+UFih/hWoZ
HEn7YNddq9QSnZdG44C/6yb7GTE4++sExxQMysrsg8P1CAiI5W7EBYPSZPr2t8RwcG6+BgV5rCOv
lLS+kDKDdESiE14QHpBF44O4RRb+m4JPqTIf0SDpfETdQrW5rhvNoi/MeA9TE6vtTR8xUVA6L6lM
TSjxnhybqjNPGKUVUgC1MYi2KcQlmI4jSk1/EUdRydMo1eKosWzaVPB4sfcalNNzugiyi4gGhYoe
p1jOgPuxlFa3Hsz2PfT4HgRL1NeEyOxHXe+APQRA9r3lSOeCdXk3mOTIPlnyu3fA7DgkPC0kB3n0
e4pqJ5EdiPp4IH9TyvUYQAJEkTVeNKceGEUTzcqb5u06Sj5nudEtbGuncYmgflFDtuR8DCnrYjej
j26GnN03s2G6avIM2BnJsMLaELMFl4OHBzTSU3HjG+rir4t6e6GC+cL38L0YXAGmb785TszSTo+s
HEO5vS29hJutb3a4UOSPCK6BX74ikjGhoxMhFeVJRQveabVpAc7oG7dAEUmPKaMo1NTmx24LV/UK
/v76vOAgEk4r0JyzD21Wl9rstS86Y2Zc9ui6K3Svetoh3dmS+2mS4Gs+Y0sU8xuj9MbePuSjDTSW
o4tpLOw9K/h8/qR5E72eGuOyT73BKPLJAu39onbyVkfd+R8rySsE2JmkLfjsTYHnkCQ3vzKVjQy+
kDNspwB7MI8fVPTbk2xzwMpX2vx03Yjj9Pjqh43ssXMCnrTEJBvKrRMSz9yAdbbAsXnosMRbPgBu
nfJcE3vWqciwCfuJf7cjuAWaLaVhJ8wGbOCsF56fuumbaGwdCOkx9+CmPS2HiuzBDd5FnR9HQtLA
GDvyuUKqWS2jQwa1EM+rClnr0yWiJzJfXOq8QAxQ4bFPGJcIDGX387ktbwdPVVerSOH6V5yLewus
gwT+JL0tPlVfYTm9mIDRNiAf4pfQjsIv9zKPXIqgHmRXoYfycCIUpC/52uh/o9ZsnoNMYCTHxUAm
jc3E9AcUHunMCNUAaoxRmjug+QGYc2GU+4WF5MZk/y7i+HvZN8mlSeE0g5tJs5JBs6cvxqGTZflU
zY4RN3ryhAMcaDimVlx5uj35RCjLUNMr0N7SXnzL4OWiiu0Ymfk+gwWtWR5OTAiPe5P7YEKWbPQw
Eden0dNIs2+GQhSNYKZNbsMm6pQ3ST1aXUvduo5fGUu9rwwY5ROJumBe6ja6XoBqEXzm5ivkG+Xt
WCFIpVffGPx0bh2tHK/y+qTOPliE/YkJhQAIwr3NKusUmRzsfxXDj37Wns0NOD2uvhbnGwa6z0Yd
ZV1CoRDPjO9d1O20g2uYdrdD7iMpQYfWjraIXonZba+5SlRlafUInICXc/QI0l3jm2fgHc5LbgCx
ybiG7y7IFz1K8GrqOqNXAJGuRWDjk0k5r/MwAQVCfIt0lEo6svsLgjV1kTD+8Almhx4xN2HMf9it
bSTWqi2Kn+GLnKwjVXBVNB6pz/SQUwN/Iv1gkA0J9hakAXa4RFbtTRYZN3Ah0Tvl8a8sgAswV663
42WZ+e3dyeHzI4dsgp/okQBg8jAIfjgyt9avb3K+NLQ5Wrr6cRutBseTnKmWMgOwI7HUsA4we8lQ
ViDVZuWKWGv0+R+txyRzWG63EeKrEgJ6dGNN+YVu9m5nyvpyze3fp7Vcqeo6H/23/DeCoXcK6to3
91QpsXESxiDSWh+wrcMCXmkMxhX/I3TbTJBTX46weFaV7AmgF3EqTZs6Xdc8kP9mWMxzRq6nhZlo
aL0mKxyQkQ7uMYDDcRH5ShId7Cu5ohTYNviBsvUNmuUOrdJXt32N1rpTFY6jh3bF54fjz7eYsElX
u/9vFnerjd9Kc+FP7vJPnACbJDXJX73izwDDynGQftW/7grziVYhU/wJJasuiRrrTiLo3FTPISjY
Eu7sTVBvvhXqAVSHUt9AxakR3Me85WVaIxBmQ8KANog39LZIvYi47OjRzZYzR3ttE54goAG1ihfY
fGpDYA+5t3w5AmbXZQipW6+r/ciz+4RLa54JJucgB+JiMsU1NIE/z18GGJqtZ9dh3ELiBnNJ79G4
PYRD6nJg+27f3kyEW/JHHgYRV97CNU0f9sxQ2xJFkIottYppvfGith3bGHHMak8d49WQ16n5oS8f
r4/kHjn5xdqbjWHCr3XXAONWd1BjXHzD5Amr6u+lWQpqLO22ldctLN6x/YKqwbzXuREuMhAtJhtC
8uJ8bkKJni+FpWOcmbwTd2zJ6lz7zaIl/1W2tsaB+wq0ioO30i6rjBM9YWbMtt6eB3LwDKhQID+O
j1PQ1TsSgUKFiM5z3OUbrq7MP0F9GRG8+JmayMpdHjWN5R8/zy8+kHmfB6sf5/b3rngUeNHQq7VZ
lTKv8xC7nYoGYnWR2FR/hnWQVJzW4cq2mCsK8aCRf2dnUGqh2OHbHGeFMLzU3hj/5AyucnVaVNFn
UmfJN7Rcx+QkhdySEe/E6sT0c67QQkwAfgEOV7jHl7ac3Uyt/BUBPVV+LXBfkxcwPAqRLi4csrh9
4pI5Ajs6UtWScx9ZfUEbHspI8E7mQGGLc1ixQ1W7hOzzPZgQLIbF9zJuTAgl14ijQqIqnfqYZpTI
EHaOslhdErRsRT8sr4OPkzKemS3JOD8WDLmA3b4tV/fGEZegOCb7qgeRR316UOz/pOcrJbsalpKx
Y9XBiPka37/6BuIe3kqtrRbRDVgZhqSKo7OYb2lojWFEBl8ZLp/YISS/fGJVg2bIMQl4Lgj9pNq5
ryP/JGiqZma+GH6JdUlrW5Hnv2CIlwGzeJMu2nEWPAMiXe2mKvY78+Nbw7imdWv292+Y7lsC/DkN
XsuZOlFLnXcM1Z98F4B4Z/DTs+n05gc8WQRxHG9ZHOPoB5AGvXhsS+2LjtwEY54N570j5IuAtGcx
XxGFOC/Na1XOmRWbW3UyXp+6280Nwe653mk7rdRa3eUdBmH0hkNfq/bkVXc+foh41SzrM/j8ukBp
qHbtDH/ZAGtWa0fHiO2BHi3B/nRx33QFFipRIoF5M18GST9IWBSTd5YiCOTFVFKzYtZSjM8Tm2rX
CkHj3NDhPWzKBAMjazw85yK0VEgcU5rfoPNJa3a1MERlHDLEzvq0WKvHvEGH6cmLUCUNDEJZCdb1
aeS7JW3RaqlHr2eHFE69eFFJ0hVa0VYqZtQescXGxZS7t9Yi3jUgrxtnP6Awabgv6bPdFRQZsqW/
PJWDqg2f5942psxNj04FDHMnrJ+6sUDd0H8xaYjc8IstAvwnRVp9u/APnlCTHoF5u2437zS945MZ
kitPtWtxzWzV8IEKjCONd5S8v62RtdrEfyq1cayYo7ZQUNgT6gjI494ORVuoSgb5b6nSOZpyBz3D
kLMaQh7VkPPUZ3Fq2qlJVt6tWO9nJFW4LqPYFxgnDLUvsa60BwvHQ1D93NvZaXyOu6mYVZRl2AAV
h1U+dhqoMClp7QfX8KZGx7QnyyIDlEPD7xIBInpXX7LpPMJJckzuNQiTLU3Q3B4wEYC6+nGH+Zgj
PEskCmtRw9IzMJBM7h7pOPJb3KCdS9tWAwZTXJnTpAW0JaNfzfkVsTRWyFV5D7iNoe/EzkkqwCjB
1mmsbMBlYtX0A2/5hZBvVrK/UkG50cjVVYz69hZSHsCDf5VrN7bJ/2Y/A/mAoHYmq7c+d7zekQxp
TdX2fvYxHadW41Gcm/mTiFEU90LOchO/3j1mi193e5MkToLJ8znfTKo5FQmY6JrNvYuA3mx8ViFT
1cKR3F8ZymlVO7XfiHjWwS4aB4o8w692IOgRpb6Iogh2DkEUyqOtW7xctVotqwWXm0jcPyV0p/ch
eQDw2gIgAz/VnOOFZwL11cHcR78Jvt1Oe7IXDmmAHpOzJ8dUyfEheLzYWmDCq82n9hR6MlJy7b8r
l2A3ih528I2AIOyeUeQLe33jdXphRGDg2ZkTV9d4sQ5vF0X1IFHm/+1z4kqKhBOE4DlqMmNdif2q
MRRxk1hGZXhvNo5gsdZF1jOlo76OpaDpAXQiev2AyZ0EqZqpY5S37bYwyLdkzgDeUmeH5Bq/2CpC
oY8x9/2uwmdt6+28lA3hJEv4xvO+H9NROBHeZzXCShr8Ftyb/6+wg1g7H9MHtLwSUlBwB/1WOYNt
4DNz8n26pXHYtzlBFXkKOE/qE5D3k2wgccElVrU/kgNTgd5kYxFu863VUmH3BeWhwVdVQWoyYLVn
wJ06ogolEjpQtGHXyhGOVnWQRgax1X0OPCLOFO6Yrmj3zlZRciSH2V6gVkAWBILBjQJCNq81alIr
n91lD2UKK4uXgADLGh7XNvazpnzrJGJ5e6x5SWfXC38cAaGiQx25fSRfGvH/bXi+PF21E0XmCIzy
01fjCDpSOHK9RFBluAuXrTOG5OTq18pxRh6JMKI2I1rq+8l6CB7oQLA4snJYICv5ei4Nes+OB2jD
Vw7ff5WavQPM2EXcuiNXUBxvEMi00dnhg3er545KO5I4YegyihsZxjw1DrrVWMnZr2pXNz4k6ycy
Fij2BSSMinAojJrR0GFBtI9F071+GFcko6hWTMOE35FwIwzlCXkkE4UVGcSUkQbe3XLCkg9hf/tR
IPMMWb8tqzUvy7oqxSyueBKIIAsi1sRqRjfmnVTrJP8uT1owN5HfhZhw0DZJ4xpQ5bQGTRolFCp5
bsaNHR16Z87JNDT5xD/MH+lDEacylf6bucD0137WeyjhWH/HNMwKoNixUx1nczA1Dv+mjAgMmLBd
5FwZo0z2VJKRw61CyD29rOjsRVaXG0un+PxR7ObdQTQf2N1yeVI4KYIC3At4lY2UCKOY63oVZ/2Y
H1ek6PtsqiCrs9kSyP7UXm3/Wk6j1bksEE+m1zu9y4IhBs5J81J7nukxF33zLgUVATi5L1ami8YG
YNl474NbpKpGCRDbskV2KL7Ay4/V/gIjlJNs0qvktHxVGcN/i01TsmhOLG4iVif8HcsuhlV9MKQU
Po+Xmn4dSgg/SIOmNdGe31eWl7f/qXMGdPUWCxvTdHnFEdPIJLAFLMgIhAls0JYRdHKDi9bYKsG5
17WK4yhEZsjOzx8EUfz9FWo9mdtwilNLeosjURBmauCGjfKejDMoUKK6+kTwh3Rn4ME2aZZXN8AH
LyT6ci9sXQA4KVIEv94vAWYvVjJdENnuXzZb3CzhuCClVL4EUBBCALpEB7c0VzbP4VtBxvfW6hmD
cRlGOWCEZdLOVgna681gXqFvmNe3/Ad8Y1oIs+Qp8LW75j70xq7/nmeIvxBQpz2kHvsicU0MUqq8
f0ASccTuj7K8twgrQ2ozh+Qzacxxi8n8bGdE1HQZ2iVZqEJpG0f0smWynXOjzjbZYfxrR3NvP9tu
ktymNkBhLP+7xjRcsUI4tmsWjLmqWqsIiOx3iSkmR2ckS/nvfjvGBZDK22bRTxtks1DjLvTvl5Sq
GiqauJKEHZuTARrDhaXHYOO2tc1Xqo8RhNMXBh+8CkemDLHp7jFMFn5gtu/OH/loHWTcfx6rZPY+
r8r296i9JG3qoQN0+P6bpvGILKcegoozq7Ie3SihXLCoQY64Gkq87D+IV1sRvrSW+MnNcWx0CzKj
XWy1EI3S6DeDb67uZWz08Woct1wEpReriPZLk/1+xNgIGALhpLY4gVCKt9TT2rE9DJa3KLOgNY3R
szvXokP9bYYKRZHZe6bN67IgK7p55FKp4vqFByfdsMw+DNlOeYsuPY1WiDD4vbK0dpajuLRrFpoJ
1++i//HtxeOG3tyFO0V72qPZi23HTaMSbjuNQggZTbD90C8hmim4dkFvwc2AKWvixd4jcJgmcJUA
SfffN7x1ypir5q6c0sD4F1eYtF/tErNgIvbmaj8aQv/cZQ7cgOu4YTtYrsY9AXGN/KWPdKfMscKk
nkQDdzpP7suBYqtD+ol4g+MQU3Y8C+u/AORpfyszwBLWSycn8NZlJ2Qr3kgEpo88qXHmGJGAZ41p
KZ7VGG4enP5aHVGmnF5M2cQ8OQe6GkjJQDoLUU4hkV5gDVWVhG8JWKlnSKzLrFh6B+VWekRLfUvh
foFbGiyMh39zgm1D5zjMyD2bxVIfnGgeeigECzazIZsu0Baz+kkbnzSbReWvwpxEKVMX8F6hq26h
/RPVLyXz/J75TlC2ESc0bzsex9YWRRl7y6xna350DZEn42WOGUhJWUsX14RPsP8RQbkqfkrGD0Wf
59SG67jO8CqYt2UeOOfidaww2eXAnVSRZQ0na7Da0N3ubvTGknRRVle/SW1Izuur4Eb71U6oxxW8
7OsIPKOzDU1SfyS/CxjmUprGLp22kjmo3BaYoHYW3q0/2FecSHT56dujQcthu3AtZflDjRaFEmrZ
lpMztcqXZ69q7kjei7lHJZyd3VqjDUEHm8RU+pcontCn89EnW3kHjjFmn3IA3wmOVwqCF/V/7n1w
FE56O1vmuNsGWOaKpwsMs+kh5b+kP3DjhPpBsqCpoYhL9LvbvcHYpocl0QrzY+TbRKH5q/ENOCY3
6kmfKdPUStDGgs0dAPZfPvAKF5ul0xPgezt29ivprd2+ZtoPzikcuhK/zRdqjcWojJdhZFDVVJHQ
4l8x+N8JXdYo0EhdjfR+1gUGIoM4Xf1L4JYaSxzHxLseILIT/qTZFRuJmlOHA9epzEwxARh/Ib6s
D+bKMHSt92VEXE69dH4BC9Cco3t5lkR/8mvFSzMhehcihor1h8fJ7jn9uNhRHf+nqCzhGdpQaM2f
pmqv2nr8tPj6pxYK1axFsFDYZmyDWC6KDDdmLN6wHijrVWJV18zVDsoEhKwVIIE0SJ56Fgl3xOFC
DKBqwq7YDhQS59mKGYz1ua84j4jSc1+t62hAPVLOJQp4moV+xNf1h4P3V9dIHAR+CiUE8ZVtZkzb
TbHmm4ffLYROmZoXn1v6bfY2+MvDXnq9dRBTsbXrVbrhf+3sB2Pe0Sh7e22R8opUehx/WC3f4Gqv
YpOK4E0CmZ5GI3qpckfbsJSbN0z4k6REdeMu2JdzcFg/uEs5jjjwiCCt+0K4V7QhGmseWBU/3+rZ
wXBa6oaMEsIfpg491I3Jbloxpay6PYbDHO6xlwTPzmfYRSlRMN3fltMH37mO7Ld5Pm8lhLmdYN6k
nwX3wjtUwI5QK6kLARmsxWdehnC7RpVJNHJ/jEoMjuVb9dFz4jjuWCImvSAr4r3nleOx7lMxeYpv
AyZOPbgi1jDJIX6+O5HGuY9sKcGclgltEBUNFeCAgK0rKX3+URX9uzN1SPdrB+V6IHHEd+E3OrgN
L6T80TXTCFp4fW3fcEJNuqAG5mj0K5HwAKjwa4CcGStbdWekR8y7lBhk33q/WFl5gGkEXAkxh3C2
pB+hSS03HWjpQ+wx6sup8Tdp9SQpHDIWE0k0CjoU4AXu8QUEuHDgNcxgtP8u48CqQk8AL/lBKlyF
PubbR2ApXjVGfIb05Kj7pAqm4YxEUhVJ9u6psHVa6Ut5/W/zR576hQkv/H6AYAgZIsa+S+qn3g+c
pSXu/V6p3syfLabYBDd7bkahJ3cb0urzFP6SGDBVa5Eujc9UGQQ1paJsVOmnPfAjTCvsyf7czEOA
K2iJdBvQd6jLd4vBTu9mX/8dBEKDv9wYOy/yY+ItumsLiVbxHZ8TzUxeTTFgv8fGF7IB48yB1PqS
JkMN9M6cbcAEDjfQE8nCvnNqncbE7T+OphMLPdScanNgmBnjrRnt6EZ1bkV4pZe/sO2ti+sKU5kx
WmYUbZgJ/pgXA4/L4mDVNRqeQ7MeVh/k6ExcCkJtmR7XnYai21MItnPf4rVDAdrnB/XYnjpkF0Oj
sz3y+IVTAOEI2T84D0v9Vf1zwk5ruEYt+U2Lh4JqVpJbxd9kJ4mJrvZ8YVBhXRS2kDVLBIPVEY20
bNrhV03qbQMqeVhYLbYptLZ5YfJ0W6m9qeOuq1xmwvYLTiBBPlIgQk4XbcvFiXyt0tbf63x3FHD/
4/KRmjeOKo+iql5h0EMpLbxR2BFwA39A4NaeLFznVNdQrwhdoN+9jE2sqgBNjetRXGCVpSqFZUk2
pMtfMGNLFOjVTHYnUuf7+d6zpKww0olJbG9K2dJqw3CzRt/T1aMAXopCqF/KeDvneeP6GkXe5Wk2
qyncaEUz8m+DbsZi7lkIm2iugKchxKFpCJUzgD0KIClMmIVgTQAUag2CfTL4S0+Swba1y2zCR02s
IOIq22EUT43Bw3TE0k/XIFYSAuUJWZlQRyESbKgAMewBBm0LvOT06jJcW12SnaYW8hGLhkYsWyyC
9NZzZUY9QKGh/zc5cgYzndh4fy8ji55eb9NS3fU0ueWUn8KIIuaajUEPyWG7rLgrszHIIPPNB7ks
cg0MJDk3Aa//iiXhrw0t4X1EbtO+yFwyfy4rhOE2J+DptWoQJKWQsJ9jdV0Jdt6qxeCAZIdH3vgD
WeSAGswfd6sDCKxxcu2UxzuNzrmGujp0L+vO+VwAZFzzpE0dSkurtfc3d9IyhciSWb1ZXkvlpCvM
pVjKc8NoWufQBN3ec/a4MEfXOkT+KbMdJ2WT//jSYp28Km1yA6wWxQAbBgAD/YN8GeuYtk08YJW4
6qQMkuvSXUsstfMSecWNzQspJxs1klH91AOYOzuQW2aaR80r4AjLJe/X4NHcPBKR+XaXZfDqTwgH
m0qvaBDfwbEc6BWuIp9MLKiNVIg36DAMgj8pG+/NSAFYINq+fWnoM3hv0+FIs8GN0Y8V9thx0DU3
PuSTxKFZ0sRxrZhGLk9PMKs3x0KXDb7tJEWBGi6TiSWOn3eQmicqPITJ1aarURypU7PDEUltzEAK
gP2yVkVlKKDNa5pdxIt5xcJMXf2O7rTz5vnVEYYgKJCDSuQTN7pjTasea+dVFFwTVYvRtft/oRp/
md/hc38lojVemg9upJHs9MXWd1V+9HdHLW3d9YShgH1NgwkbCqDd6pxDHuZdq0k1wocU3WdguDxK
+P3j+b4N3GIsTno7PGF5Zt0EGQi9MDgU8kC5LompXdks6+p9nRsJ/dKSM1Ef8PSUPctv0Xm7e7o/
YvxnvPqLX0wgJhQsqcEBAxFwfnUaGaJSP+TGyPc7mbt3vJzIQubwmKCW5wni49sc6kHHitqsYSN1
KpKnI/ogu6WuW6OICoowcAVdmJyw2cjGnUyHDHXMwB9OLnzyyiLLjrLkrkRGibua6DDtOUiRleU+
wRhgwxjD04V+lMkWl6/j+tB74CGgof8pVohgfezACwssAGnK7jW1PaeIKRLvSmng/aisMz006Q5/
N78OzVVhf0B33A4hvfQGYIP3XSlwdebICUx7eiSJoNW4lhzXCqx3OxCfEJfAaQLx0gBJVxeRXef8
XbkndJnF7XOjzPLF860VEnumGG8F/CIK2yHCckd5w+oncbv1YLjkgnSUyKTOYitn+pL7LS0i1wYL
hBuevxmian7W4d9h3llU0eHLQhrHBir0pNnFk1WYM4z+b/u/sPZon7btVDP6W0Os8wBrAahml3AP
EPpXbmjONDSeDz7SE40zh5w1RaPgkYacy8G5LyAqUdQufpd0bTBjlTkNeHcaUoyGCts0fv8S4/OB
Rll2+7ho+CmO08Q4VYbqEnZ3vbrZEun/Degy5Xny66i1iy7Cv0kuQul41ejwDFiBDDHA8L9sJkg2
OoiVbi0hgQzmIQ0n29yVp08m/3oXBEsPPBDJLIruRmbpydJaPIePEXEHbT6TsaxGbt0tG6iR4gAJ
4icPjz1oujhl5ADN8hnPNMgRM/BY6Lr5a77cRWLGwp1jSSLul1b6LDnY2aVuBOFNPURss90jXjQT
LFISZaxI8hCbT/iS4Ui0fIGlCdvTXjVTXlUf03/67zUnu0IszJGmw0AOhn+h1HC5LqU5MJDa9T4d
2k5vR6fwh1tKSdBCinI4wPrbOBi4BFZwcWdFM3iuvc6UFLRdNpaYyvSJZIdWL/ePRMnJ7TUTeF54
LBlTQ5Z5/BK2MeLXQpdpg/C/YVX8W+c+YaNf9QfczBMNG9XAH/VNYUdUoFk+yspnc2b8DtsCBb81
O6u8sdf805UPmZW0OKCrzyqN8I+ZeeBXwqA0dMNS+9Hx/PE9GKhJ1/xLrzdiL1bEXOmes+JOm1gI
S2gWW7j4gNsqtROZeAMfalhVqyWNTStRUCB3XIHWYyouPlhDjoj+iJLWuXN9QvBFByNso3q17Xt/
W/OnQB4Mm56v4DzewKaiI30NErP0AuGPjSKtb/FwBc3LIROJ4QQrzJrXX1QnMb5ur48C6qkItwa1
vVj6VphwlTD8QydqMvC+vSBAC/b5gMIEjm4uq6cMAWNEAxWd9OPPqF4KILND7bJorIwTgdbXLzce
zbbWmTwvM6Ow8uHhrOFoqX/s85N9pSFfVwnyLqh2nyZzMgyMNrY00fMCp3j56fFCaxMROgl6jD9O
dE/K7ork1NxC3ONc999J39uEfsHAgpw+INErgJlIvAM8RWVtvaS19fSUG4IDg0pnWb59gO27KR4A
ValGrkfp1zn5EqbKoXXcmZuTGkThsWlaBmoEqC53YPo7G3y8fSgOPdAPsMwDF2nXd+YCIqE2fduy
L5Jm/Pnjl0202KkA+yJcSldLf8/hyoZAkKvVPWEx6gaSV5ZfO9LVDpUbIo7m7jEjpSFgiKGjKsMy
0cyYlCcOhDOpv1AJiLG/pToOfdGdIl+LCrzANGtUvjr7ag+Eju0za3dM8XZZdFQsdhZ7LGNQvYV9
uO9n7p6Sd1MYDljxq8D2/rjQnlx1mLj4VRDuxTHNM+aJMJjJBVCuZWfMIM4OEBHpiTKvwkONoZfD
ToSkVYHubHsYBdkFlTW7fx/heG69uF44I2KCsiP4RBhNZRbVq1FdinPaaiwlHHS0Za8pWMQWu/Tt
i4SfooQFVOQL49jw3p+dQ0v96NC8z9NmiRLiqnBXY21jUR08+FB1J2AJKhscSOxUnlcapwYluNn/
X+CLP0qUEIyjucnAttzZTlBWUjyrVwlmgHpZHxnn6j9geiNrh8l1zlI2qnhNCcoaXUyYS17SScDy
xoJ9Wme6X/qPuK5M5wLYeiBdfW6MCKQjCUHLI7t6BagJacAN315MnW8+Fe+Re5pVrVnJ3jvMG96O
V8rOyGQehHAJQN61+9hrGKB/pEB3R4kACVl3MlE+ldxmFoEP2ytDzaLwWZMLyb9QWDhx3YlBkh2X
Lx2lSWtWEjLxymtPySreuGNhWuilV4du+oGsq2jcr+EGhJOUWL5y4PEo1ZSj1e38AA5n5+AiysE5
vKHCEi5aXpZ6CCgDwvfg71XI0PgTRLrwsSx9rQKA+CxJGkXAe3B0U6EX3shjuS42LZ5a2sl2blsm
6pkOyRd1AjvcABRIjRWFM3kGmOSMv8cr4HfXmbOfXSwGzDjDvymWb6hf3lC4PgR2hfHazJfQ91uT
pqYawybbRBdTAFoeiKQ407MmJiN9H3FH6EwNClDoaiHidpaXxnP0pb5HHiNEPBKO/NuP1Z/WTFHk
7cqCmmp8pjwfOnRifEC5DvD7+GIEI0ZxNacXKqSc4LRwJy+kOGdF1s32TWQiIm76wca7cJ+xGEW9
agFOi9VHnbCW+U/Xe7+sM4gKphtWsrnGaTd4vdc7IwCRTBaCvGgly1YPgreyC8cj0l4F2458nRXR
IdyU8R7ga06Qu7Oxc4RykIebg1BDzGAnRwSpn1H9uc6IbVBWxa9fGK4UO5j/pQ6pmu6MI9ADI+cL
XpJoV+on6OcK9TuZada5Dk3Q1WjgTi57uKcEoUcFvKUacvMaZ1PMZKG0Jebm6XdWnduHN0hUq0qg
EqlFJfawOP77P4tkKVhkjlvTSI5RaDvHFELLEAqGE9YTCBW/f4OVooWFd3tFljFiYZlofRSl0uHR
ubmbiy7QhivtHkogAZb2CtB2LC4SqQJrnKW3qTWVNkM6/pQSZtuV+6NgwlaTmAAo77BII6ZvMRyX
qfMfTNkbPWmDzzxAkavQvSX5z33Yxu21ci8o7hwElwCz6NpcH/SF45vpnLmJremvquXx79PCQlWX
CxkmrQpqysecr60EIqOv9yMFsCCgzzJUZLoY1uBG0ur1SyiIlzwf/Ce5B0Kdp6qPp5uXpUrc3MRS
6J9hxsRAJ0cVHxyNc0pvsdd46WIwt1XG2mmREehZqb4etqCQhBD32zKItR3Pg8tIPkt5U1YNKpWq
BzryRgg1eQhkYVEQbpkblHfdfrB1RIaENiKY6mGxaUkZd2yQrM5Mc/W7qjHC/2lBlpFgSsaIEmW+
As7LVYxT2ewmVGGhDLQHaNPzJe1iAk7XzP9Uko2isgb3xyTDGk98ChfRQBpWRH6o9H1yiQdK59oo
Do6+vlZxVP8EMFgOvLavcJwAJN32HH9mSAi90KpRvfofhTsEZIiW+65J3lrq3XiJOern5iIjAE8u
XVaZ7yw0cI5cWkVfWzJUyKcR63cGNl7Nn2IqZXe/EiKxl1f4wvyWDw48IA7/ibEjrnQA3LW3FSp9
CKuxdBm13H6R59oD5YkRkfTW6XqTpAdq9/OPy29Mc2TOCGX/n5GaOrMvSuZphbNWivZ/7QXlJsZC
BVxNtzKpJMVbI80O6O4nqfE+8D0KVi+WIHKO0KB+HWT+ND6YfrJ1lcdsymJHnJAvaezJ8U+7zBax
hXpzgC0j30zAO4Hcu+HP8ao6o65Ce5ZCJyueicN3vopV/hjhoJmB980+oQucV58jAGMCYzC9UrCt
vE3ZG5Dp3JXNa0uc8gRFXi2dxG22fPGDo53/tS0r0aopV4q+Do+h3S2kHwmmivmAmTPG7I1WowVb
0rPqqCB4jcFHEBs4qFtpc+XgECvmlQW6VL0SSLwrf/M7QQd9CPMcsQRaV+kyluRW8ZA1TqFbyDKd
Cd34/ScaHY9qKPNOyc9slBs/aLeVbu1nS4wCl6r4UuyRm8jNsZ0drREN9m1w9TkBFi/8G796L2YH
h06F/TnPNoP1ltg52YLcDhdGD4vXgUm42VJszitqZfvzWMJtv5BeYK09DFiMQonQYeDo77gb0Ob3
Vk/zDcERXTXZJbxwefSQdvX4YLVztod0JkPMMsT9gv3pyWgBSoLPRDKJgxjKZdyR53nwL3FfVAPG
YYsov6iUu9hXpDPFqFMQ0TiyELW6v5qEos84xYGhMPXReMzHiu5vbmy/mgpt1B7PcnTN3XPLsJ/7
R9uewTqsNUDZvz/BorpWHP102SMdFmU2KGXTHzs3BmbmvJmBnETYKMGKbhOx5rhoDmEwzrD4bBoQ
xJuKhyIh9sbm4OmB8MD+B/Hwj5cFMqg90zMWWyc1m25mGPlqCbe+NtfwvfgCTxX0G5fiS3lhLeYW
r2OKzoZEeerXgOjjtVL3IxLL+JiCzpL5/flSsM/t28IH8cLwzBIBmFm4AdV0uMzpDSFW1x0FFFwb
3GduvwtT5mMmXDX9U5UTkBBEABXxhMgAnRkHZQqgQtJdA2uvnsZv203fjTkXSPs4eixdkHAXS813
wo3R1BwMPCnnTRdqyp3kglnHdbFXK15c7W2M1x5Afl4+ZlGl5JdOVBS4kCMD3mdwwNUUAauS34KC
KatoQEMPij6Eg8qBq6bzFYhG6wu/ogqkpqf75Z56iOwT0LD8eAGdo1hKxDz6rYWiV5v1NKmaUnVM
7a/1LpvSJ4qHqKhUoAOmAxjS/gm2sFyF3Rd5mP0MmL4xOxTTl4AKdPROwQWWdha7sj29G1hm2EXQ
DpayNfR4lasdQ+XGCFxNjYnvH1ZHpJ/aJpwItKxGhh1SN8Ea81q/X+2Pp0DxQSseMJdeBZqhNMok
wf/07m6LiuBpjU/+PC2suj5jQADDSa8HVUZHyLjW2nuqIaCZqbrXAIcom7Umb1ujaUb1x7tDmrOG
ybiUFHRDF7Ljex8PNfrpdTmDixhS1bWTLYNcQdIlck0he7NPB81T4bF1XyL+u2VjsMHS7nv3bMlY
jOA02M2Q0VeOdyRP5A+ECYwWs2nmgmv/xXB80mrl1aNR0yUDARUdJsT09BKDErtd8lCPZbt4wVRK
QBBOWrQU8yOPNZZ8vp3Z5Oq5msxh3sZg/ovDIT2VFarFmIwQ8HhsHt2mzfVZHatdAJOHdbdASMSK
GRUI6yLxYXYVCxvz19rBD4uLjD6+EFI6oKLG016DQX/AX00OD0CNmJFT0AxyUAy0RIDGr0tE8niJ
ghNnRBg9f4txZk50uMVHbGi6uNtGFFU25Itbnti0aDBfdsd0YqOWfPfm1Z6pqPEqA8hXv4Te84xM
IMOBPO4lz6JiXg4Mi838mDrLdzYR7SHEH1h3dZEZBjudmLF6drXhgSjVICZ3P40IBMJYXyYsIIBn
rzkNKBPfQb0EnIuYRnV2TpdqQYBCvfzf3N1kGigM0gYv77EiU1VKOLAiL56JB84cIjL/NSGO50AG
0SWyhpQ+qT2UcvWb+k24sMSvN3ys2km6DW/K1aa69wuXtVnyTuss3IwZP9tov0VND9R6XBCvTWqL
YxVeK6qf8i8yzFacSy9EJxuKCoDHIe1Uo1fD5jF+m1S0QaRJbktfeaQI+gz29n0IbDltVo9KlG0T
cbBWxr7Pu5Oi9DKNM4k85IhJ896qnuCFKMhccTqhRB/OI/xmKMpX9T+z51a+4uKF2X6/dKluWTco
wYRmCqbf+ZxqWxQC1VIA3AP7wjnfPKkhNK0OAZ29evpgsmL+UCO6HLxxIeRFYZNVxrxPMgPI6Y4f
HJprcEesBqO6F7ssEVt5XrMCbrKx6twhII1l/39hFB9SRPS7D1jLw+tPoberuAwwSEAQMFaXChiZ
hFdRvKik/nL1ZlEKEFEc9KWNPNU0Y/bJrsEmOa3AhHi8sq8YrgQAA3/4PQRzcHKmaHMqOSCPuCwh
xX470qZ+DjuFuh93Ny1B++CVXirO1N4dE08WWmTjIVyTgiOZcllkbRGeG0Rl9ypCvdi9/iTmWkpv
ZmXhSDXb9BcEH0WkDzfgua4d2n9mst8cT+AWs1K4Osoz5+Ta1pMkOWvF87ig3hndSHaGH8ylG36V
XoFOghoQtca4xiwUalSity0sgIdpfgGjrY3EC5zKDk4Qr90nDE9U3rUJPNeWRJMmxoqe52GQ4b82
k6+NvJDdR4Is4LsBDOtZN8hS5kJBYhki2dzYuPCvhvoGLsBoKTDsYc4GWFM/+bVHZDrR1vwz2f4O
Ta/Jj3tCRyK7dDt+jEc5tWA03Hm2sn5MMMH5fmuYL8kFAv4GQy0XRFwdYXhJEoZdJF6jDI/xtAju
h5mRPMIz8+fLJuZX2nHyiBKw87Lk/abSCDJ5ZS5mwlIT9kDt4hjAYR/1Y3QG0G8HTlSPiqc+2nm2
aYPmBDn3Fm8TMf+exEoCjmc2mCKRvw4cPBZZugZb86NzcNg/xhBP8gbEFT3y2IaVziQvLFHcC3fh
I9cmeDiUEwFPLuM/J+JBdrl6bPLUnqDRkJHpK+CS3/S6BnrIEqZ83dIAo31cnSTq8VbPQtluudpY
fvJtq5+yJR2dBQjf24tgYIUVKlDPqpkuPwDFObg131a/l5Aj/gSAN0E2AxRB9WnhJDBLotYFYjQ4
uReCIVjkEwMaydA6KGWgXkT5sC3TTLSQYTviPdgvgvSY6vZBSjS1+UkEl8zUPAQgI7n4tayCeBDI
pJgkEQwGpWohtcBGlp/dFsaBO5pR86XFK6zLkL2NH5nZfqizkG7pPIWjlNE0kyVmcewkYrDFEebn
GSwtiIFPO7AoOzX3I0d4Q3q71fh8XL/wuf8/hYjZRHD08s7QaMvDktk72+hbuizbbzoCXOhfk7M7
naNQcUIeobYUCXGKXxE6I+yDrmAkZJIqAFxgwf7gsbrnlmVB+oGkERrCaZsZbsNdBesJGWyKBuwr
BMKIDVE67Aq9iUkriSTZf+qZ6aiI3gvMZN5Lyi9mrRKFc8ex3MUL1VC3IHYSxQ97LPrBV6u//0rt
9gBF6d7pqSeNA7sUWL46VsPZu6hJqEH8BVdprs/TL4W/ujmo7oKYUlgpaUjNbNNByHisT9hkTON+
aXzDJ/aax5HV0kNyZ/z7GcBez7csSHQ4likCO+pGn6CUlIm0kgse95+uEKD8nboI0PJBtmEBg6Wc
fQIobi5BaTBIi9P7A9M2O3ersGQZKfRGzp2lg4pxENc/rNPL/nYxTCciMsw0KnjnfUyF3D0KprZ5
6Edh2nFnGfLKs0upsYtOSLhpQW3NMdqJFnirdfihmDuyR4Dbf5pT+QyOxapDwdmZprbTnXZutv0p
7AMpVh/et0CnYOpK6Mx7R5nUwK1n/rClnyVw5QBJJ+h+T643j8pbLTaXCgtM9R/Xtvr3YMVAWn59
C9RvFzqDmeqRkSUQc405wRg5+zkhtKx3Xfe9HKwJydfG9ihycvePq9ZxGjfHf0oXnuMKg7a3wIlI
5tGpjPZ/TWlxKrn1fdhQRIbIrh43o9v/6cO//4a6uCu6kOmF06eg36+J+lLTz58AnAmPk1yLb0LS
SYSjuNk6vlVkWfg4I94ME4/VOA6vTXshBV0U6n/hr1aLl2IariRkvDmpicXxB9qFfD2HNevfV88i
I8ZEnO+p30EmxI50G4nSMfIhzaf4KYKYlbhI5T8EVpewEJsCBu/IZyUGiZe5hDOEB+9anahim4d9
yo4oTtFaJNz7eyqTTVycHPqBpgPlE+OmmJ4g7/aC+t534/jOzQbX10xwx4sz+npC0PHS43+jFg3e
+poFswQBI/aGcz5fZcAG6OS7Ejn7QofKygUpTAc+SWfVhlYYgGwyOX7TIHhHccnrd0zvJTuPlvId
G0+u12k/ZLC+SwA/IfK4xodND2Q1g2Y1m4tCQLYt8n+HS/rUrKZocHHIEz6xDQJKUzaNJFxRib/6
94TKiaw7yeGhhEYc3GPinMWgQPTHRKrE8QztbWj2Zky4QVVVdElFiaEZvd2vSY62eR9N6GkuAJPk
KK6qTwqkn7+xB61Zqb9tMbr/En/kYw6mrP/txhD0u9fT7SLMpbb7aGxhaPERfABrGA4fknms6tuA
USS+LYvJBaSdLWk9gjPkI02u4y0eSTzbYZKknrZlSQ7EESACoz5xSLJm596X0UjinpF+zKiIcT7Q
CrNoNjOsMGYDjnenA0CPg9gfPnTsKflGzYfHRpiuXH/I9ewUhT+p+zbtURstra1OHVjLVxmo21IX
CACRqv9jIqOfOmQui95bq/sOq2faEg3SaEMe7roKFtkxjVSe71dzG1iyqtXVljYWTvki+BKFChNH
LLk/FBQH+iqH/EdcHk0ZP5J508uqX6qLpky8ehD8ppviCZLiYxMlJ1xdwVmQ0//JOKs1Kj4F0dm+
lUyy2yEzcAJs7Sc60qHkVeQNvGSyzu79+22Z716m7Ip7rDBa0e663d9ioU4NSEd93d9QQZUt5USR
KH4K7gAVcOv6fm/i9i/gUN41aAe/ogDHq9K+Vp/C/Glw2Fhj+xQJNgiJk8zhQFdoEu1rKd+Gj+eh
PX4huR5E6regGn40WQLTe5Ru6wazSHfSL+JJVHQg7tXyr32TU01Hi64e/86omODLPWINk1UBWpzi
K/CdUfAJ7c1RuIPjPq/yxOmiexH6ITx7eNsjbzKe4Av/6iakgU2FnDshtUYD5ALic0Qc/s0tS6De
o6RGffOPPAqABbl7rUCkJDIJVIWB5hxpaxybkUWuPBWWVonb/sRpMNlseoPyveLL3Hpv43WEvDpW
xbawfWuv/WmTBt5RGlhfkaIRmITQZYu7p4JLbdTOaR9mcQq4ogylu2W8C9PezP5KptCl4W+ipWLD
oy8zRM4rVw0NtnZlo393S71gFRnmqh6aX9Tg4UawtXJNKSAUVJ3oZy8ppGnJGM6QH6lkLPuDPrlj
DM00KiDr2MqyAZW438si3/bZcluviKW5XGM4r9LK2Hwo9gAfY8mTdtUbTJf4bFlamLEWj/PnZCOm
eG48qvloulyeDTh3dIDCoDruG+4cTPhB1IRUyun6JKcdB58MnQdTQyGSYrj3fpRt9+hpnHzQqhjK
jYBxYiYN/xIuXszyZ8nonp8dX2IifqhjW4nui6ds1HP90eD+4sij6OX1pyoN2/+JtFc+GLKmGVq+
MEZzw0RH0mkD7HW2DJY83cYVWJTFOjsxlrofBZZj0AHaDRFfmdgRmu8BZ5f+YbHIX3bFYhOrLjcL
OV6e/EDvMYnGCV/vooAUu8P0Eq1qj+k6uhtviULuYK7i1AzRnhzTYglVUgOU617BN2jdrGvV1lTh
UyDn1muK7VZcNAui3xDjp/MfEkVncp9Ttq1KwFUeRO3zKXWku/1FZ7MBOlo6qBiVstU7ESQq/if+
MO+QQGzs/GI6tC63PzweXur6NAAJat7hPy8xuGc0g7QguZm/OKko1UmLVokDOG8cIYqhXS2cM6ht
SB54lO3NNuiEA/RhX3p5oLbDbgDV+aKkpxFW8mfOsSYAD319kE6MMS8F5JN5wOmrvnBUDXwjrCOL
wbIFEbMyz37zBjFTMSPVGxLUYW5LR9A2X0nJgVjS1zprnvAL05Uvz4pwCOOxW0eh0D2sQ1/Tal0t
SJeya6GYESi8GFb2JNwM5sa2iWwwKJD5yVrrgvmsbF31wvG0sr9YOIunqBEMZ2tyhYgRy4nfHrpT
a6VG6zbcjqSM3Oq8f745fSmrqC+7a9qYRk7IS8IWOXyyYDSlaWxSyumuwuBV99HiMTO489nfGm/+
3gmkM7D0aFEAE96w2ktD5+ukg7DdazcWsBuUFjEKjSh7Gj/L5PdsLdVuVHM/Ixm3Zy/eKf89w0/l
R6Ctu9RmqEC3ffTgZ3kclUNIHpXxLW8zoL85okaq/WaYY3gDO3nwt0WFrs7TdwP1xT4ACHUBnP47
DVy+fMqOX5mLiMQh88pvV2dOPGcHrQN79fKCsUm245jj2Jtj2ofCHneAoZ9nmnki5uhRvZCk2mAx
Y5wT1DHlnQpsncIDvoMhzcLRJwz6cB0s0twHgp3KHOkEIzjs8Dl8+pO4GMe3yJOV/cFA0GGVWMDY
i3bfMH1pvyjqPJobA/DAq2qV0J2zDyP6ASx3F0iS3JNKxS3VCOjoWPvvBPKgjpvbI9m9ekcO/dcs
2T41VdK5hlzkK94a+WrDoapLq5HMo4BoGVZByc2fQjw18UOQcgwzjJZwV9abT2wS5JGc3D2IYjrd
sAp2g7aNUp4daxmfGlkK7gokWZz5lS8P9YBK1gdDcEHq+F5F0xkgW8avENP84bcAUvVtxT6QjTTz
kAbzFuJwp/4Cd7UotLucKE4IKNt1pi3U5FKwIQx2KHAvDdQxg7GUcOtxx7+pwMhqfzfo0uM0Kjll
W2k20WB+EnJQb+2gY2wK1N2uBJ+x9yNsU0244HwG+4oQy14g3z8DShh+k9jV+TPAX39JQtxgIuMc
QEv1j+THOXGmBFxPMQx0zcfaPx/dDIO5d4AKsI7zbiF8gtNKKogC2Q7yX/+2xP9T3Nq4ycDj6z8s
qpNmStCAxqTPX6LfKMUMAyGDM5MQMwVdMQG2bAmQEZyQ5+7BqBlcHW2O9TOCdFUI6x3bymohGJCy
7PNj7TpJw909WKsMvjWbwdahLW3i7sl9reEQiQUEi5VhrlkzoZPbPW4PWI9Eo0QveTBUyaAEUFpe
RZ89x+WgTerYRKsT2r8Q1Ce8IjYStsgcH+nhyBGWxMTyo6LGYs/lukKAoVBiAzuz5vVguNJ2J/92
cVjzNNYc+9P5dZX4hcAx/c//58ATVIW3zrmlKc38P6ANRfbfHzinpSgOHgqGs7OLjNrd28TMasKi
Esa+vMZEXsMvog7AIg4Wxa18Ce9PXjzZFXDZ5TsYYreBkc6f3YHfap2p7Xcad/gpZCPBHAwMk5nG
UzMnZNscg3rRCIuuk74s6coyoaAZlQAht8/wjR0IxRE9MJMd3YnP3eYnS0Wc/DHvhLH9jh/75nUF
PDyuFBEnWig1XFa3SnGcQq8I1XqtPz/BZLVTXz0TRp8rA9mE8FGxcZbhOKgiYkuV+B6q3Fc+PAvE
9jr6NsQhzPKVqYik7tIpP2VXYfmXAvq2s1JoT9zh5fwkgYXCPovq3RQtQaZBaY4CeXbWsvzDPd8F
fV0zMw/FGli3V43jmXfnoK+XDZ1OLnF1fiVJbk5Bt+bCNXMW2UorScio4c8xEd8Q8DJsgA3s+uQX
xUlL7N/fvqa3gcX4lvgz5riPorkw9F9M01tp/mYtLCi233kh9ZMGQCs9K7mZHy2vw9mCAW3zqj2F
9egUjEOkc63C2zo3b9TmWSm0so6T+WbR0VjMu9dkxdMXhL6/ccMOEIWHQFnoPPyHTzl2/pbyG7hg
HM30G8OiUuQBQa6QSEd4ygjxabqmyanzEj56utRq0ZhJko3GJdwIxxbTl2UyW++4TLS6GzJ6yXj1
TF7qJaU3BE5MWpfqhPYnLFH+swDfJqE7QmOj6hp29TggNRMgbNctwhBvtY3Z5M0RhYkZzz4scwMu
Sh9pxCU/yzGgGtrUPnWxiZB+yf1AI6YmPc9lPxC4NQOMPYqZN+uqcCagAQJ+ddq217rugKb9flqB
XhWoYiuISYhoRIFIhTBvkitY91tIqGH00Tr6/LEhl9u320ZkVh2PA9OLI/7q6Dfn8NGE87MKWL3I
JJ8HZtiNAyMCwFIuH2tTND8EB6GYeAklVRhro4gYo3Ps5PveHJRzC2DvLBhwE+x1uqv0mW4uOH6h
L7kc1Fsx4xIwx611bpMjsSYltXFyHmR5mn+i4dk4FtJvEuu+Z7nDv7NVHHTYkC5STKr+wSRZJsZj
eLnlmlSsJGblmm7yegFDHxAT60gT/56Ph+4E5o2u3owvX1tuK4imkk8YoMI0GHVEr23E4HEzn0DI
GOZqKCTqLlzKlGI8vrWpwBY5Fo48gqLsDj/U1BqvtYVhi/c3KPUd39rlq5L4zYLBX606zVSKQ4ci
3pT1IUi2hMqfadvUSW9k9Qalft/G3QHEb2KLuZzW/JnFueW4Yx3L3FvRESxNkSh8ci8aBp9VEMqh
VK+BXwUoQnvhcqvwxl9gFbRbD0SHGGlJUv9CRpKyQ/XWLWNSKitTmd4prl9mVL+mgASD9CiArdWT
X3vBziwhO7gOYz7qkZO4/y06vJ9ehx42C8LOkNCLuSi/cGq9WNM3vmySlinE1dPlnpnGzUogZXuI
FrnWbnqGFSftJPEVrF9HVdoidW7PvdO4b8vn+MIil3+YRlUL5z3iZTgFSo92iTY5mxrruJ+XrgY8
nTTV7IDAPwAbEQG7CIsKG0fWaVZaZb6JKMU962X0J13Mqhfvv4IaLsCYjk08EpBiAZEK3T0Beh5k
+F4ntxP6typU96sOc6NlBrJtjQFmUMUXRKvPevNLVJ/5A+hPzYfYwUNzyxhz4w/zLoMbUycMzN5k
rEaYSIEveRC3s9wtu4vE2DjBHJDdeFUWAIsjwr/woyv5vr9BQq4rrSY7vIGGhv0g22pvV/o4AZMF
D2LIbH4ZGGN0sB7ibj1bvg8vw4YXVtTp5I0a1zocjW55kwO2gz0vLgkn4eCvoPohHLgKnk8U0Dzb
LmEk3r1JHopxrPlSYWuPhXQXvZWyeXC+fuT5bliP1z/dh+nUp5OJ/DnPMYpBwGF4pIGtKm/H6nFI
w+GLP6B4LuGZrlzGTgRSiDO0tlwQ+Flohy+A2ajQBdIHrdeiLx90i7IhBZ5WRfz+QlYadXGVvOh/
7seVBdNZDJqpXyLjyOw9Xv2vvP3xJL3F0gi4ZhGPjCD5B/GSAocZ/DbhkhRWtocVCWUuIxrj1dGw
BzwrrPhQIK0qeA3pmot+M51JzGIZKHH8qISkVXMDknMjU9f/omqe7i/ZJsrtl1iPJDOOVbQc5WYJ
N0sefyxA4774JCRVT+MKHf6T3A9plP2R4gEMn8rSYKUcpqb5Swb+lueDwk6LRQe5SrEWnzH527T5
9LsKu8sZ1nbfBxfTWz/GFwadybfCp1/Bmc7WXi9QjdBkaj066kxNSG1/cesSLeFGifRdEZQfDklx
LS7OfmryEHQk9seZqL5HaMxV3aDW+iceNozAJBuGyb2w0b+9qdpJZpNqnF+BS+bcnqBc0yRvEEG0
zekTuxMb8rocJLJg6coFvkhw4vdwI9XIcPbmrVAl2Cz66HiFFAj5W/Dn/OFtQUDYzzCsURH+vffC
cvWUDbsWKPVDxLUPoM71EtojqgJ3UFuaRLZzx0sgL9ZRrp+SWqSsx8CSn74M/6xsULFxX+GUvvLf
PvxxXSywPmLV8VYFv97Psqs1VILqw4oVWecLb1+febCXJjn6bV3jZm6HtQ2NFm9VlPQR6Y420k6Z
5CEQlnFghimh2S3RrYYguVJWsWGF/OQw1/MvVO/9FnE7lax+BH8QiqVcQR2Rau7TcVgMEQu0FAMy
twHK8Rj78ohdYggc/KhtXr1kOB3h9AJXiws/oyHAzq/CThh+P8URpSM+ifsX82s9rxQPFdcd0git
GJQ7tNRlCZgh1flLOgTWJGbtFpYbQKwpyWCFCf5cGDRo9YKjhKWynqP2/Kxljgiah3VXWs3O+1ia
3sqyHoN6ks9BEkoMMLWVzqrbwPiV42tg2A/6l21ZkyvEor1jhMBhTJ3hM8P8/GqZhGTur1pHlRii
/6pydvb0cTwgxIdHe4S8Ed3BQmiR2SPYW0TcXPX1XyEJU5jdxGaPn4ueyXIqdOhX2x/YRPMpwZMS
o2uxwCf+cRa6zm8+XFyC1mnCgVpUK9O0uvGUdz4AuiDmznrPhhTQGBLxQvMgnMwRo1nTAnAunhzU
W4WFySxQOO2i2s6awUzwvQc1Vv9SpJ2kA0A+n6nRB3lu8nFhENYJS7HSvLWOgDbpcOiFfBsyAzwx
N4GiPqhsBshnOonrvKlFxoPe/CgP8ul4hiVxzvKD96wq36I55bt1YXn9IxBkkeOgeYO/h69kzCrx
Nv6oA7IZRSYk+J8f/+07H/s7VGwGhrpPMeBzkRmWVtep3Olrwt+MkZH/V1bhfl0IU8r+UDBTdZGp
rPpWxROU3/sHVFA9xbLUAeBI2e2iDoVXFafdDZq/qSFYR1/EMK6UqlHYPRIQyqHqvvEot4hcCkD7
lbCrmXptuphVXBbBw1r14ShUyezWFx1amiEfJUBK0LZTzVJ10tQGPISy7H6QCRUt3QnuYgtH5+0W
Sm7yr2lXU4nDNII6flYC8xONkov/Q8sVN781DOYBFKRvR3o/6pJcN17+vO84lCTs4U4jm9bNPRJI
OuPmUN3fM0/6mLYNS0uslvPmqlwR1VuUYqqNGOaTY50Uif/ZXsinXOoWmdclAvWqOBsaaxdWGqDt
hkwQCtD13oT2K5yo9IvYSNg4+WoXRMEIe8K+WU4QmQjQXEuJJzIKAB0sy3e+o4A9j2c3Ktw19Xz1
AKu1c03x64p7FX+WcUCck0t/9KMNrFlYpHzL0CpdHnuR7t2r2EHo4dqDJEmnrLs02VD17ETyjsNy
RJORL6E5UVcuKMjZ1N3zUGfZmccU6Bohe27+9n9PDnWdFuFu6r7fg9ovrmHZv69KfAGI8QEiZ77x
9kmO92nvQs/EM+XIyzCfhQHv29oHGylQZfntSUGgFwkrQMWsNUOgXJrbxXOttPowzWlPwckLVmPk
tvn18hpmE3iYVwvbqnBSAliAwakJ4GltNCMZ9tUW5sQEclT5O1HZbn8tpnB4h4CuiVDTsCoJl+1F
fH7EZwdYZ/otgDDo52KQlJkSSJXFRKfpQ+pYp4cRjq10ckAtd5Kcca6MpAw6A+FZvvCRxDAYZu7E
DvgjRN2eA8DUuySWJARgJUWzxtIBHEjx1kYPmUW6h97tqdxbQEfioR64UHZdCWTVfs08KCphcSeX
uMrvvKRU7jy6lEM+n0jQkVuEJShErzvon3Mu70wuwPVJNkBWBSHGuXRqp6oeTK3DDPTRLZTvkWDR
ge1+mR+33LDG2FIOEXPdsryhcm17mwdAKdfba/VIVoA9uMsl10NvPkDDtggGJHVsFk7VVPFZV6HS
hbSfB3IZJBiirguFp3af/ZNw9Hg/S3WMtUvKMkCcUiayqDqjU4dMD8nDFhP21s4QVJIiqg+cE7gC
XCUgYMIOTHW4//cFKFjj8LnvIUa/XC6vKG16vCsZjU3PoqOSEMYCuxU+2wJOuWJJ1WkT9Dxzvkj6
GMd2sWbMaSe9oPsPq//4QPfXRIcDP39KBdrsF4eVjIwcylJepiflB+y8Mu6dWabD3PUVvfg8QZej
wXh6r/aUPfyHKoMyAEpHb5pzOVoUZH7h4E/wC1gQi4X3NCQg19lg23mdc9zWcnfKPTLJIL+cpBZ+
+5jfHI8BVo6Hi2MWPFR9jeelOX9ztG2zgSqnDo2j6+XoCBH+6NDNjFirNc6lEGr88LxFIkRKmGFX
jjTViOYsbu7qUytGyiCj+ovDPHmMsaaRBeyroGumZ+pDBJtoAwUJ1rMPQKu8IwBR4wBl4mbYyXgy
iS88W2XFo3/ZclNd0RcwGSS9o/mSulH6Op6SfK7exJ5SXMnhtDdm1HeFAHjGMqaAWZyER4or5nMf
5Nb/BqBHh3CzLyqwEMFPEF6toZpYgQZvnaAI7nqBNZ734EX8oZLFDVt7CCBxzOi2brLGNUXXPjg4
2cqvVFmTBEhOtYmgVweaVKW21a3JplQW3kOwGpdzhpVC8kP197q9CAVOHZHVjyIwmXGCmYX/HOnI
QK7Lp9rvl6cLYcn+T421ObAbFz4Ee3Sqmvde/VFO8lLRwPAy1C+HUbgsb5Rlkkr+x5YXuzAhyz3+
NCp2SMuR4AQ1UuYFY5ADW0cTQqSdHhtVZczHcVvAYLoZRKOrgYFOdCG0AbIeC1vGpx7YX7WUt7Le
1hwPgsp3DYReP5Lui1W+YsWWx5IX0t1cIZ64fBKw2Ae1fmgv45lDJQeMUpjDlIaphA5ZPK45l67+
j4miS8k0lnPbDbH8uh+ccyjDsVBj5tmJyA0L4DHu/jymDt0DkO9TprSv9sZJynDpQxa+dM1ErSHd
m9E5jypdn3jsbgxwvMaCCTpM09m/u9Ai/oXoH7/qBQ17ErOnGt9i7cL/EZ4Pv6yUHsT6vrO1qLC4
0Ekx2MRq0tiHjrYH2Bcf6lWwhqUsltVmRKQitw/YzzCy39PP6/t/DwJ9arcHtuCJe8kSP7q/VrBe
qv9kFSmE0AhIqY0Is2Lg8hX9UdmaXX4i3YP8QNPw12+gubgQkKe26n8kwhdJRW0GRR/B55lR7aaM
6ZFayKxb02WhQvyNTlIgS4717QyW77Nqv4y01td4X8THu1h2uZgxN3X06FW2yl3XD2PXUAGOBdCJ
asNvdmHzJ8yPtU2HvL26Dfa+Aepx2XFAV8MUnpDarla1sOhxxts0+2+94n9HrbrgW6R8EoGIbXNw
IwBkP5vNsoFdRGzdJTkVK3Y93d1wg73RTzllyy6Zh+rVDzWja/CCMMdF5uM8wTQJBxiKXqeFS/ji
qsyK9VnumyI6xYd4+wgDB1z9RO5iTSK91HLgWEb2fodFZVIQMZ9B5cfcPuWiI6kbsCkcbv7yfDn4
trxsMh7zAd4bcOtRRhAfgBOHPcT/N/W7/grltXG6Wx4E1sn67CZMMLw+LwBdKu8x33tjk8O0iiT1
dErFPHmMhu7Y8not4ynqfyti3x4l1OS/NlcDPskHhplEbbzym3X0Sp+A2Sw+0CrfYVvEcvuy3XjE
QpiYvrUPMccaqbg+SkPkjvgvZC/HQnizvksXyz1a6OtPBk2ejhhI/EBjd3nTHrtiy9ItWV0D6zgw
uTZ/YKJq+DOVSKufzdlLWQ3CPTKKKejHu4BTm62Cd9aj5MQAe3dKf++i1YbF2/p9sxR/hsU2q+Fa
641PfIwD9P8AZoVQbs35NcwBHH+auTMWNhBRBrIVWVYF+4fj4b0tsCs18KxT57sDiZb7k5GtutVC
Z19L5qUsE0R8K5m+HikwwG1mfN5wKblpLGBefYWtTyL4X/zW3Z0gn9wK38LqYQuCrY00AXidEvlX
GRsFQvgslUszXIdtT2mA+xODNAXLoCJ6c9UWtvpiNBtO5a5GrxINZY98g0Joa+PRcKzCUzvPQHIi
G+GTp9wd0v3kZcLIuWpnM4Im5Jn7FEAvJ4Qb0O12SYeRbXODdLWnqvNaJk9Mt4z46j2RUPwSYedo
IxjzZIIlJ+S1HQDFSGeNfztkLSvXyAOaYbayEeCXFjwwQw/IRqPiNcWJD7azLEdCYmCb9/oqIaZU
ug6mdE3PgATYfZ9kgUuN8lXqiAmGpBY1eSOCeXSF2s/3AQr/4ywhY4MYBJFr4kzjp948rnyy9QYG
4SIU44RXoe2+1rnKQqz/2Givaqqkhacta2YNbMbJQ39hTfNWa1plEhbHNNlPTu3rFQ4sK/7hJWwy
Yq8UOdzh1tydEGPDCRSD77fpPhAGjqG/99Aap0Q0FnTxDzdGuEXtlWyRoPNFdYbWDjTZWaDMUzKt
I70tAICbdVxu7J8Wi3rcCaPYXWicAGHStdu12+l+wwfnu/T9oPawIUiMgwq7L7e8gCmgQfAn64Vo
KYBAowbFT5F1vC9I9ijrHIbkhSspdumkbgFvfHGOuhUVGcwCNExjhu2ZD7kKEr8QzDqObRtVp1IE
lsnTw9+llRVsbKBYyuACtO98g9kde0tDuw0wa9A8I5o+YVkcM1MEuH5fSqDAUfqzZvkRlgHkmpR7
Eq0HFGTqift/myLUsbbo+GGHRxg2TUVPqBeZLgx8Lq3+JpqmQbyW4TjDYYY0QPnJEwvT4z10DWIL
ldCmqo1f1PnkEiJgXrYnRfVIFx5n9H1YnNGs9W6u/yKclxAQgixvjahyk9YWwk2SOk/ripMBLVe1
51xjONsPxi+gnDCSsFfezTg/Gpai3EGxrKlkYyguz36sw2fiIbqkvOwTT5b7ePXSqw6ThSiHOlWh
qn83tIMM9zkLYeVaEi2Bm7vVM6ESCRCjKx1y86T8VVPQlEg6lmX3OUiUkkQuVJTFItClDDOUuQXl
1B4MmapzL+Iz8K6hPXjUe4UNV2V2ODkkVEo31/ebhaIZRVcApiZAh88BhgmKMz2ZCQob33IpNe59
gI37+v/oa5N70HznGBCOBQNjkKNUxZz+v9nG3qxXHjm2tr4Qs4pD6jbLC1ZfrZdBXYThE+eBRr/w
0C+uAzNWk2dk1rjTPpsRqwxqiwimz38slo5UOSZrkNVOWsX2NSILU0j5P6CJhvFPxXcQs/qAfjH0
wPqlNvv8DKegyhwtj2UR14CVOOHs9ypmslIsQfpIA7LL4Toj+jQF6J18yXxxHRSN60uiQBvsFkXG
OqPCbLmCvocFkm0w01zN022EU2SFUMgmSabOUd3IhWbg3bpB8Cm4bPvXSkLSIjuvb50No5ikIsK4
UGHgH/HJxLW/FwOxJHiBcsyxYj84itc1Prq0UL7RTaJZwsVPoNSfvo6TuQmK6sw9D9wHwR1kXEKy
prdr8nXfbr0Xsh4/ykknV5DlVe73NfWe0tILdbWOyvZNmD+YPA7jafPlW8GdGb6US/b2NVVxzdZ/
UhObOG6glmZsLjVrnYJdwfW8D/b/VtINHzq1KL0mjTwvubsU96meOOQaGYkZanpAwpzV3zKAu2Wa
7kgAss6u1yCco0oG85tgYNPXpGws/iw8aUXj7eLHUX67lbDeFnoS1S8Q3izHhWXoicUQ8C6UwZo5
MO7ijUR7fZBD/UX7WzWiM4dCCa7mAF6TnTcmpuqHd4ZuVwG1go6U7c7/CmJOEzaHxUzT+Tqk6OaB
UeEFb4/3Ls0D353WP3WuTpfp+dwMvyIQWzUC1HdYNfp4/O4Dn7305xBaaahVSnXbC+mUT8+Mn2lg
4eppYZkUNR/akvrse3fFd+w2CqDzXpMJbrce1vxdMQbM4KbkX//EyVitIsAhDL94dOcYhaEyl1sr
SZsfst4YhAT73HQ3XgUyND+Wb4e05QNv5ip5d7j9rDypgEseit4DuX5yOOgIsziOabni8kRYQURR
pCHGhLP1Glyhcm4JDzYNzgWpsumnz6fVDzO62lFVLQnCfLK+MtKVIpEUnQtGS2er8qR44uQE4ADN
en+UqM/JHl97gxaDD6wQhgUW+QliutGNk5nVnEGk8MEfHQiCjxCQ1J1usSpciNhqjRuJS6eStRsl
oeVw+Vaz16j/tqWuRPeF2Z4xhu4EtZTyJ5nG55YJ9i/FbY9lkFXd57pzaLDP8eL5uKjlZNSOUOb1
6FLyA5v6IL+W/82WsKjB+gF51kqsip7yzcC5tlXnX+PWC8kF3vMhN1Xi2R+8Pn8YGz0Pr+cH7t0E
0qoozUFSQlkX2lcGkJZxuuQXZA6AVF5VVBaoV6AQtF94NqInXcSZ+YaaxH4Y0jilEF+ZgA435L96
E0J2RzQzNwM+6+HzrrdimkMR62wng0uUn34MUCtNKizFfjAL0V1LmJtP44XbNczoeY82KRcdeBmO
mh8sdDZiNxWnibLxs4dhtiAKzlB+V8P86ZTKpONeGAxZKJ2SMHd/LUz1Ieilqsf/B3hIlQaq0WNc
HYmM57Y9owZGE1sSA+i3Z5g6VzAEdG1VGij4Zu+psLnQJFSv98+jY7pgG6NoMd4ww30lP/Iwrywt
S/7+MdFoKDQAIU9RoDpaduNJowGNOWw6qn6CM+Hx1kVY2k7hYTLpCjIwJeyCKl+f057VyqeoqfGy
vdVfZ5RPFBWrpTpv3joos0KPTJA1/BVT/+MhKoXrJwNQGOmFQpSs3Q2zR07v3Cs2fyohKYogl57b
iCUw+g+OhSLT0zEhr8AqLW9Y1nGt0+HHR0yb9yQAEL5p+7XfLgYiE8q6wAJMzZcD4ISdQYBkGf5H
ClvkFS8soKdEivcUEfMsOY7LJuZZnkj5VEQY4+irltMa6rkImZNyF/x3Q3IvVFCRQEZFsOH/YlNo
wObGS0RGFKY/UDGyawX9dCAFx5Z6seAD5peGaqa7EZ1Jd9tmVkg1cNpRZor+B74tbSddcsrOsI0a
EZx2u7GY4ERDYMeqxllPXo9F6HDmjh9+fxy9LLXM4qx/CoW2wydIXrfWIeJUSe/n5g5Udv4tvlIn
Xi81I2eALj4dItVIJOwKA6tl4XYxOgbZpR+hXZ/II3xa36R+L7879QMTMNUCf/S0/cxd8OEpKR9j
tuaPRlX74vpF9vFJXKVKsbHag81rl9GbhuvhUM04b6sPLnI53S9WkdZ00yG5cHhFjrLXL+4NRSGL
1HWJhri3Q1qvSTFTQTMiLaW15OIrp/Rx1yvkvRIEkQN/cV1FoW7Y5ZTrn0nfBD3rNn2yjg5JXA5V
xKpCN4SnZ5OyQAB2j2bhjvMFyyRf0or0eLm8t0aDqo8TWpvT9iU+kkNhHbTYwC5aca9RoxvGPwIi
Gw6rzxWazkaTRANx88F1DY6tU0S3YpJZ866aU9dCnV0OnOvyJJIyVs3/kBzlT2xDL3iP8BqpF3G6
DsOCqaIZZ2PgER3gx1UPRJ0nqufvi5iPw48x4qKhROipclhnPE+jwP1P0XfgrEbLw4QSUwJU2X9W
H38bwFyoDElDYTJ8ETMjsDe03LngBYb7Rtj01umJbaybRY8A1VoBFXB6Inty/wlv772aHslwsZ3H
rk5xK4ySTOMwtARRGffKRPBz8L1HnwlAYyvOBwn72bTIHMtFhPNEiTT6B0knyunJ5SyWe2QKr7ds
9fqu+T5O8NC3ScSLXlDC4+wSYWiXCMAaYOhjKlrT25c2crb7h5xlaGDAs/uK/w+gXatU0sT7gFkr
BmmPyrOuBJFffjZGyR4r1akvuszwh5fgLKJ+iM1SYjujBMTjMxvaJ6K3uz8wwuRg+qhwHaop+jBd
Go/QYu5bbyzNqnNI8k/fJ+M5QKnJ6ls9qSZLyhFJcS2kvTxbXh1rb+yp5IbN/jQzfpPBosjtpSsg
+zQgyNrY+VUGGgY0HG1bpcPjKLqh5YVL5H8Nrsaqeit9oVroyJ692xDRELBniyFordxJRWjc6f4Y
3uxHb6kf5bgeAug7nF510uCZCxzuFDhB8vZ7f++jyg7lbxaNJignFzzrtM+bJYb53ouEUHZrqHMq
V8KxGxowAeXQ+Cwa52nzpSl8nPUrICke5y/QvLhLTFO7C867VW2KUTkC6PzqWBtF1GqWeG8xhLFb
ypAR+oIgvNSjvjBEO+OTI/RlT7s+ZknL19MSWGIjtT1HIi9SXxXsVMXr1tIaW8VomEaS7pdHJBZH
ABjCh4pMSf2Wo6aQT/4ZJSkEq3Y+PMvck7Wt26BzmxZJNr5OimosKqkdJacU4/A7bwT3w10AoWvS
7cjmgwXt3NG30/DNeTrR+3+MOfPuI6M4V2zl6m0dSmtgAsxITx8g5M8hapR64L9BxhknykmmLivy
Awa47JLu9qqpA8UIrtSLDJIl7EIKvPgfs7bHKCQwLEGO6yJooftC/pVAo+6zA72LZxqCZiyuEu4o
nopucbeLt/FFb4nrq7qVfck70m3ESJkxMC4CxFbr9/Um/ECCMcoVfgvB9kAdEvhEHAfUyTlVkclC
gEt5CWlzQL1FoycOEUXyeE7bSL77790pCo+Fjv8Iyf+sMfpozwZSyd4BV4zvenppXuknTK8hcyjC
VQVXhb72DsOGdSK1AfO8mnDSrwkafPEadpNQmn5a4e+D7see96ou6ux+zRzx9adTUGSTVJZgRJsV
89nIzTUleFG3uHGK7Lp0u1XdfofwlaG4Bi86cexgu5n5DPn9V5frckQ033ulbJGfUlpSaT3GrkhX
yTsHFqLa39n8CALfOgWdUirNDCHU9YBT27t0QqH9abUBRAiioH2jsQ2eWqSSrXeCw2m/6aUpHM3V
bRcaeP9Pb7KeaQSnOYygb8+dCJiOaU8MS6g1J8hm0E4+XQc/YG2eUrmbtSCQhvI0B0YhwHSuUZTo
9yCnEEF95waExCgmxyP3GZ5JlizVbMRmcMJOa/9qdW+Cn/NkSJwKAb3uRE2fteU5miEGtOl9AKE+
I621HO/Nw39X/v3i/MehNGwef/yzK5s8tHKshSxlBHl8156ohTVEQv+SBO+RZyTPckGfD6Ey8v89
B2cvwcyurfK/i9v5sy1xkbFKdN4HH7VRZsz7REwIX364WYDbUNrNwacIB/0V4gDufKJbUXjAV9W5
Il99mh22w391dLiZt7xtuKNrlGMhpA7KcXrYLgJQ9X101eEU3jWUfJMhCkI1nISAVcpBE4O3xSeV
v3foG+oixLegxi5H5Dp2yeD5BwBUb/+BqezYVydguhJ2ebS4F861cp4ifF2E3OoSgWkBqyEYC3aP
ZF1qbLMkzQ6rYiKxS/6HUy2IE7NzwtrbZnooa2ZC5khpg875t8562U9JLK60PnNvhZuLjHw9WJvi
F9R7QVTkS/jhDGXaAuwmruvc2kMvT7iVaO1xlIZy/cVcjHUi/guxFcEydx57AR4RtL6/xc4OVIH8
P+VxStTIoAXzQ7yfUaKp6EF9W9HyuUMtNO1WhYNuAz4ePwpnB+dPyjjk0tl7G/gVcLIzaBpcbD6S
MpziM02bY2jHyw7pADc91FW1ar/sFnhyhO83c+s/t8FCdoZpHD688JrOtVUiqP8tyLjER7BaHizF
pEBJ60PSkOfrmihuzPQepCROpo3O/ibAOWZ+m7STwvciCM98Bq0NagmVIdEkq+TJVh3NrjgR7ZKe
Wd8mkvv1h5pB6veQ4XMVhWXroddzNQYGxoqV3q/CYcnL3BjBORyAeXD4PTy1n/pMk00I6nIgT8LC
KqHI4xPOejA0QuST8wz1FQbGPnP+6+/x/Q0VD1ABT/OGnDgyYeCP/yOfnM1THkbv3JuvSvX6d4iK
TkEBsCp4YbCNTmTBEgpnqt3ZpM3aZ3qM3CMMpF/lQW2oKhsG+TxD8Qo28+08OmpZJYZ5FvGsDU7f
YimbXGV5UlOB4ViOMERM8+8Ik9bWEKU4OxCr3jEotuPZqgWpB3Atl4gJgG1+u5FnDxQeg/PnsIPX
aFvpFL0mN6OSDl/LxrOID1eRvcAIZlrQtk/T8zp1iGSGFS/p2TESXDuIsf7PfT4H4588Z4EFOE7P
/jHoIPLGPARX3LmQy1PvKlBlmkK9XqIyTDhnW8G8ol+wbAPCl/xDbIz9N+CbVQgbI9r4XYxwfMLX
YJrqrLyuKRZCDJvs25kapgnTluPHvFNZ6MmzAafCvp6lPOHVdkgpZJdcrdIMroi6ucW3HepjGqHa
colYu5FMae5NuSIBgvICJtC9jGwLAmedOCAOW/f2E6X2Z6mAzvsY34YEzKG+1puXeGkhL1uqa4tq
excUw0AGW//1Jg9rv6UtU35VCE/ZJu5A33P+NuaeNhc2ZNl7Zcp9SU3m78YiuS+7Zf4HF8jSrihU
jb/bhwnQ81jZvF8sIfevYbDRDIxj7BVV/vcfM4BG9fui4GD7+TFzguvZEhZpi2nduuS78SIjrhHI
sHYzg/mIMnoFkVE5atk1xvFdke/LAUfusDAqNwK3PKCV5PrR2G1LpP+NA1EXYEik9rLgGEJV4yS4
ndrw+aZlofL26A2g+WS716RvPjsK3ExBuzRFIpVNEkMLE0VKoEmK5amxz6V6k2JfUrkzxu9+69SI
9wau28vFmhM1tKV51EK7plEi08Yk8tMnXPfTaGojvnQ7+noBeugzziev6tjVaYqfgIENEed6Mmd/
lYxuzppjKGgrqsiGNDmEUI1/m1HFvE+DLNYeKVPNS9DLTzeQUw1ffYMPfSnxj2tItN5hoCclfT/r
TGXhnnUnghJnkiiRdoh4GKntMFJFetEsbKCuRuC4sniS52Y/5sT2DStsOpsxpVRT3syNAvLA9He4
GFDkxvklASPFWczelDlCoL39yJ5ejxgD8YpebzqxRiqpIcg+FQg1lerfPvO8A8TBDo0nn8FU6JHx
l+k+2fk8oJMExhYK7MBjv8u3PKJqSTRVvb0ZSN+fmS2qBYbh8npNhEVQJapfupr+UgMhshNhv8wh
8R2zZVhGFD+NoILD84pFNsv/g2OSCEbGq+I6TeHi/gWTD1Jw2WWz1c9FakwXftd5uBB1mljsCVIh
hQBhht1GyQ3BM1NkTE+bycI5gnbVyAn848diwyy1caXxy2rMuX7lLN7FHNqNto2KCWngv8IXCPUr
BEjcEEYFkSc2VXIKQUq2EMDlm0VTQE2OKJ2RwTHnX7romOsLUNnor9Gy8CBA2OtFKsbrTc4SuvDU
plNaPnSNHF74v0tx5K/olSaiSkpOQZAh4PY25txnJerbP+QePp1XhJh7sQ70ig2F7vA+D1Aw61Eo
fMuYNU5I3zjhgyDQvsCXiNzqVYm9Q1PK268qyurzri509gdO8L23TlVt9kM+WSqvf3KQ2RvpoohJ
I9g7BXb4bfoPSai/yC9zwAWug37bHNhDNjtgFkBAzp4MYUapo+P8e2w0ZaoR0avdcUhODpSUZrcj
0GlyrlqRPyDP1tDm9/FFnHqQ4vKmqUeDsRbyU95GK9gNu9ZmRdi9wB5VkheFo+p07zKCarF9Z8hH
/C3yZTlfG5/p/fgUnKRDejkp/Jx0LCpqUxftbQp8cmFl9yOQXB/ylJ5+rCwADc8rm84tNHVYoyS2
CvyN1THEHROyMsdQc6m9lvFW9ECIv9CWiNvSTK2oco82xWtHrvMLvOCI1oLwrI7z8BAYQeQ+xE3/
pBRpiMUpwuUBNkvgElxyKgzsGxYAln36vsR3IXTVHyNv6y/f+1RbfJ+rmvBxddczL2FHpprac/IT
QkN4cHXhY/mOPTvFCLYhTdB3RSnUkgsfWMyBJLe67VWAU7+zumjIBhlDhd46qBrWsf4u7Rv8++Fe
32eA7LqI5CvvXN0ODu8blzfZn5FFSXeEZmUyOQaPOXPza3iwD9KbAUjmuIy+U4FRbKFIoSuryhPo
MM2w8TuvPZ455Q0zbewpF6ldoS73B5pQfBCQJCoMGxLfOVj6OI94Xip9pMpWwGeTSZOwjqqzlprd
AkkGqxI6XH3wCcNLQ1Mo4C7iVQdWCb6HjTHRCrEeaCOa1aEziMPNSycxM0NoXjFE06grDcwkIryw
Cry9TgotmwVZShKSAlfeCaeeyRdBGlpF2hvLzwYWO3ATHRApSeXv8GoA6v99SaEHyJTjhYZDSygr
iipLx0lWAPZCp50D5+ABta3DnTXU4KlgDsy4vmIMSFA7fJx+v76l1RZ6HGwi0+M+hw10QI8yILzJ
Tvq/IM6LWg5iVqyc5p4WINTE5Ym+ua4gVm4HLNhBuBVqfNzs8cYyyKtyL3Ec6aGOPz5MpDbMv4h9
D6oRORLFR/pd4dQREoonJSxnI1BScI04nSrIlRznna+5gQ7s5jEz1RXMvl26m84DwmOcljfbi4mu
7RFQwxO4MIzr9r/2dZHv7GqFpF4YWLC4CF5ATXHIuMybYFIoPEyJFbikVCM/tQifkfgpciMn/xpp
pPlz4u6kjlzrDsiZbpFVEypecTSiKl9xgtHliqCwZB7rlLJuepYK+B9Fzww9gb7cs/AEbAnEQvNu
KWinvRuipZGHzq2R14xt0eup80mbRNVGmBkf/tAwoVp5jFfAtVOnFuRVngV0VBwjP9iYZLXqtJQn
v6GROBbmGZqVNmT3SfrZtt+9RldpXEmMve1+AFBtfLIfRXD5D4J7YySUgBRlto1lSi6zh54iIY4N
z7Szov0MHuKsG/2lpqpex0nsbPQBxkQtgbt+UcpgEeSVBZhOuM6NuFdiH0jBE/eHtrkdyDyfc0zC
e5Bw29ayA/HXllakeoZwwqIEdz+XcmXeJl6u7+05W9MxB5xJv7aT8n6BzfJXCR0a8IYI7kaV68qL
iYvAAnqtDNJdJognaNVQgI2pM9yesAJVEBpQRI58tAs5TSpKj148ZDmJpgzoaBIKX6oW7U9VqWiy
DLYIPYRfreva8YyvzVXBvQu366mYnw223hNbvr0PX+s1jR2MOFv585kR/XpDzCUJWKLnFmBnjTyy
zcvu0ivLi9cKdh7DNejceHhCja+KwXWijOPCrzMRlKa8UIrKw6N+R7Jw3kSvisgfGBH8OZy5/2f7
4BeNYKpqSJblc8cw/cGGQC10yw0xCgt2kyRGJzpGFas3KdBSHWbW8i5EqPE5FiGzRPNMPn7ETjmU
scZ5HVukwtxz1p8SMNVKqA7LGF1kV/mTsaGBY7x23KIbaDsX+QFTsekr2jklHSD795RmimcCl8Qh
WvUm//o3L+kMwA0WcsCiiQnll83+J5jkKaTEBDwzny0ZdjB+iZFNl8eCZ1un9vj+VplR8UImF2mv
QsFxkxGhDTgxQc4atdznWk3XgZ6/6ru6LLpZwY3AyUSkXZYSchXnLnS8ZlGP0LJG9a2iUw8ijO6t
lEfyk/zh2FaY2Og9vWfAD4D225SWkJVu5Cl+K97yAf7OZR2DKUZZG7E242rhoG+RMY6GabgGlhRi
o3pTn9tGZ8QbtEQnhOpk9awZ75xO0eR8gjOLovLc05VllD83r4aomPkzWvusV+blQo3xM5E06SsB
xOkqeyuysmVEXU+S5RGDB2FFHus4Yn+lMVFLpaojcWaGMg9qET3JPlOVkycNp0EsNgVPCv7QV5J/
5H/2ELo40YCOK2qwTyxYMxfEWDf3RHczZsHVrT39FMrotYqvbkcwfWFqQeAwY2jDFWgKM8sEgEFi
h0U1W4v1OzR4KJUxLFooD3bG1RxZEoHV+xyCcu75Zya/5gXj+2XT7/+jRrEGED5LtDZyWRI9bb4Q
Zb1pB8gmlYhMZIVLw3Mlydk0zMRfAawqiBn08RagFOC4pgLj4ilRF2NNrP1BKtX85FTDrVD2mngw
G4iKFwR/QJ/QBpTMlHNSrQoBI/UgLcncNC8d75BmOc0TgM9bDqRWpTqSIfeyr4SN215QMVsqskjf
TiOxvwMlCBLRxcRyM81myPRoZpN9k7jIaW7h1JIE1XhQgz7ZDB5vUKmnzKGeJwv56H5rxjQ6hfnc
oX4TMDLLQTVEKNf1+A2hzj+GMUlS2SWsAaznqMw/nLNc8lZMOWVEPjDGq4OlF0ZvrW8ojL8L6/OA
ogRAZRJ7db3q3WmrDjB6fXXqWbPnRfLfdmQxz8et9YL1bP/YOTg0QK9MLrirE3obuOdOrtPW1s1I
gs/HZ4s6mdUG2WpgZW6kjChL6+CNPwNATUaQG1ma123pxMnf36t3AyHm1jfh3CRYb+yzoPp3I6w6
cIj/Lg96TDjr/BImm3o1ZslloREAxcGaX/dMvmnnpwTCMFMfYFc9DVvykgK7BN3A4VBQd3vgwM7S
ywjL5+Hju8tkNw3RWft7oBXcnA5ygK4novvt20i+P1CxCWLEXAjJ7go/uezY746EBuG3WXBrB/EB
X+d6ToSmbJfPBzIo81GNxGR45jO1F/2FGfhmzNerSX2zyCzVzO5eobfk8YVBm3sBarvYiGDSRZJY
7rYgdPrGXZaxbECKg6fAfIlyZg72bFfim0tUpT2tNoOcainMSRlyMmGX5uIq/pZnVGMzZq3fkRG4
VHbnXbHXy2OYJH81TPtF8a3KUIe714tUD58SpJj5viNP+Kr0kSvbk4RhXDWrQDXXSWpefd5F1Pa5
6kjI4ZwgHBCv52daMplahonqhwtRq8sZ2ehF3fb2fqyfxdUfbHdHu+/HEitnRCnfTtaOee2tvw9O
PR1u3p3rmKkYWIj48m5XZUHw+VH3Rh2hNr67u4PeJDQyK4z+PYGZTKiCPfX2yxV2adVU8aoBcFXA
u80XZJZ+rMP+PiPGBhCwNgWja6LL+DxBSOywkmLEyNRBB7Ex21e5IcuICeX4jU45+CeZCL/As8+e
E6rN5Grpajfs3IvIvfT4fBc/nNwH5QHcdoj3WY2OLLHni2FGIL3DZ1K3DaZwZS6gmNy9ru+qZlwv
4ioLge7MePwp20dlN34R1AbWK+pTFhz+x5Tg2UXz5jCQCGpDZZZhZJJgazaK2wOPNVNR6zSqBg0R
P0/ldi3KW8sxuL/wu7ibB6UOOjarKlA/FaUvTvIx78oJtkfgr0C2tFxDDZBuG8i4s4ESrlruuDjP
Gh/ibK8W+wgrcgPa5+r1VU8ZK0tLLzbF8UACHRsoGk0ZHkzwGuQmT8ZwZzHrndxsFscimgV0gxnp
JWhX7OMyEtLMMImk4lcAC/13Cg0NFWgspXP8r8mVUbn67fbESFfkEuSHXQHbCn8jXkY3lf6qHjhq
+Gx/0DDd8HzGSGwIIRMHpQ/l64nF83r4/buphShJmuUQ9vcRuEiul++FaiZZFFJktcvEM+jRDmsC
vUcgPkva4a22N2woeESyuMtjj52N50EUArNG0hi73NUUH3V7xSOZzlbPB/M7rNwNp2Sg3pr+iafF
3vRCGWUbjLgLRh5ENP943OQKJdVYOtJiZvLeBEaD9qbiuOg6lADKi5IMs2CgUkXF6KSsSFgReKQB
SL13xplqd8LnbcvYmBFFvC0ee29nr7LeUS9XSQfLaLqq7Y5uCTsCKeH8OrZ2W1gb6JGrCINHHskO
Fc6WIvaL6EJMHyHbpxVx49HLmQg3s/vjbnqwIyp/gb++SizW5kYnmHOF3t7sLmJEwPqRtAn94NZV
MFJgFqnYrmZ8eepSS4T5HfLB6nYSMsGMDxPRlfClfqLvr4CgSqM+/x40u3nJXBUoVGFLgmswwvov
OGFTdV1GIy+O9i+wqwq8Eub/KzZJxrQ7UcUvCF4ASdAJaVlDxhepugX92O+pA0JJouITjwE9410h
COLBjQJ1UxwwOaC+iQdZHrRy20DgFLKdpYmE8wI1IX5UhXufANUVquC/ur48QtwGTKsO+ac05eul
03EREV9JlUytC4vBfpYUcYMhDn3lF6lnT9TydpvvhT0BnrCpyTxHMtZU4LgtGfSS+lvRChD/0o8k
238htFfuXjiNKl+ICTa7WucPdDZrmFsVUVZ3nxD4Zx4SU67PAFVfAKvBhIqL7lxNAZhmdsudv0Ys
KmECv1GpVG7J+zQwwd2GR22J210enltVJfaJO1Lv89FVZd2R7NTWrIhehQzO1ZeDIuKkmh4Wl4pN
etcku/TO9FkAT1KaVPsQAXs351cLVhcsBsICHcQdKEN9cW0ZouMpp4xXQoAv3wVnqc9+Lcgj2Odz
hBgOl6TnAkEXZ/mw1crtdVF4wREQb+oPgtnaxCqY8fY7Qst85zz11AZ+F4SvlskrE5QJlSH60kyD
AdtbgTL//DIi442X7pra0McnKeP+79z539Mry/DH2OHzUMo8PNe5LGarUmCKHPEQ0oMcpRlXGdh7
xn6fyWbHAzDgti0jW2NUltUEJHurKr1aZvPn67lcRhg3ZA1w+cDdKUWG+Y7lFCTBQChgoNzDQnKH
v9L3qNQL+D/piVwwEVoiGe+PZRkiFLUtZJyvbjOu3ueKTIMYrnFdixJfPR1eTc8j/A9BSeOu+7FK
+YS3H6K4f5D4Z/agbC3B83O8/6ROTGcg52KvxaaZXtz0b0FeiU3peRRiEAm9GqM8L25tYN3eXO6f
8D7W+lehE+pnSlexWsnSezZJgbUQz3zNNsh6w3IxKVDfgDSwNjXMMTzLZZlSiMVmJGBCbafNE/Y1
aRFWAk0G8YUqZiSSXz4pXxRmoMeZA3SHKT7cEEqO9XkCgFtQZHF97yIKYZNBt311einBNBwRPnmm
IuWBkzTpjDPJVi1Zzymvo9fH+wiUBMishAG58sevoyzFnNojYJmYiPJdYZuJNdsKb4nGtnkBptNK
/4NxiMe/XTAcxNEFRNy5lpC9f+2yF0vfD6XWgwO5VQzf/lQ2v0ekVFFycRXh9L+g1abrtyBnl/4G
yLjtIP+rsh9uk9E3M/Jl8RRmvOeghBld6wc529Fa+yYybL2Y5qYN3ZZ7zxNIA0PQ0ZOjKsBthR1C
nzT1Mjt2anRNvPJ6u+v45KSpfM1duf5D0YnMKQ1Sxm25U98JOhbMvXWnyBVM0RBBd0yhMaecJ70V
xf4ryaLLttY68jODbQaLSEodlVSEXtTnykSKhq8Ab2E0DUBgI3BntGXqg1+MrGXjC1Hr+G2KEP1r
AUn+QITSMNUvoYtlJPvQX6kWVu9a1mV57IMFCX2bsMdmcmfoZbx/WncGKlmij0Bi+f1TfX0xE1eG
YUdN0QZTvE5Dv4ECVNVKuQ19Eed6XtVsv0Bj/u3EpbiPlkvrKuHYkuCifrdrKqUAAXuyMZPOzw0H
8EhFXSDL8Hy+KiTX4XDLj8+0yCfTkI0PpBWhatzXByMbAiwCm6Fsbik+3KkrTH4frmmlvwKZ/+Wm
mLwI38NHIS0ECBwiASdFKE/ytpHvBWKHmr8IazPdQoA6b/a6vmqGJsWJkTC8DssFH58ArIjqmp5D
mfUsfrSni3527SVwqUJlC4vhK+//7iid0OU++NmnZ9Rg6zoRxdwyR5lnviWALIp3YJsUxPSmLfF7
bnN5S47O4VeKvcmIOx/RUKJ0JAsGmx54Ofg1jOxpvE3mNWniurL1P72R2RTW57y4lpsZX55bdaXi
fBfksJVG0RAyw+VAT+Y4TFo48Ms5qzlU3M1a4CNqAYEyjIGvLkkLha3FqTqFu+twUJYHUAWdVcd0
hu/beoitngWUJQ4ZQrcnX1XaYNfBkZjX2XvPTevsnlFHtxbgpRDB/A1EuG/DZuK8+ms4aceTSoLG
GIow+J76Dd5lsZR5TtiCpkcimkzFAc/PlLAwgEr2hXvbRjlfQ0k7jtsY47prszMbLnv1di8tNRlf
OTT03ueVm4fp+JleRBtCiX2DhEKejAdT6cF0OtGgFGzSzmyXQ+LmMyWFy7LrvHqjAjsmRn7QqDj/
iCiH7G/qtg/CxihNdaYjD4iMetqAz8guLVXjPqkXbyAVJqpFvRZAZ77m5o0SHhFLFxCy6rwKgZCg
TlV5s79ieDGwJy9b3uqSO3zhNnvPs4VOT1Bk1wsdoGfDp9F11Xq9WPYhNL3Sbhs1SlFdNG7M5o9Q
IGURJIXe8VAP9KnuVbp3SP0jvupH0F7fcS1U765VF3Vq/34IfWxPAyeA0mzgwAvpFydd781UD6Sn
5gp6YOI4dJWzNAEKkWry263L6H1+xoOY73+JBSaP5epQniBX5qcrviRRvfZg8gKuaj9YWEhy9dZ0
qG4myiobKYLicxzy49HO5ioJn59qf+enVTtVjT/S9ER1DRLJOfZAoQ9QgFiU5DD1e5CLFcHH01k4
hTYubhGDSn2fwpL5EJJptNqaYjK0aOGSru7K3fMvTpgJDP0CBAC/A9QqOzLL/fBGMZxqw6MM7BCT
bR601HTM0AbEpa+ic7MPdomm8xWZgxpxXA60H4paXD0jNDIaZ+xmxhA8C0leeDeZgtXVtUZ0IbSL
yZBYrTQRnacD+QrFJfPb6YGTZvsCjRW05n8RSssAOK4n0BVY/pThdLFRtF26633KKw3KpLc9Vlga
1vReTbFW9npV6ASdRTzgYv/GK4HOuJvKJc5n4RNUVoqWBvA5IsmqkbS4locXlEiakRtyAjGk2hhg
hrbXT3NFWMSSUVcKFuYX09e32NaXNxoIhqKaRBO3tVEfOolLirPbVWFFzkyFLaLE2GwOaoHGj8Tz
8Bo0v3QuezQEMBrK4sxlAKdAZyE4+PBUXhTcSChyujCbUIAvcagHDJYpmITEFLPO4kJ6es1XHFqC
bBCALKxoUcHyEZjuXBwwYGlBQ32KWeYzZRjO3BlNzZIc+z41lNjCvW4zGWgDHdLovvjsnwGflgX8
gaKo4UX9cxtUPbavDR+J9kxWFG7S6iPKL6g127wRL0C+ZLmYPpYSF2vY5kz74SVsrS8Qy4pMy1qg
aXrIQip8pS63FyHKhYtHWqwMhaT2bz2nYUg8+ATmpZ4V7l878HcUalt1p2HDeNTb+ieT6YXG0AIu
aT6XO7ifQX1DbMog9F/Ca4QJJb+FLfjQMWT+MsvPrt+vdQehqeKDuJabFkvegxjh5Oe+i5J47u6D
iUE9jy0UelP90ZlUbSgvSc+0/tD5S2NEWNV/Pgj7QypvrMhxbbUxhOz1p1wKGqBnN5FXqddyLi7+
23mCjx/nli1yeQYuBQWyDRTzZpTX4+tXfhEwPE0FUxHJFXPTQd9w2QPs42xttqepjjqvNOYTLmDV
tToBCUJHX9NzrDYpjEMPUvs3tCjwNU8M8ptcko3qWtRi3hYpb4no5qEg9WZ5xkZT8RtN0HjLLxGX
uXguiOifVS2PN9ty8GB+adZiSdC4qQ0c4ZE9Y/ZagPPj4tb8ymuMXO0yKOZTnUK/kDiI/NcfRaYI
BGxN4jWUqNS6GfzxKmormGjhp8ldhQFtUn9v7ZLngFz1zpYbjCzIDXyTopwIRZvaYkESYWGc3Vx/
OAfycMSv05pnKsdSya0ivyNBTyqdmQQ+hUKOOx2V+rwbTFzzUfZ/B/psZLWPJioinc3NKHXUVWcy
+v6EFaF2ZaPVbnycK2jhaxMb9mlqXPqgdBUurgNCzFwX9WH+tphqZ/N2qiUn8+ft7+KTeym9rduu
eCbDlmD0RR41Z10g0bM5HaTXnfSKTcM3EkcBG4VBzRDkHSUVUw+9zSztZ+/e8nFl9FcRfcXm5I4A
a2sT/f+eyhu6ddkk/4Spu98tkIi294c1hX6JyKgeQVqJlMMFFY1Be+bL4KfMVyeVb88/L4DLUAqV
CeWMhcQ/T2BVFAl/XI0hGT5l/YV9WwGKJhWc03yA203Rjqh2MRJdboCfpfIs+XUfa5QkOmHF5h9V
JdBdDPzK605aza5mi/q1AioPugs72aYQgpaIWIUd47ETAKHE+cUCMgXULGbN9jNewOKe2KHM3l0V
/wwQIejQTzS0tesIGJvBu/uu7zZpESWqZ8Mc7J0xz1EUvbyvzuWoy+QFor+KBuFAnYKgZkNZrA5v
lXnnu27Nafb4yjDsh+bFosgOQSqp+24AnYM25HSvyguZYsOc8o1AjJxmfroTipbU4SWv6ibxlvrE
9hjLdSNsQ5fJuJRhvNYEvLOnxnj7lan+00lMHjXIbA0vW12YZYNZrm+5mj/Lv7E95KBQVXAFGKGs
ZcECivKtOoYB7Rep8ffKnOFQEcLi4ZA+43S0yAN7fXzi/35ZlTNWwgrWXM9PqQzI/lzZx+rKdHhf
ED+wekTbWy0eSzd6wjFnnRjcDmmh5rVx2Aw+JtVgZR4ka/mmKC8O4hQbSeoUP9MI+5xos/0wsDXt
DG+qLHyg1+ZteCz8ZTetY37b28hS+USrzb6ZE/qiytNKh3l3wbuJbwdMgI1gZd9fK9yJag+Oflr/
HIfUsOX+oiWLgiIxx7ImnWYyPc/IgyyNb+cRTa+JjPtnaIrGsFP1l4y/JO/m+lHU7SyOsG4KTCVE
rXJhqKFevZDaLwJYK58v9et4Oo0CDTcS8Y2SDwzt+Qht6MKvG999zB5ot9ckbhmc5mbDmlzPgPbk
0iHDqITsJ75EBjJZ+JGxYm0FNT4F9kR1aKcZQLfzGIDVDaxyygPolktxdx6FZ2pEAAz892vV4287
epI1qQvXUyqgneAA27yvkJk6yZDURgDDB9/Bm3BX/in+dCNebbDb44RzTejIYJA4gsncuoOqASgr
vkBkUPaO3y705sNIFHWjWa5XA+qGifu2GHRQex3Q3powcCziDbI0Nh8+3NEvwqaG59gsW8LjVOS7
4fzVFlgClKNBfmp3cep7uq3VmcXcLNvtWCzAEmUt5MfI8jdR5jkdxnDzAjz9D43nTcd5dn6A3oy9
ldvNxPUXC0zSAjMnYzodEpRPurGWaCX24pYsezo5VAkvM1QBZpiKwkRpPzBdKrnRf5dZ79RBBXee
kH73XdARtI4fqIGxK7gJjhLsCmXyRskjd3ObkLgSqowhg4enP7oePYyob+pcFtYFog0JmEz6qZ0j
6c4anDI0zJpTApSWPFcoeQMT/LCm/jfW9MZoPwB2l86xwyE8lBQe77MqlMVBa0OwmfYR+oonEj8b
AOkTduGdjIRsy5bwrteBxpcNDe31g8jTeaB858eupyKeOVFlBHK5iLsRtnjRfF7iaCPSjSxVve8F
xYSRvt/zsRWcYoyauz4W+w8ETBLnzwVtFGsZeCvpk2FjJWCuaWPPrYYG9n6bJmLjb/UAxyO/lK1u
J5nVpy0UCYZHNTvVNisvPCqlJgRMuRbQFVr6FXTX5uiyGRsYSw82BFvnvU1a7/r96tpJrApviVqZ
8c9z3nZLxjJonX+YcXleJVjRyZBRupqILlM3LGNGQppcIkrSFCPM7/aregh8nVp27ZQ26lzaIPEg
d5PwGUdBakalvgM9++QUQulM3vBTmRVyiIOAFPQrZEVJD1V1qimJtTSuEMeHZFpxxhF2HldDCN8P
8Ag/Mw6n0Qq609LiplSA42xVNI4QR+dl9mcSd3bzkJJKyZSKZJHAPAyd17r4fBkAbUt7Uqmkka/S
MpXcdfpIp4IHzDBiYHyK61VbbRPq0CZSJGQDj7vLCJUa2sr5ZLG6EhgxPl4GXZxxP1nRwJta5vBR
N8wjNL+diRnw+8CWdCirewf4CxdkC02Js+XXTxZpLWVXk7OlIDDdkYQ0IKPUqZIW8hx4d4+EhpsS
Pz1GtHqUU6DF8qdjCD/XT5HPV7ts7lZ9ltnEpBmN1ivJiD+hxmri8NxRaC5LgGIimMwXPqTTOANP
XWl+QnblSUvgBzci0o+aeabxFrz5Da55WX3bo6cxf9Ku+HmXuAmUiLf2NvV9z+HlnoLm8eeVdnN0
wZUdpzlcfwW9cAof+tC/fQdqpDJC/IqyU+WWacBcR9addDOKuI81pZZUIeTSk/PkDedb4gAWrbTb
28RDq3nO5m0UPmxZCK52HSwHJWOCnrjbVFzeNw6dqKzeomx8U6+Gt2pZsCFiJjuvjCRvXYgEY7oZ
DYTKG4ah3fY+dSllatCa6b77bubjCqisoOpyuAacparcW9jgI/Q3zHHrH30TMD3M0XvaAy25G1W9
WfjF+MMYMkcp14QqCFv0w3ASIimy9PwSft9E0JEw79TlP9j5sevzTyebenzIKS6LhfpceCqgoxGT
o41w+m4DspVY8ZwboqoQ766GncZ+B7MrKjRQfRW9tmah2xAYrQ1A9AmcP7SNY1wh8q3b20wUWQwU
8mPeQ2BzN+ftsX+hPIOA9Byva4kpZ8Tl0OWO+kGTLC4PcFocVlIh83gR1cTf5IBQD6sWT1OIUEOy
yVBBayms/3OYgPpU3hYXxZw+nJ2NidVvpz8zJkgpNIMK1/5gHhhnXX2XvcJIF7wXcR68T9ThxBNa
jeIWeHB3ntfrrq5IW4TW0j393srGMxwHtlCdxLRNGVkFRfMROUA2Uee2Rwm+lI5WOWA+NAZ3oR7/
vvPd45ktlOUKTsK0P8W4lRx3o4UKWkiYlXD1f1Xe1r26EnoezlXLiZTvVMIlU6bgktvI403HIZwi
nldZYKJJmRUAmsXoEbMxW7wUENbTbZ7rA3RbuOeN7x4mVHCiJvaVyiXjzh7xSkr+ijTs6+/cgPgq
EIb0N80c82ZPXX/xtS3d0QzuARIg3X1WN2s0pmefwE7JuYDvkYb1ljRK9iAcykxdcPyVBIYN+fbi
iQL6ioeytzVd9auKDprSDhw6JnCkzWKqTwaoJoEgCURrvWD4sRB3bjitV3zcsqI6WvtG33eHP1kN
Aziaho9TaTctfBKKYeim+4oPDO84o1qvZPrZgfAwwFpojAAY95qZWiJvTduaFplylHyCEoQRZNIf
BSClYketQViMPbJBLzNN15zj1OGqBD/P71YXJ9MsWIY+I8h1cD0MDjY1AC5K/stV5bLitcrovY5q
7anJTFWdg4xMBZoiFmtOKYZVQqkDmqQylyFJd7J7GALZnhbq2j2g+HyzJmXbYvGapCXJ7m43RlTX
QCw3VjiSqoyg5zWJEszyB4qygtUHRnP2lf5zpbNpOFwQSJlGvlSEKOagY55RhWdEqcexW/bQia/+
rzq3sii8UYtI7TmWj/nvTwOD1rJzVYHs1uMeGrlXEW6OgQ1Oxc7qKDn9ipM+amJMgzMYUZVmAcpA
ptnAOnFxgtL5F04mZ+auQklU9r7wLv0DWwcyiVjXC+Swlr6TJrWvHeasu/d6P+Zw9MMUIjIvIGge
zZRO9V7Fj0mwe9nw0nn6pG+r6v2UXVgpzHTn8RH67pKNh0RhyAjtAGQffl/Zc5sxl4ygqJMTN8qR
zKA4e1ZV4KzM/Jbue3qvvRtQ0prr7hnPyrmityNHz1by/kB+gdZ8YQ+c2JdOjuEZOgrNO40ycT3h
1Q3GtAseTXhrKOmUZFsEbK/F42bHP4PGgIChQQ+RcP6jFXnZ8FNStXCgW6aFhYwoxCY45LXOasCo
D1XZVb2zHejSGaTRKQqSfG584TS1c8vrZ/wUlsIM7nU14Z1DYMx/kq1v0n9UeBwj+BEbN3aceafe
0HEUXeyPNaYL13vjxZcwT6ITgs+bBScOY/IaDWrccQrB8EuQ1bUpo60uK0NZ6mz6PYtqHgo2Lnjd
1eEsX4rP3NWOoMozfXTmyljwkU7Ie94G6oj+uKnQOBEnf8A4GOCL/QSCPCxSyIbtEs4AhqUhiKtx
INcSlVkr/Av4bquSsXqzR5Qqo8u9gY6u5P9it1E8p9SaW107jtv5nrNAE+q+IORKUYMRvRWbniRm
6GbjmCiWIwZjux+lvov1nmQ9EnT+y5Q2SvB3bzZBJ1TdIhJTr1R/6CLcZ7Uane8/VsaWDPxd6k1O
4PJHK6s2sNCXjCOMq8cIO854K0eMILLljCIRW2fQ/CqxiQ0OUxgIXH1w6wM6W4tTw1gLsiUvg0wZ
ks4rsydoWIityy/E6QHjmkD3AOnmlkdJXo/xZXwCO714IQ4Gb7R1W4jS45h1ygbu9fY7t5lQ/OHt
Ig6YDj36Kw+/Udqwp+CzdmzaSDHcSygosXrtKmYGQ9obxn7vpTkvJG7ISFUi0SnEDxzCGofEQOFH
2n49APAkkV8tmURRCW4kfeb6RJ5KdeUpa7oLZRxEZgCHDt2LTqOm7hkunaOgeCTOc7dSiHmEUXiA
t7bGk9nlRJEOvR8amycnp/TnhAlFTzxH1pgESstC2p7cjqE8fbaO7iryqM6sFSSEzDltlx5UU1r0
fe8tVddEW3mLY44vXrQFsnT3/fbUjVC07ud47IbY+3fZi67PXiaT4ZXXqV/zKTsdE2siUzF3gJvo
nDOM8kbE7s6olsFXBqZoBQZa/4uJI3Dl2CMGvx2mJFHZmMqLhquasgKtupfDRsGmpvlhcRA/DcZN
4aJ9PGzAeMNBwOrtmg/E0bGDbMs/lmgG5y039MrMN0A0KjRmDXVK5AaBIJYOioTTxXL9ztjL/5JA
+r1743Y63VY5SKjgldKZ2QPgox7aJ67RSLwMYlYmohODCafF8SYXNc7Z4l/V5izsuVj9fw7cjvWD
3aWs6vMxyV6EveaW9vdg+jQyoY502GmDA+j6s6FIuMyJuj66rZSYQTjzu0FXMR9mSuMITiwRpXwj
kR+q6XZLMNPMFESgyCe4eEd0S48ygt6ns2krQ1qF0Zg8edW/OqL76D9R3dCRKX5Ic6uNdexQLjpL
eBvZX8FrAC3KLkSzcidLhFb9dci8VwWhhUsM6Z/qBaGVxPqILsTXXFWqRR/Gjl9VAl+2+MA8kQj5
F5iYpLh/ljulNC6YLzklixLO3UASDDvmh4A1L5F93vCkI6q2G2+K21mB8UJx1Mt0ellirIONNyM/
siTlVaWp+noVbfQjSXSkWnjZ+hbzrnjYO7xG7t2CIQjZG9kqw45u3TcRKHvDJjCbl5MU2Um4zjwo
SYcJAKSeU9ULFa4rGOjE5+QXZfV2BiGOCdd0Vm6PY7y9r4lZW/kACU/vK33gqX+oWb8DMWnwksjj
PF89Bwy4MqtVglReHLORk0QkXZOpRpDrrdhkcPHeQyx2dpjQD7XXBYn6SfK1t+Qh8jpPf0gT9LTf
ONpQYPiPudisEUlcjOeS8VA4k3COb2i7himYMqAmKTyonHWYhC6Pl98/Ix5YJ8M4u/8R4BOJCx61
jmhZUBFT/pOR3c6CayF3C5NNq85O5iggwb8BuFecQQSzHFaYujDO7TxLLSvzvaDf23cQACu1pq3i
QAzRMB7pOLyNf6DA96w9agg9OXyLP5QDn39psY00SGkh3110SXjbC3Qru4zZFEA5STsb5reK26O/
t6SY5tQhJiPL80A4ly3L9KU1BUYmqjnavSj60V3THHI6vVGOH7aSi3R0kIlqRVqz5VHEjuxTAQmQ
/yK2WvAr4wYZxFr8O1rsMeds5n6UHRaOBcw6/mJJ/eBZjCFQ0OnL6LZD8rkwBYKHe0wBlYR4Y8ua
blHyI1Py/ir+hZDjG7PjNsQgChrQ41MNoycMOh17fx4VGezWZYSHVYBCuQDSkIidlW/m6s0OMgsq
You3c7BV6ZLGXINAP+mZfWn7+2ciM4Dcg4naobii8xAihjmHVRcnRTM7zRvNefLmIvxrohE8dKME
S0rT/5qCEZY62QCO8aWn/RZup9BgxYaL7dpjlPPyax25HNZjz0ElWJCI2F3sLYqR/RVTjMx5TJjj
OT8P5PGcjVE66QkDVEDPTP61QFy4b67nWQq0bTwXD+mAmliOHJJmP7ZWwDbsR4ZkEfvvf0DTYGzU
nEzqfuXSZ7zRhEEf4OdYzLq01qowNK1TEKndb6E+Sl3GaPAdba7lF/V6LitqqYbsWujNp0Rj2odl
eJjVqx4fALyd3XyAOiU0FILsZ7lCIjQAIHO5iWSjtxXe4K4qfg5Q2sdmdVq3kcyXFoK2XlmcWsx9
gqS+QcFIaDQ2MDtOdsM3PrIRYRVz4P1NCUk5uxIv1FcMBZdsDTYpciG35IrP1loFYNU6aIRefla5
qiITGXEZNre50eOdfvqpw2S3GAzLhltYWGASufEaQLBGtAFDQW7yJ0FgcYS6c9h7MuezCCE+BH4Q
K4o2BkvmSdFA/FEjMIyUcM2fK1TRoW9NXpXaWUeyDoTdj3GDo3edkBrdtOdhCI3fEOfB/1SMKRsM
m5AAdweV8InLuXheCDSpa2s/E+mIh3qftUwpiwaTphNpkLa8yPyfaYSXah8bWzTr+wN0UZozbZPO
gSXI0FFigDehSgRFPlPZMuwVD/Vjy20JL62wUc/++ds8obUk9mYulrli/aHdCf48LdtFaEARUVU2
/pVMV9YjVCJqreZPnQxRdi2x9aCHMjVLIIJSwwuw50mIk0nF9CgbW+A6I2NSbQOevrj04dyrfzpK
02S5H70/aWK3ykpSNHc2mQYReheaFnyhpv5TExAuCQNLFg/APvR+xAUv9J/8Kz5WPPq03MuwZAGy
dxo6Oc7yiM31YZ0BeWBY3umPRkN2iXt9kAN6CnkBiDa8+N9GYRJZirxeBbWE60fz0uRU9TPjiL1k
B0IJr8A8AKaduQ0JzDzl+v97sk0AolOWDaU3hw4wte/a77Xwe+iMUf1bPWMxdGZ0Bk3t+bgMMH7P
PNRikKEv+AaPMLBCvtHdEJWw78UQ0AKuD58Un8F9TTBMlNPMFk6v5VjdC+TuQ9QNVCjJ7co25BnI
NtW02Mr23lYrf209w4aLIz70lw4RtK1rGM/D1WbnuM6nNwkEHJJT0x39B4l2TY2WjvR1CN1TA2a4
KksD6K+V9flvCH2nXHSRJlA9aCDVTkjrKBOp+rezLHIMMT94nyeMCcVnswTjGPRt3zmEwNaAjXzb
1IpoPcpVHIgf38C8ruMOcLJqJdsxR4PZTXYw+fSHKB5gDmZ0ugwhkOzkCkfBdLYFVJ7zCnHW1iWQ
VExgdeKTAxLY6NNzvu/oTpb5WK96vykFDdhpDSSDc/a3BuIl+67U4LWyxafXChJPSgfKbXy6xIB/
NAs5qkLuXJgO29iP7Du5vdncEf/7KWXY9TsSnRHQmbjgn/SYT7ocoNv2Xb0+NDeeWCb8v5yqd88S
KjTGth/xnFe8pQY5YzND0i4zeO4WtIUiqJGAmpo3M2bItbtkuSaSLfa47zF3T90kBugGuElRFxt5
04kDa8LyAOPY5hV4wncMA7H2DGlB3fLLzd0xGL0SfXT9rQaKPaorP2Z6SqOXYTdpbniURhDXwnW0
lmNM8V1gHT3G0ltkC4U3t01H0TxYtqSzd2HKFmohGiqMnLK9qII/R+wyYtaHQcS9vTuB9r+Wk6Dn
IbUpTrSz7YDXEW13UFQN8JiMGxBH9CJBUiRdud5PodL4E3uOO/AaooxFz+GancqYJ/kVolgXfqUC
Aj75keJe9N4p8QJfwyT1nJR6Yf1FKvH/6tvC7SnFDY2nFnH+48N24hZPSZhyQb4RslRY9LEFcJC6
CeRn6IR9IVGh8rBlaRR938AFrhe0p8bRH5BB6/yZa3OMnek+QRPRm4+1ao7CJjy5+1ugQlTBWwVh
TFKNhgUnVBtZjbqcreLaWfiy2Luo+7BypGMwpP5M62/KbsymLlUcpCZkygS0UeYHbiDYF/zdPQKG
cqPbuQ7Et1clP9hB1ab81VG6OA0YXWsUV/mq78puGktMjr6hGduCTsMPHtLOrVhj4Q1BTRDoXlZl
muo1OUQ8TeaHqux5K9An0g/p1UmO4DbTX/V5GjtuHtDj4xRcEdoSGjaH2mhWvRdN7uqpdFFKiMx7
4wDNB5lMMx18NzzE/i9YdYel6uQBt+WHiNpAk42iduer3UWtUjxAlq94BqDOKWGTiaZd/tN5K9IN
5QR7dTa2JrjvBRMV5BBy/UlavF100s8ndv09ZD/rCj/oApxrUZLvHTcyNhKW78PdGb+AXngPsccr
9klhcM59ZLjdJnvhB+DeWz1DUnoCo40rm36YSVeItJqEMVJzaGMRNt6qOCVI10xILQhA2p5RYZ6w
lfN24BA3Cqizy3aUNnQaatGH3LXndDnTRKqzIELnj1FiIg1ogZCKFSdIKd2MCd2E7YF13CbiUz39
76sMR3NKmu8LBkhxo2aHFnzAqlduNGQQKfz6A6Zx/iy//CX7xDqwFrAO9FW7RDJZ6TZYphCkLq/F
cDgYoVX7RlirAFmMmjD9w2yc+5juTrWAi+tgzWUqhYixy30uY6zOqzsbASnUjpauZz1ZI3QIHIQk
LHpEGQ+L5nRU2hM1Re9fxZch6ASAJHiuf/mbW9YXterR5fPAhtmhECrpMjaraSooAVvmQgn+aFLo
EsdzKIhHF4bbC//G3AmQXJEVKN5nLwkUFcxxim/kMopsqwjc7jrLb9lEZryTN+9XeEBndGCa7M90
u4dQlmsfyMzJ2WxBFnwob84cjjts/NGD3266wky/fLabgnJLI5Up+MYDXW5vvVZT3Uo8ZHOSwbcZ
p1omxfdi0q6kcFhAONdQ0qXB6zwPEMEqEEuHJZe2auTOU7x8nE/YtaR3Fh+ntJEoxvN2JBWkfkKm
bbJ6TucRQulE2Eetp6cTsqJo94O9GWyIqARaI0cK+WJjGZoyqNcZWtKThUH+Sj1ei641FtWwrCBK
C4NXR3XO1/MBaBitvrgQjmi18ZQYWZiZ5/C6Dm5s6Zex4y/QUcfEUeKAc9H404on21fRjUB31f24
QrYxe8tXNirs72tjFYA0NX5sVOs/zkAc6DKt0DA5E7wFh0OcPWQ24yBOmNTzswfjCcKrVPr0QbvI
eh+G5Z+syc28/GmdvQXGAXCxvWPcsCEk8D4VmG2U7CCGBLn+eAdX21+mlpWqOB8cEzBeIl3DsWc2
dd9j0fOQ7rFiuD8nsCfVhwP7rx45TdfEEgi2HZ4BPYVw2wZVcNB1lW9lRMIiuj/XJ9KsKDNokBbu
3MRxCnR10x4sJFWYWVgqr0Fp1wNoI9Sll2Emek6UmRk+yZQ25UoCteE3RGWgkPphWuxr+aA0eZKl
ZviFcxTYD9IXBmpjYqR5Max7cn0k3tiaQOx8O3jKRRjac6bDIpcfyACq9jgpl9EOYayBLsFBF0Ki
cW26oh6uwTFZrswfHPHDPyM/Hza/OWG8SOuMfP8csZVuohWn4HrATOUbJG6N+xwbpWKUocHwk4gj
DuCKb7A8rPu8rHYGq6iBIOH4Kb9TlC6Oc3nic3FZjopYL8ZVzINl+WUjyXjm2UjsKe40gZcWvLX2
cZyScEyvOw/I6CS3z/oCkuTBLkR3tV0cTWpiHKKl11WnFmndP2Fry3cWmm/byVLY6i82152BU/Yj
S+xoyuuyTeiZ1ZF2u14dDsbxCWLUPBGdvIjD3Eagp8Jxtfh+4CXZSr/5dJoT/ZY2wyP2sdBjsRck
GXn9rBYZN16KslFRnJIJ1A0TwQTjWjU57yOemnH0OBuV/JzUyjHcaUIEzt1SZcb1jqYofhsYENat
yfTF03EBK9gcbk3C6h64sGLTxI/KLt8FywQbI6Se05yqeFCwRIUnBy2F2OgOHh1ZbcRNTHZ3dlTM
TOcBL9307MGR1VD+2YMnxjCQowFGwy2X6ssGqL1VWUguFLi0fb87nDKHbv1ybTAH2jUsYps/V4pc
LbyeObewWZ1huCHDICXPFYv7EHkLOOGea5YgI2OEh6F7lV5MGyB0FdjQwskjx+bE/FhG9QnYxeq2
iEnXRmGp3Slnso721WIsyXjRoeCykQZ0vvg6PPKi0QiatwPcLNGvyOd/ZajizzflvKg+eFtcQOr4
cxybMiePdCz/jjMBSEvSP6foupNvJh0tMjCjad2icG1DXQnyzTZMLl9A90SmcaxR0b053EpjdgpJ
j4onVZrxEHx4OZZER1J/tUMab5FSym+5etUVho0V4LNu3NVIOnBM4pFJLP2gcfVH3QdNeteob++C
grXKGnec1NkT8YhRU1F+oXBNrlm+SwyZXIyp6txTsshj2z9S5h6mNowisqkAkH0HoXMBYoMli8eo
T8KiZ0Vn29U7vmHURTmM/v9F+3wTaQ5DbXug31jmkoz/N/6fq1bsfQt+Jk3Ka3KmEtVpkeeuAI68
lZapvsypID2eavVbMVG+0rK80VLP4aL5x8eUSZoW7hV8mXEu36JwT3oSDozcDAk3RVXD2GnjSySN
rLhqe3Da3pv5jliiKTRGGIIBKrqIQjyTKpavtVIbEqioUdDb490lHjS5xY5mZNr8A1yA9IKNlQz4
QrHZjGeILFw6orEkmutVakphQRGD339wY4f3xqAj7YLaVl8KwOOti0l1/an07k1IWSSRsoKTbXWG
w6eripOTfkMym2LJEMVBC7bLbbcO2ouRxD0WD3V12wiwKguSzXbs9huTOt0bxgOs/h3OXYfBGZYa
0+xuoTUd4tfq/xcaskgoWH0nAYMDRSqxxZ2pV/76I97bw4cUc83OsyKEAvF4FinExIvdhgKODzeY
cPWHvqY6tbhP6ht6S+dJfd3ES9LVGEw+VY+mGOr+AYCCVxEm5SboIqKmjNa38pVtAQJsc4rf5PIi
IBbn6ESjzvIxqxNAlXbwnmn7zm4iZSNdqMTRxTPawmtA3ofHyOG2KGy/HkeQ88AL0AyD3ocBf6wq
zHVHYTn3l4v+yVaE1AxaX/chWicexqH77uzTMyfdOEWz/NIrS4sDasJ1zIm0Rnma03L+17fMwj0R
FKZjkCGUjbqA7XjEEcUHspshMyL7U12duCwobIMrxySvQpLp6dq785PMRPEammNodYhyyJPtgi1d
ZwrHAMfNK0sXROnOLFoSCXYByGm5thC8ANw66vbammOkHx+5H9jG8xXCG+FL0vAMxfhbgMpNs/ho
ZVkD73QwL9kRsRWhuYTcos8npFCUUAVCA07CiH+fhhN8517W/WopD7qj4Pt8zlIUmX0JQHmHZOll
EZV/wGZOuoQOetyhywKYh9RUcUL0BI/o62OK3tkqNUzDuyJ0J4fKQLxXIeeNAV8T3lpauxoQQT6z
YFKZFhjf+uHWOIO5/rQq1xW50rk/Erm/JYgSGcecqVse40zAV52t4Aun1D9sUWHdT8uT5hck64Dq
WuNXl7NBdnlKHIjz+OZJ+LpRe1QluV+6yUqiUxGnNgZmNc7KLcxEW2IZhh7fAnk8pylCeHlB1moC
c2qAuHqpI17tk5tPFr51JCeBaayVokZlXh/cZoec0l0Ho1NxcsXH/IgRWbZ4A7LNI58573OopKWw
kLnpBMuU/oPBseGoSgXKspkoAmq2E6efjdZCA8lK0aEiOv6Ufm5J7XxzHAd4dEYb9hVsZ2o7wAWk
0dA7OmGwVhO2/VfL5igudoLY7TGWDprWS6GiIK8LwXG5TOMY/frVw+HawcsvEfp8g0XazZnOKg1E
t28olwtwD3xVecCB0c2xc1H8k/Pbai9CkXfrqW+ZCpj1IRvQausTSSlnLm7vFEoEKdy1Lx9vrP+p
1ZWzkqCdwauJE+7YKr3MkutEgHxB5FU6OzMazqTOtmEtPoqAXHMoBFNjavhxIFVgojsxhWHsGkFY
5DFdSLDqXFvvB3fmee2oSsveJlL+IqufrRNt6xTJJ69DH0c8+qX5rPVfBttI8ZFiLhPWihO8PbP0
f3ZkV208JES68v7YQs7FDGSMnuMGU1tFgtlSPOTBYUPV/LyM/dGqMWi9vHNVNyuRQiPEW64I3H/k
UHzSAWxhEQxKkCcPKxk+r6KTUGE0yyobUWKShJhXCPtmUUJEq7gZRNsF5+uc8px66YeMIMVzuUub
PZUeO2zEPAvTq5+TES1DpCm/+RqyYtUpOZlqjfJU0blCdau/YNYf9DplXxwSo+Sp8Qc8SNfwthDt
F6k4ghVTFuuwIqIDatYjnl6SUy2ME+uJqtDLM88OfI6/MlLRjap427okJeBEw9BfUSMH1emjhYxg
0up829LH/yGhXbxW1lz/f9T4v8IQO242jRguieRvBeUIYVdF4z7o3y3fnDyvfGzuzkALMsbPpvMx
7QgWrucAiLr0GAuPXOihBYEAGkiQTlcnV6RAMUWFxyO0T1k1sktNy5JC9Mnc8V1/ztBYewyjQaKo
JWv3rZnPwbTBiJ0wgZuCjZteR3rAQ7QVsG+J9qMRNgyew+lFU9VGBnd3qhCDhWE8Rb3EbC86cLMj
W/brCYN9LioMD2R+Nw6DIeDeJU/dpqsrriamg2voRB3djeVOora7OkMjUk25fNNbY8hoh0isuYjP
3PN8hJC+MDjkRtCQ8upQGrJQbk7oArcF+6ih+eM10S7NqUCspfnr0pasSJYezd5xw5i+qr3CoD1V
dcPcj1PHzEa6sSoyqQuvgnssG2G2Ozk5UgurQys0qBmE55OhrT/kqLGujQD6AwlmdUIUfSyYlN19
JpggJxN4LJuvEcIu3+wh/Vu1sFGOPP5W+CX4D7iCVieKpU+eYI9yw5w8PWDVBd213ZL7to61gbzX
XVtL94t/j4MbvIzPV37Sx7fJm3yJ1TFE/GHrdRtskXSWh5yR8fxrgpAZC353XvvoRg510Nu/rL2o
1+a2PSVP1g+cqPMVA2n3i1UletsMITiatL/TvXlqhTON/2jKkXt3Mg6hgdeYaaFJfRdSKR3iA11p
aQZVhyX6K5seDX3+O2BwV0it3AJQ7s8wKZRM38A8kLZElH+rkOQAtyulIRAL62tYnh3cnzxhu8bF
kFEqESvQVPXkimhiWcPITYBf2HpXYztmzx+OSDrzsoq/KOHnPTNUvmnVc/XB/4998kqzUa15Z6cQ
em5lNhUQkYNg9I2P/S+Q4bgYApGr+zIyw1nCMT/AQbtHmDbzXTAkqp1XTXL7p0j9no/VVcSZheB8
F4onFfgtGyYNGb0zeSp2mlbclZsGmeEGFFN3FBg7aXewxSyRCwudDbHH0qBcCLnAPfq8rufwh2J6
8ljD8XdLzztYv5s8qTG50xUZ+voE/MGoS840MDybVkMnnf7hj2h3CHtuM620VUkYAV4RJ6bADcVB
sw3an9MSsjv0JtpPhB7+Datk+V7L7ysS1gKozeraDJVwj/fpErce8jXh3EDVm8ytA5R6gU1KIJmm
flECAtF6gA/8UTDJUPgM30VGXB9KkzACEHnzul+gZoVa08XUDBmcsN1YDD30T+spQ0KmqWxuhjka
VQeEmGDy56+zxhCQX8rCNvq/gAUPIK/Ly2YVmYT3i+J614NxyDwlkKOXqDadHW7NLwNdThKI1Wgi
4oZJogdfxs9trcgynIcR66Slrc3W9pXtrgP+VJ0tG4sXBacIxZzWUuhI5TYGY0dCswTjhr6krVgF
igRY79oiZ9wqRZTrUUze6Eh3oaxvOC6tVXfONIa92wuxFWjYmOaeK8lbm0C3/hAwA39d9849cneC
9Dwt11LsBC6QD6L7bFewtYi5ab57jk9sLU0PXGL4RLz1j16UG+ZQCVXA0h2fAgUe+62BbV8QJY85
PSSReLwTfE8u80+tNuBrrOUt9RgM2W2qb9sPhvjR/1cH5ZHFu4Ahlwg1W9ZUmvEDb0ePyDJ3Tf5O
0B+QV7LEDshKV2fC6KD8k1xbB+o28LDRXK/SLzPSHzwAcuwkS2o2e9F6pQUR7f0ZtSeOCl1+0JTB
gIcluAOWTnpuANvMiKNGnKHNx1xMgiTk1NNdkgXCjL/x+l6xgyTqQIyAe5PEKvecON5sFnnS/wAd
gWd5Vb7GJeOz1bwt+RmyDuM0KhCxDpmHfnnU9rARu+U7jyfBtxBz/T2hnOMZEV15KVv3WXb8S0pm
fzfQO1U6ReOvxijGB27yNL538OTR6ubnvZZeoxNZ4VNekadRKHy6tqiKh4AezLBqDeYEffE0i2wB
lM+uX5cCbgbjH2BHBBn7gLyPka+awJg+fTILrOXgds0IxVUiomS49/XNZfq180qZV3tiwofzQl2U
rBatLz3XC32rDAKmeoxc0nqPF5vAZ9aM2bFvyCa5uZ4Zc5G2/qeIK+L4VIqEwtg3E0ddKsd8wGAd
exJsfj+b3ulkFMCYU4886BBgBhQsr2Nql13ID25JoiiGWV94b6bpSHXAHxpEjBCk84eTIhPJhWHW
tJJxNd824JXiaIKIa30i1mnS3TlRKvHASaR7I9Lw4BwtlZ3GwdGS2FDS5/clpd9tq36stS0PyS/0
8DjxuraH585+g3Iovx7WTo4rKajZlrKNrMkXYLZZ/HIPJpaL1n5W6q4DWlbNVpS8JX7K2GLtMsG4
ku/gLTPar9tq+5+b9gPxukDD2Gh4j3005aAz/kAnSVgWfFINuYHof/j5BVG/+608Yf3sB9MkfYKL
UmQUESuyH+cBzd84XzSIvTdbiMH7meE7yjkOMEfYPn86u83+LtQnlvx1HPO3gBSgvhAjrCht+yYQ
wsPmOPb/x3cvC7my8xAw8tK4u9R4b6xhxoS7lQsTW3eRbTgcbhMY4rbi6AWOF0aIFUhuuCEiBBWU
avLSL/M0Sc3r6Uh4HU5FgMGxP/HAGH3193VriOsTJwrf8PM2xNAxkS4bc6ghthbOc79b03r9fcdh
mCCuY2O4mmbn8nyoeZC64WmIVijrEj1j0+A2Ll9Wuv0MSkAvBJd66A5gIyEbxV7gtDa4MBHa28wp
oQRTezpA/icn62835c8X2QmQkShqQh6m1OGzVAVXnI8KDtbOkzNpKDfZvKi2HPwFcYSrCus1bCAE
5pYqzK2GZEsHgxEjrbtPCI1FI4ZEHhaRolmyyXrYwS7EjZoz4hjzlwJutFaDn7tjzCzDiCJU9R2C
iUvBOMxNbVvkCw7NtT2RDOPurbtLbbzBhQeGIn2nvqSI00HQAgNTgZzy+GMFELcYXxX+u4fyPeOM
Gb9E8i32/Fov0B1B5k6naZvJ5Ax6ub7WCRLM7kplIPgiapR5iPZLxIRluVx3fTllqcMG/q0Bc6cs
5pryCuTlNIpA2sROmcPs7XMrAVPG4h7eGSPD3qtiKD/AWKPeeaFs/dofuzyv8mW0iB4QdQWpA2/T
ssZnIcZPierwac2InGDQCTHqd1VTFj2lyeI1N/PVh+X5bLoFRZzXt2xbXeeCv6FaNZgkyKf46ELk
TqhDay1MQkskaZs43OAhVpJYHctToe76PDXHQSbZMIQHHniX25Rx21GeOzfuduivb92/WerZy4No
/A3qGmxfKdgeTYQg8bTZTKHK+x9l6h/LvkIbWCpJV1dIEOuJ2/LnqzIFaCVA7c8qxtgDIp/2L0hw
qvMKGqEh84QsoQQlnhefUKmIGmMXDrTjqdHQTOsfZ7Lc4qoeWXGDD0eRpBHBDWbyf5FgztANowPn
f+eLvk4/VKn5QF8245SRFgXu4HFJ9rN+NCB1oIh3UEAauTdLNdGwyuNgJDiQkpqZKfnQoNWWnMfJ
eFIiahQNyP1i5sDkbgclGZ4wEV3jG1+fhlFA7QTQTlcGhwLJiYqEqZcV+zc9BmIeyd0Zhf7WMgjQ
vqElTQR6wR9fOSjOdSgfhatMHGFzRFFUTGSNorM9TdbOl6129jaIoTIvHwk0p2HSuWPGt5t4PIJN
CvjHKvTu+vmztXWum42vk7g6Cq1PlmwTnFzkzdWBGYL8N/jT7Xb6MnQxT94s0eeJjLNS236B/QfP
RGlZwnto7YBczLHtRhLynZ8ygP9KrQl76nmOpkbJVus+vDqlu/Akm8128g+3T0Pqj1tnnUoKw2Vl
c7ht0DeT4nyLdfdNmoddcfp/fGMw4ti9DzGzNHp5qDtq6OgqNTL76BMEk8J17A42mkAODueNBgOE
x4fXMYUvpYQpDUr1Qwlh5EfyLWgYVNmaTS6ZExldnvMf1w+wRZAEXYxNnfodGHNQbXQ/0sBa3tjx
sHPNXI3by96MeGW9cw0rbyBcNQpRLLFpgI0Z3SToZ5DOSv/kfSOkOUDlj9eqKkEYYGBBMW0+zD23
yWiT3wqSbQpJ9VZXA806TA4lpaPnXAIkEDb4alzoBlVSRq80nlXOTFxfStYVg7SSQ23r6FRcXvsP
JHU2FRYGSa53fep4oiiMZG6BvxCarJRuOTyXZ4D5FbIHOKV7rgmy+bLUdAM5QWeUk50D+LrupxNX
CRiQjhJzdyD4/kJtMJzPNdk5q4PZypWhNZXJ+4R8oQpMXq/KZDX0mRj57X7VlCfAfsvo+tb23VYS
07BIf91uEzroznOyOW2ws3XdCMZHea/fZ4IYDnLaEy5iiBqYUKOoPhAQif9ZhpzcMZ/yaVNwOkkr
cGGVtFkudVxr+4Vac4dghURqTuOc8FDJQFt2UrClmr7MkzyPiRoadfoRNMoA2frmc4sR0C8l66Gl
2c7dAQhmWQawHqaj1mwiy0/QmZf7dG1RgmSPJQ6jbisIFMru3zVmo/to8YkVrXmntYG+QGxtvMLB
zX4i2ldcR2C+4NDFeMu5ks/wTgVO7d/pOGDmdfpu5ySxwwC/3YxnmsEXrIYXZ2fiI7bNF0+UTLMS
k/4Qz0bgpWzABEQIxAfS/NbdLzGsh/RFItsQTyjP/3OP8n8ZjNIC/gBxEwlckfoKwxApqkwBvbbp
rmhU1XZEHKEbAuq47fPCLDhPJr/GuJxkxKUuOsZjgQM3YiKVTwevlfh5tQggkm3dQ/3KRmw2DbUu
2gBvfi1ZoI8mtzWbKJYpEIuQAq6RCVvbK06iLOrtbK8fD5NK+qxFzv5veue0pPxSilBJnOL3ZcS5
Fg/1E5J/37Fg0INGmXpYmsZqMeMQGSL8ZUjDtcxrMBQnCimuIeR61whP0fXYQ5xm/gwkp3gqE1bf
KNOVJT8FUkdnZ7Kswb/rKb26xjKWje6Q/N8vosMeHCqJIt1FbYL67LyIu3eIo9etZ/y6W5iaw8e3
4zw2p6X/ERU6hWRl7OevU8wlK9m2FdAEtp7OiJnqYLpmYIrJa+kNhMy2sPGsnNUw7Qe9aY5v7yZx
znb9gcDcCYIyrRCAJKJpPYnuTIiab8HxSwYupZJWAmX4AkuEFKHyvwzr/uUlZWj5FfIVR5VG+ttJ
3oFhKwc5SG6PiJhilfUqhM9bOfSuEhPracWsjJXdozISPfFwjmxLzfah91b7gYLK59DpR+gClgZO
4EN/x/wlmN6Npul6+5R/cmTpfdXSSSHG9N+uYnLVvwRUjasyy8UcjMDOHVkxHIkMI8BqzkCtP2w0
ji7oCPVf0jFNYU7FrDV75YC1ClYK/5+dwZcVE//vvfXm2bF+0ku0i73PVa+kbVxw6wgpdya9Dkis
YovNrtoYlmrMdQdPDCDwBF2CTY+MYDG8Ex5FHhPdN4YFeobHwuxXWUpW9qtyVEci4yFntXGVQW0e
7UAz9fzPNmqHvcobyKchkduNppDLTH+5qLUgSKRF8WHjCsICVYFcnBtzEZ5WZPd+nWcyYi6Msgg2
U27LIFfS5SHhaWjIOmAk+KSVE6TbLHS1SpAZIyN37QtmcVqY8HEqLYdWBBXii6aKHhOuWufx4Cq9
/fBvow9l/4HnqwHl2JN9L/SK305N2xZfcx9qHuUf21rKFqaZpCfI2W1P2zuvJzoee9IhdrCDZ13d
ug0Bg6DyRAvslJJS/B0pbXnLlRKr0zY9W6hArsq+J+evxJlpQI7Pg33vj9AxW33A0s5PLrrnn+BV
WE1g3ORixD1f396QYV9xcV0MLwbVvROqrJcvOQmDKUzlXX+Jr23j90qizr/GD0hwxpz45y9cDYSI
la5zA8IIC1vYijBgr9QYKT0pJfANH6znbnd/3vh1Z5LKdDRokveYkq7MSkQCAiLW+Ds0oymy/4r8
Sjv/j/5+7puaP4G2uI2Pr9nh/CRlRYg46BNVfpM2mRIe1/qBx95uIJ60TIYDxB5d0J3pYTmAaic2
CRt83+8XWc5AgCTb5FWp4hBy8JbTH+BGL/XwxKzi9w63kWmM84HqMGzS8ThETwA9Roma1Wr4pKaV
XH6U3cug8X70sJfLOJcoUmsAL4lbbvWECBlgNfgQPb9PCFkWA/V8/LkmyDF64gf2LiEK+J2ujGZ0
kNI5gAfa2pO2evOekPDQCOybaXeQFSXEP++iLgOHAYjxkM0weXDzDstxu153Ua7eMU58wwNe0NnA
ucW0xPe02fy3qrU1b4eTHUYeKFmkegNAcJBOIHLO4I32A81u3SvcrpeJc55taOBf1lQfLtrWq5Ln
3KK7UiLox3o46RG7flbwQtcP+i7sXlp5Se7toO1XpAUolEwV6e1++xW7BoWVFWZVkKJrNSvIFfZz
GfeaSOBeOlejsLTyWD4NPl5bVXX0jhGD5GngRQL286/RmMu/RGUK+8zjCLj9B4sE+WMOZVdKjF89
wojmCuyogfL+7o3UV1Bd+f5/ribBODqOJ9M4f4a6Z2wyCv1xPGod7VdxGbUwNlM4UDwEu/ksindM
WzMLvcgQeMFxQxNTLlRW69J24KI+bJz7zsgbE0n7DeKWqoIpjg5pkJ9hhQgm4CXioEAJU30vGJS6
BTNGoGnNTkoDhVyz+ffFUpaKbE1VR0s8Gk0y7fynvbYSZ4lxWEHhpBw83N6o7dXEucQYzcM4qQBq
Ob9z15a58/O74sAarMsxNOurCDtFzU3kUEvL9Ji6W8zqhUYNpom/aPaz9xzn7jPM0UktybX/v4fV
e/jkyGDI1JSoc5EiTmMwlwyKknFndGc32EkVAvE0ZHuFLJUXZRt2+bRT9SptmjBV4XEOfe8Acpbm
XSFNLA0eSKtml8HJMlQCXM2iNHsIi2UU81AXq9F7P+wzJvLO5sBb84BWkdEGhrh+i+vnl4clKkrj
3QRX9ewmYRAMgAY0060zfoGtyrzp5ZaqQle21WcqgARqj+OJCQcP3ai9RkbJyzpidzy+g6eokQeF
DXc4DW39D35/vcO+opass6HzpUIWrIu0xLGNkd/ne70fqC7evzxuNrKsjpT2Q6FWiHSBf7aULH+7
l9cgKTpb/mC6cgpkbnOQYla8cZ20BMtQnWF4vAdC7SjDRxlBByMnzTReoHQfIBEx9ky0b9pwXJSq
s10YopLIsyItJXxbNzV8onas+7oW4PVB4HciBgo+aTZvjeVGDviCJWU/82rZ8jdPR9U7MeyvBRaB
D19JHILSCOyGWXgnum6OI1pAexEpFQX0NxrpR3JKNAi7tdxd8FW6IxhlVmtwDvTy/Yqn+SWDm7u4
Tb8+cI/1nykAclv6dgq1X0xQmEH2Hm9x0Mpaeptbmzf1hAbEJEcJV1+gkUIihjhCMWaLv3AQEG+n
tG9d9LVHMcCrY+jDqv64uumvSKxXfn+H5Ku25wIBgQzREvCi/yAlHqK2i78xkYNT/WRPAjXWmd6F
i1OcEjpmvFz656dvsATMyH/nY0Iu96ENRYCZWVl89+0WT18H7nVRg0j37v1xDmzp82EcTqBGjB4L
i5Oi/Ifu5DcpRvDqAQByrG2dWFBpzOD3ryJZk42ZR2zubzi8dxFWB6YN4YNDgocgkv/Zvp4Y551U
GqDwMblHO37nZtZzw/NJ9UDMpMMHKgFp/TpGU/Kn8lYU3DkBAh8s37tGhndwZwbOy5XfGLWN+wAJ
BrNzzfrulh/LV0LbGKnWdko7u0L4Utw3FkfYj2+kQ6uKmOazP3aFChEQVIwpTAWE7SK3DfgB/YYJ
Uz+SMuyQPRamZVsObz0XI1bdjdB6Qi9y65SZVWPnlqpw4iRtFclCreuzVh2INKVHCweXSL+EUsGA
qZNDIRSVG377/7F5JLyY54vfZUkNF3KM1t6S82ku/2ZaXv+R/m+MZeduswKeRndJUh+SP1KjdR73
F/O762r6p/srioJQeYjqKw3fZHDiquy1CyrBY7wgI05MhYnMrO9YXYWSgpTvcy7qBzLxqTHMwuJ9
PHi7gxZf95WLvCTz9Ob/u+3P7PkHhMWDV5MKcdujLBuJbe21kP/RPInmjhcvj9P3TRRr7/G5Opip
W98QWxCHC24UszxuCMh4bM//wt9jrQKWHsHes+Ndgjq1SAal/F1p9jyVc+AIqh5JJy2pDidoow1Y
2w/CttLRZz6pHFk3l4Gxc46tBSVdUKP4IYK43q1h1ZtuNtnplqLtMPtrgWPCvxRWwXS0/W+Hpgo6
hDot386LCBvdpd1ouK563RxA+FGSccuZXijgI8l2L1EQbyXa+RTxQKZTPZ6eVgqy3SngVhtZ+WgK
1GSp5VX6zqUEObH5dU9eu+75ezPsCcLu7rfNsZ4/OqlpFa4HZnLfb44Zbti5QMwXYMBR3PRgncen
reDVkhaIxYnrvxax7pLowmnoSmYqi60Xch7gWZ0jyQ8DIuDZfINcuHdOzi4xSVm9XuCSbXIdc/zi
UT/05RkBUYX03ScGTFVIpRjcn2h+Tc9idRJDCa/oBYsGGvJbX9jHfhWgvG0YMBnR6+hB2bzT+dZQ
kc459TaLkua/s63heNlWGzo0XM+/LDWP4nsrc4kD18TocvnFEWFY7xIii4jfdm4stnXf8a1zNWO5
68OfCBiCJ1/Uro+3W1g3mBziVwTh+tnXV4PEZ2eQhJ621TsHhuLjeA67owtktn6vc/ifdwpGCGjy
tjG0cU7QDqN1I3G39w9Pg1aaM3oMRFAYjeDb0DwRD8B3AmlwgAK8h5F73zLzqCwW2H+cYj72wI4R
M5TZboP19ixuuP/aJZPIE+1pqX9Trb6xdxB+Utzl9FoCZzGGDpZ5S2UsEHA+2sMyycEQH4uHjYZf
XPy0bQ/d3wZ0CeLKHgroGRGuTRHmo/Ciwyb/hPd+ykjtfpvHhgJEQ/yp/5GPrn69VvZ9o92omj2n
nVzuF27Af49EfesLOCPtAC3ksV3FueCXL8QaRHOB9ENimmiYEPR6GrUVvMBaOXq9rXYRHQSZlgau
Wj2pNT45pH1gULBhpZ7pUND7X5S8viMpN0yEoSg2XtTZqF+tGPb/54oKKq+G840eWK9y9IHYD0Py
8Zgek8Yn/Od+ve9OoeVGqaIdGu6zNvg0c2abxzYfD/Zstj+7hUa44BSDxsysOk1EkVXqR7oAmV2v
7/HUf8XeWRd+58ezp2eUTj7xkTg38OSVLr3iutTXTukobqfnLlDfjbdaSQ71nFWDrRo12Qd0q96l
EO4JFbgeiG8xR0kbtxwhmJcdpeIalR6v9dk7qZjwGp4YJLmF2svhGBXTCyBCs293fcsMDgfETpgr
Rom5u9wszEv79/JGJt1XbSi4rlYRpUMn9Hh3wy0+o+xBqEIIuSIa1Q63QCfD+Y/msyzO463xHTJb
EgNeENddpKkbSmPmyXf8l7I0kDa82alwR3V0M8o2TrbTl8wTMJIdc7uS9IZf2FZBehw55kqoVM/d
XVwpTn0GrMYP+uul0huFrq6VSkf+qVrP/EhYxqbO8qrJBWrBBFGGKxavu/DvPShPNhHkuyArTXhe
SYreS9iykRjseSzXBfTKyDwe8OdX7K3OtRw12NMFbtWwfNQjAurelOrOF0AaKOd2lPaPiSvLJZDb
dk3aERhNjPTmMyp0keHnmuzedlDfdF69jgI3+B+AN8uLpQh0Vsqp5rmljjCgkYZOD3WThS9+GnmT
el7iVyJ2a/EDHszOeSyw85SwJYkfH/j2KJhYFlwbJJ93RYBHHKa6yg/ft+3n8u3TEiDP64rQTwe3
4SmkX2Qir+Iz/kOYbb6n6jsHSWJWfS35cC48Xq4eJVhgyRCKk41eOnRgBzW0FKGAd86/iBhyTi/s
2R75jriVwugXMs6oAehckWdAkT2fQQll2SARAcQKjHyvmY8PUN7quEWM5GejY3V40yONPXfkSXOQ
kpZpFW3GaDnhxyw7SVzdO/grG2PVzb21XL8QBWrOIjLJgmK4TjGxndAplcp0c/ImI9pyptVZl0B7
pEMxH0ag+YrAjD+oBtLpAtRv058oWlDLIKeUauMsgt4WqnTjbJ9+DFdkoc4g9wVdF62lS3CMz02M
aHO62n/bDO6SFe+a8Fx3deo/B/qErRnRjmHdHd0iaY/JNSarGens13rRMZEh115aTX5FQFX/fqs2
iJLLVhPNms4tJUNwV2Vo4oCuaDgC0GxnOhf22xyA5ZR/vt+aoPdE21HH7QurKWyqsmZ1Y2IGyPxl
4sraWwKQVOjVyzakUzxBp2fnWUONIj3TnOy0RbUKzmwAvIrjaR8MknrprTq2t4E4ZVZaluo7FXaa
i6EDS9kdKaEU3oLqDmGxnqLUrRobsAx17hqmoZiiFlT7QGIYO+LwDMwdJ1GrHLgo634Z0KGRsdDq
gifswuQ7D5csqXtpnTX+IminndFL12mxA+PadzU5D4wMMiimfLmG66oLYFjDi1UlHm005lDwog0r
iP32pyUK5iFWjU/nEh1k70vLfZmUiRmrmP1foA/I7V7M3GJ5CYB1/veF83IWRxntUOazHA6WxgCF
sM8fk3DitqOFLCJlGuVujgwN1FuGw94/ZvQcMdndvpTYM4yb3FGalq/Yksu2x8mOKe2mMWrTKkYf
jIPWoC4ipSA5ksFLqw4OWNoEz+BknEuiL6OQZnB/pxozTjc0pTSukYGTt/Mc54IbP0W0kWgYhO/d
e2EJ6tvwJeg3aAvBDR93nM15J0Imbh9Mz2WjNv2k8crSpzvNsVE5uCU2a8HHuc6mwOhezERTOO8T
ZNkqYv+LobsJ5WJ+97Eukbmf6qn0lETYlcw/572lL78eSJawGfxJn3hpAOOXydY/EXH2h1kjCeD4
PRBGNt/sJgWMltUryP2GLo+yAOBLByVVDdRJBENqvVJ6sLKa08k38wa2WgRpJMTC5kNp1RmYw2WV
sawyJqBQYmKVL94gnghaR9ok1zjX/hJkw+UiVaJd4ktF3VrV8eHT2bMUoysr+lvkkHGXvAlv1S2N
XqCQtfmsDlTp+PZ/w3ZiozdwpLLlAliUeipOpT+f6sXgRpUG2AIyydt/PPbFu5vyOWOHSKrtKrjC
x6ZgBq6CbhkT9Ln4e+Yfx0Po7U6SEAyDXffXKCYvstyzC+9a0GlHgg52X1iMdp6OC85iZU5M8aEp
ar+bVa2PObVrYyyFaQDE3ZR+P+gXNYSN+B+PFXjNzqdnjOnyEFEoDnjOWotEYfUYPJEANVga6ENR
XEMyqmdyRFKnzjYiELaGi1pg5uKlog6p38TQ4VkKTaCBNYlvkxQT51j+bmuj0+nMRJiKPth1H+Z3
YtZiEAixtvHrxNxlu//Oxqw9e0pdv5uoy30NNboQwijgzniwEswuJ7fD00uEg828M7uSdQdqfGHe
5NrX6UF4aJX4NsbbphKd2lQcvxEJSa6hZ8Hc8CqcAWxMi8M+Adbpw+4pJgPizcMB1LCL5jZBRDDf
sSo+v077cF7H3qbEI997aa0VCD4xTr7J9P2ZpmZAmQsxGIgs76iew7M9ywwz9CFe09DKwU+B3bLI
wUxBiy6SxG8p7RsfWm7zZWxmkArNf691DyhJ1R9q+PNdsaog690qH597kaOorKSwubVjRjeMfL7r
y14CWpCRvhAhPWv/L3nLdRjar6vo+DoUFRDSp81KXOT6s/O3OuBsz5kiA84RXlKaKpoNWZ5UO4UF
qGAHgTaQVj2JDy3RqR5CW0MsjKg+2f/L1PXu4VM1fBwBG4KJfi6DglWViMmgBJYtoJFNm0gjpMWL
zwofzkG2h4GMCg1VyXmZbFBsIUVlLkkRzcFHs7J8/jf839mGR4BbPH/UXAOXQXwvaACyOPY/rp+9
RV9AEdJV1ZIYKilG1JhKLoBESUH9dwpUaMVBp7jNB9ZygfSShGMmKaQlXmGCK45ks4tVSL8WzYkE
PbwPhbjnvLNunEQCZkKo4brksg5Hr7s5TLMu9o1IK+2uuA8VkOLU3WJUIfRv5u1lVh/57cwT4t0S
dwH0qIHAiRiwnimyvU0+EBNKkbYFv3/nnuueX8k1TPok8h63OaBmrN/n+az9+LHz0xbbUs/wcGRy
Z3cqbLsjIFxMMu8NHe84b4Q9azTpJk/qwEPaXybZKwPz8FKp604nYdHz0nPZJE87OYF12uwXng/0
qggje9r2Wfy2q34JiTaih96A9s3R5Dx6wGBlP2EWBcI8o38SUpaG/HKSl7KDu992DCdd0E+0nF+s
rSmGWDUSib+GPHdpRF+gbTMM1Jn7iypnLdcKZ/v2SWPUhd7RBqAk1qIhan9bRQWhQlibW6H0YrAZ
cUwAqEmNNuJGjie5+B/xb74b7RQvAqB2wh1553mIVt9mPNKc89RYM+wte8R0aGq51B6wBfhwdkVh
ua2T5ZF723t3YBrn9+9DOrx5uUeINPxNUPT9vH7f6QCHREWIiT+xjnaBk9Sx53KGFmTN8pGPsv3S
ZtKTlhWL20+DWgJfCEiZZx7F4zYsruHwahSg3U1M31OBSGJto8zqp20dL7VP5PTLlcP2N4br8U/Q
hTd6PWnFu8GhoLs966f1VxHCycVfXNHtmgZQBP6hKKhGQXhL2G2rWRb/jyBpq7D8zImJTxY/sIdV
rMBSxKWXUwPdjpjpZCcjO0JNwZ24euEkZ0skDta4v3hKGrI7bmamP62eAsxAueVmL3PmLqrJysW3
1fDAFs6/GfHyjVFS928b0pubo6EXyVKmHISdiUi1P3IG9PzBOJjIEedO3Q23KVdklvEfYkJUImzg
mB9ASkQIqH3lCgTj3axub7hQ9OGN28kN02FjKBlxWoIpIsRVlz58x6F26A5QU9ti14WSafFUMC1Z
Mgzf/MW/8hNXJ3xSVVUZ+phOOdnq3XCd/wRvOWfhuuMvnRKCJS6h6zPiQRp/PMohbE8TpoHtrpv1
oJkdITsYbPdpDdA6jq/Bs786gCDIT1KE0o9D6/qudHYKphUBvF+NZJGw9Yxjc5ZNo+ddNPb5RjRP
Tx3hMKdU0GUz3jqUjS3xasV1KVP0Ffp/KNP0unxrVceGPp7YynNuSB+rQDPCeBBwlNXJCyv1361f
DbUFTokIeyjFThfpJlsS8sAByvRmKTViN5uRA+zY3HJVfx48qLi3j9vC2LB1rphUKRju1xS3cO61
Rejz5xO5hz6FvcCMyXtZj3CNA+d6A6RP+y9yJGB7xGkrlw9r5fvFnsz/kaKEihk7Ns3f6WhkvLKt
qFTYgwIvjrZsRAujtcGc9HmsrDYyS/sj8hVzAmY71YtXnCnLSE5yqIo6MDczMU34anMA498Nv21a
KAnbHozXQU6JwEoCdyDsiMipc2lkUliET1w4gpk3OFJY5/5pJpdpvDgTULik1gSL0foahBkYnXIt
FLcDFui25l4j1xx5zTzWe0JzHZ6Y6BJSDKNTN5oLWOo2m6Yzb156lcRCzIVzlDzRpMm180MX1py8
T+wNNB9fUOYXfAWf/5BptHnRaYIB7hj7pkQ7A28qF3RP+M6+Cd7GedCvnBYnum5//OkZ/H9nI6oc
7Ihe5tXzvsPmKCQ/WPHMMSoPH7De5C+XJQuH4VfMJnoowV6OTeyT5jIofUP6DNgJ5Ity79ZHQYJ3
03F/Ytq5OFqf6DHGj8w0mLBE24Bs4okVAM9TlAQ8/JzZTJqvJ0aWs53J7r+l/E83mueTgOvZRKAR
KPR58EX7VMLSZqXCUgnrHhv2qtyq7Kt8X18GVW+vUCECEWXgfy5PNHIzNg/lZXuOLJYORCfcm7Iy
lbd5iPpheRxquVDdqcMmIutXuZZmV6izMq10YP9e8FCmQONWpzNvlq/SAyezNEucoeWv887Yn+RL
xxRpqUIlRdCmooinFfEe5fTRSZWK2oeVSneUsuyWzxi89PV8zXX2hlxjyHHBuPD8FXJMltm95rpW
ZrrCoQIgJc6xRKtMSAfWSojE/X/V6KBmCkT4QTdWIYNmphPxwklCUndUgTwPm+KNGBlnYsDE3MyF
Rkw0BzB8m2tw4QJ+PbuhHTlMhM53UrVtq6rfnJMOnf9A3cY/iQsJfURyz/rU6KQ1zjIrdk0TCV45
m7Fy1E45WStgajXNSX5MU1D9PrEg8CinDht1ka3xP0I/IyaaJoWQFPdklIfz5bKeR6Hzcz+tvqd7
IbppVA/++FxKFOzJOEZYTtuK8G4ramfhQd9KC9G6c3OsfSI9ACwYPWqeh++kJnKgnt/rwlIAhC7j
IwluwCwnVnhjeZwR6E+i5cIXJqlFl2BazNtrgjise6FjbZl1ZrIPRv7XP/D7NTS8T1tAl+rTNEn0
C62pKm7m9YzunwsIiiB7jBBXM5ghPGVbI4YN1ZUjCoHenJzxgjyCCCaWqid/we+NzFAEssq7Xuqv
7EXYbG+/h10sM06GgXWMp1hI+yMHByX4TN2L7G/p5Yw4+tftrDTmnDhw3h34xNY7Z+JzSWz4qb8c
6UCXtACmiB2tPkAoywhazxyq6YN/4SlKYHRIawI2mLliFxLQm8Km7Vpp6NhpEup7l+f93zQ4/7DK
cg0VQ2NVXJezBobo62WjWG4O7nEpjrR8FLJrBULBZTPbPOOJclzaLgGLzPFxkLKC0hBgTbDKe+ks
47rUdq6Fjr9YwRdz3gsmntakb2ikyp3WbQFHA7vMRatoi4EAmSeSrC305yBnaxlZp9Lof/R7WSeQ
88NCmmR24V/MlhJb0ee9zYixEQQfgWa+A20An/jX6BlCoXWSdQrCEaNvzTPkIjR+WEl9k/cUzSc7
1jp8L4exdmgqyoUN0gD4ii434qYJ3NpYs645zjQzYCLSWWGxJ9AbbO3mVXIZSDAmOswMTWRFDpvy
kfU+qc0qJyTuCf4XRhmZJCFQgu0/9FNoKOVb3uF6Qs6SprX+mETRLf3NvN/uXciW7GCuTTpX7tCN
oixVqdq74Ef4UT2ysU/aQrAnp8LQAuZa9MBQYVbobwcfZdPpACMYWvEmAI8xFPfjcBDivUK+QZzN
VD/I0WHXh8rzeRbGhIWbB7JK643XDrNoe2fB/cHSsZhNpFMTGEMPMvu4JTdt9Oxy4albiS/eIdY+
aDukPXhKDCHjaPjHiXUdby1oYt9SaNJJd8CrVhKEdp6aJXaOSqD8zffv2ZokALlupPt3MxDALDYl
LkDBu44Fklaiu+hSAXnvzL5exC8hhrHJBNi60WjZqt8SRsC42cYInA0qR/tgPoBVutQRdU+/dDcy
toOFDT7Zqc//LfgJbBDax+NOVvx11i95aZgtyHVIv7mRSvpQhb/KRBe6K7grWJBExMDSmy0W1ARh
2TK4q/MQq0kIeaK7hYKABjexaI/58Tciz3CMZXll4NfPqsX1qraWzgMHiQotv34QC5YTO69A2HUE
VuOC8mamfg3hQwkBu2RLtg9Y2G1WlKax4FBOawRhdwGuSPJFGvdjCy7eeqgMfcFqxzL4QyIz/8Uy
aSZ8/9kIFA18XkpxoHVM9ePs4mjpQE16cFQ2s9KHI8GbKbUEfIzpn/eW4IrGNCIN6PVS0mZkhHE/
4hJLBJFgVVATG85nBIe7qddjmfvdacREskpPWoMso+k4houhn+9cIj+BfBNcdYJLA/xXHtH1jnvK
LWw/75vaW5NziZ1HoDqfs7zXSpRz7b850gdseKUCptsa7IhB+yx+/O6FgR9Gg1BhRMa2dbtwdNTI
WwW3z30UNFAonfXChMWL7izpmf4l4c1m4bn+IIOF1DBVS8m1aH7SpbzVLO4uYzknO4qflnpiThyC
dZW/Z1KbXi4IRcKjbvrsoO+xITi4d35NNuAxKA9sYlhYlSNWwmiWR9xz6MttIbpfa18xUVYw+Xvo
JRxMpVjs3CGs9q5zpIin6db8o86VWpFCUCpU6KQ2wfNQtIhrpPltnNPyeuALW4wzMFrgncVlyAJ2
kFO9tTztuIjEzQUGFYk5cCq6vffcVGYlIGQHBxEcQYr1A5zKsnxoPTUu56axtp04/gy9vGc3CaNu
tjt9SC54d5+S6bl7i2y8WDNAjSNVn8qTTKzW7e0uuvxXCrcb3wfGG5j974HOfF9vrd8k4dlx1hJA
AGz/aOLZAuWFlNhE9znKRMo3fQpcg35ro+1znbmqMG+tOsmODWXbp4KnupmDUn1UZbdAaait+CHS
gTH7BFZwXlF1zafaGnmsnlT2lpBhz1Swsc0KO3sKfDeThYc+bOWU1RbwyWJN245cLklZnS4/gkZq
5nsV0L/GtPosQZ0OgFkhZuEaeyxzMxG8zsym4XJl8sG8RJY2rCu7xpASRVqwih1AOvbQwLf2jLWJ
mBVFVM8Myom6/uEr6xcRZ9BY9yq6a2ekFL6YB9WDQAPcL1KnOV0CuTVl0V+6ViY8H1xbXvYCecpo
YI9bflnqn8GkW4JHYG7LPcW82kdNsCXhwv8Mdl1dT2bYHEazflyLDfwl2qd70FWMAqEW22BvqD69
N9GXdzsK8iN739CSRFHGpl8gUuoyBK+kbh7I5+KLaX4PjiHVnlkwymUx2VUyEHoKdAj3z0sPFjRN
EgLNtTp2NJMbc+XpmSnFbBYGyV2dvtU1Y/IfFoBIJAA6/b+djEiEkCiAx9yTUF+1Or7nzKU9Gxcv
Esx//1F0fmjJrPY38FhmnXCK/hOAZhmDN0VM/3V0H6JUKfiwLGfkwocq0f6JL9nAZmTzCTD5/qzr
INYXRmqoqufY6I0T2o7LvtjYeRL7n44GzUgFE0K7wWWeVXZ9v/+BZlPBSgVhNGJSvCsSPeuVFj42
TmGCwDu8XEmOWI9NYfa90vTvVcQNJGIwEKIAN29eA0zDdcQfaq1Z71L8/CgO1QoqWswToj/f13O9
FY6+XJ2ixNbRPAMdZW29n1tu1ls4/RQQPQed6OaOv//zIO98+yFReGoiFSnWpe8abLbg+KEP/Z0X
swO1yS3uyOqGbIduHRJ6InlXqqe0SXFtVyfPxqMTKmLRFIGAOrn0CeoQeU8YWqsYEcCPO8E6avCe
ORvQtbfUff1Myo2ais740xLEqyQgutYz2Eyuv/XjEoxlwD21qBBgGHnYqaYJook9s5acsWL2A0jC
YYSPu2P0wi85OxeotQKvVV5CXfXpI5+bY7vVxhvokiwCZi7QQv40JC6f3fG2Mm6kFdxy0+uTMM7B
e2D4hKXsmNOzFhTpfYyiGnCnxfVJvclWD3Yr0Of/BEvZx9RGkSaYC7bi1/gOo/bJAQM1Y5wCjyl0
p30mMmt4lfiXAYqSSxXBS1p0UXpQeH4ydTndIaPAEv+2c4yXveeVDNYAv6k3uMAMwWcxnH9fUtqF
2rjlhtfWRqIPDU1F3B6pHmlm4afuDGKTNDwyKI6HNN3hcFKqzg4Gi7s4JtNPdSQKDlGxRvnskmUQ
r5CH4tLyGg0gm3WeQhG8Ofr6PXFsHZCy2ki2ZQ6/g+XL7ZiWSKWXnrkIB5T6PmwJCQPhVBMAnZCg
yY4ylofNCWJoOelUCYawDcEPe5SH/cHyfoKkRiMYBc+aXvPMqI/kZgNGYL1x+jQd1tJRvP922ZRA
2M1ttthWXVJArrEk0T/xDXsIYyk9y+PPpuaoY5JbM40P7WyL8AtUAbBDcRBD0uRLWV6NDJGMWuFP
gpprt4Sx7EUpU7CJKkwJ9UXRrUVmxG/jTo4cp8BJ2Rcf3FHBsJ2t/AhdGVkZ43Kr7jX1VcT0R+K+
a/ZIaQXkK0K7vPmaq+X1JLh/o5ppfzpUFtMNW81N+QKEgniS2er91NhsDYb2sllFbSyyLMN6AU6s
9XvApDGPCDPAJLA7bWFwnOzZ1HOPD6EccVwjKdvP0ehgFxl/wWx7VwxrrKtaqu71wpGbgEL/g3ao
0qlFaRF8VhOhJ+dqApsHakb5rMtdnPw9itGs3oYTZbrj0LNDwJlvadbMZuYypK6PZAz23RFQwzoJ
Pa+se12UGcySAXpQG6KvROmA/aHoxL0qISidtBaMlNFCw0ba3Udl8XiAyuRmhUygmSZ2mjfkaiuV
HFJncuIxiSEms3YQxIhiOQIgwWAXBvipnwvYNzKrbcvYVO7qzOWL7r5KfB0mKCXD71b6VRnHh3eD
BLE42VeIktCSFBEHEcdaAlNZ2X6tNL+nY+MwHWBo23Hn+JY/N98Tj52TUAlhJwQdiKIY5c2Jus8B
7mH7QBzIRMlx0o27I+6dUMUzpb0L0K63xYK1MKwN4tStznjWnRrmsUwtiAsBrUjLMBy4QOzjejAw
GyWVBDwMJr5VhHqYqi3CkoDYJ0XTbltRtlrCMDEi3cc2BKxEO+V/QteN67dX4+cRIXYOoygpcwyO
9UR2YspdKqvGsRxG/uCFdtKxHn/IM8zxKG3XBgvV9dEYnUipa0/d4qTyeTol0BOUJwxBPt5EdNmy
WARdV9BjOyCq23qKKAFh9pkB4gQV/w0eskYCohU4izFlZpm2djbqQ6kWAZhjIgHJFsP3vnsYD2ll
Q9o1Pw8Znm719oqtNtZzMR5qeq2OCVKZ1QQI512+rLmaZCya83UtP4RzdcJGV2jNPNfabgPF9bXL
8fGNuzbN/v4zzGfPAZLCx2jChyRS/E6DWWxflxEbH5ikRNSVtkpTGkhVmu8FF0KfY3ygZmWH+nQW
tEaeCs+l/pej4/opwXZZPQa758iuSeY463Ehoc0qiccES0d1Knd6o7a7C9tWGPilNpFYWHVUOiwO
Y9Zpu0dnkqmSE8LsuZwnMLXZy/b2ZyXSL8VVmx2OB1GLTpL9dIDNCIYhUY3In/3OvKj4ootM8v0Q
rzjbkgL0tn2gL5Rl1gKyQ6IzAXoAA/nR6wPojucCYvcyQ+b0W75ERXPosBPfJxGrNv+UKSPFvfoc
EheJZdRIWALu5pkeCSboCAn17mIYAcQcBlbsbX0OkZTjba3uPbfsfFgpz5r6X3C0AndgZrS/eBKI
3DhVvMV88Cdc+USBZKJ8Nwu2XSOvXGenNbjEjbmoaDmVzRTXbx5+AVf6eB0/YQIioRVIo170OPKd
HOaWbTtlJ4+5F413AdT7WuGUaTEmPMb+e9PpQa6yw9cqvkPBJFOjR/YZD0P4fmHStjiIFVs1NLCP
rjPhcFvbW5iaWMzXUNAg2Ns4iaDBwSlhuX96VYR5TFkqlVSJeWPGDxT0OyYIueiBukiZQ0pFlkz0
nu/X+WaTdPb0g4fgMd1rIWGE47KTIMenE40ujVGUGKBiH9ivYznu+4Fyur+3AdCAooEF0xh7mDWE
jS35Ev/FqnIKluTcPKG6couhc1Bs7FyCAzcYVy8BG19xiqbaB2QzBAc8jb8v/tRlb06QEAYvwHB3
xRUQtEyOu6TtuXY0VnFfkNlGjojL4iEBynlsPjzfwBi/DZPgUrV64rnlqXIATtHBKKBZhxAhtMoJ
89wS5ezPOeRdawiuqDW51+Oc38R0nLhQ8gJA7oO/dgKZi+RS+zsnn0fVxOSWRpHOIzytn+Wiam89
VcifsvCioKZ6xqbwttv/vACyg0/5AjQYq2QpvZ7/+Lnf44yfGq35K6DeK8lP61EAFg+mnnbylMFO
d1mrmCXckoxqH7XwhKIHJQJv+7IEvjnlQPZweJHRuuDeapoFqG6ta0PGmX1HjR33B9gKjECt4Vnp
l4fDOUO9WMvVOsSwblyG2hBN7N8Yy660z+dklrrwIqXLZHWOJ62C9WCO/VWOAeKXEOHIAvjo8c5R
PMPzb8QZfVceP76pi48uVJH1pqpEQYEOQroy0aKurmISF29HVLlAtGQXtlJRv0oAqFtum1k3bGoF
QAXfKUqXcXBgWELlStwCYHXlMJm+jTbIxgaKdtQ+iUb1LqvFbiVsPsE+HupwOblO9sORzSk8fuGb
B6EP90aDq0YcpMPXbtcUJLrvV+EtAFjrK83kgApImtvGWrd/RfDjxFr5NYvUP0RLzriQvcusIDvk
HG4awsk21dZOrLbHspUQZGWjunrR6Jxc1Df2bTv51FhY83NR8NJkbytCMRXCu+GfCXu2su/fvIK+
F+C0hz+pzcO/14MNUENQ/23iNJy7MBLAbZiTx5Zo9ef9xZMxRKWb2CH2XYjUnRwV3MhV3rrOSrlr
9SCzj7Pr4uxDuKPpyU0nx2kWClkOh8VHK2FVuQgFGT2fn11PpRlAw7mY2Ljk6PtLBAq6CUwg8zzg
78m7MCHlEugSvFEOVX1tyhDsNPfkcOyiNRBuetnoaQ8srGboS19b7xoI7AelysQn1pl0k3yjBxxR
E/Ng5pgrXOTbTG9E8tnIW8d/8Hf7FiZ0bjNlHwdIa1ASr4ePidQRkG7x/m+BkD/ghWU6S6xEQA0U
7n/UjVupCAg59/qtu4F+VM2aiLZpUad86gSM++o+ii3g3Xdmzrszqq3nQWtAr48XhKzNZsWxbxAW
p2XfkcP5kSfTjK0sBt03OzFYVXXtKZ0KWdK33mmO7WPLUkiO6UNyKOm/3d3UF14hqaZWYzRgOLsW
M61V0kRLfqeQ22cbIQlRdYJ37Pn9lX3L1b+Iq9SjCFh+w8NhAeaG+o1/ioAnqmnx2O5Fmu0jtMtn
q42TJNTThSapp7319ZlTrVdpdRZhMyqRPGl5UL3OOm7hirjeNOya4t0sBhUcQ/AMkilyHiytMCfy
iEiWcvfBuUctW3G2rgde9eE8uHEZN2MsrSCYxXsv6HmJdbLfTqbgcNYha7xr8/zAK6XKoRVZ4B7x
igIewmu+ICaGcsfI3eqXTBGz2eE+7vQ+whBXD5nV6bWl8taYCDPLHXEHD8U3QINYrw9Kunn7FuPY
xOk+ab57mLYubxADx4Rw3FAZZx9JurDdxABb/WEEuLAsPIqMrQXWvrUD7HFgXRgi5pS3h/VEArco
6bLxF9g7IfhPN8iEI/sXuYIGyAicnoIKw3QHwxGdFlYFMuWCmcESPGjr+qwsqX+oOq0mYpTZaY/E
8AORq94efdQ5ESF0n6arrWJWZinn+9ryCjashu/Gt5ct8cwr4baZLQ9RwCshubCjOsjgMfNzTJ4E
mqlHnYiJubUK14YLNa/BAoLTeb3HwcytNtOHQOrur+IyAgcnETjgA+RexICkVE8G8GuG6h0KseEc
agDgyomlQBQtWfMtB3CpO1ZEIakpuSUGNLQe8+lfc1lHIfLjXLyVcYfpJ8ytpE4Zpsyihz6dwzKM
KvNo06WDXab0jTpT77vObKYqPBJyBLMnAHEzusUp6El5Zyak3OiWfIxMd6eXfLWNW85D8hIWigg+
L1NDsJweP++B823cmQq/t9/ZJYiZxZ7tqzGVhOoYTgaZKQVnxkgRzjERS0WgMYketppFl2nwu7Vr
ZOhEHwUD4AImuYLNB5oHdlFsIopS1/H+fVRnuDug6usGs0SnS9zasN+5caUf4HrizbD3c0swAQul
sT+MVmAeYSJuQ/sRMRfyhq/b3SKxogDqBKfeJI8cO+2PvL+HJP4W90rdpwKY+C+NHcXUDuAMkryx
q0LnrkHw29ow7axEuyMvSBq6TUOfFFwAgbJYnXdDiVujYj1cH/1ETNg33toB52HugWxMDcqG4PAE
XlmJFdvRPiYwjZJv2ILASwCbTnD1vHu5BXvE7ZBG+UWVP4m6o2aS0izmKSUpvahcj2bcR3wOosyU
mrZ9ccaAIdXU5Y15F3w2i8zl6lkBgdOP+vyEp5V54DJFh7Dhfzyab9/i6d8QeBczM/lKbVJYV+LJ
bCxh9fDxX4e6vyr0883Bc2bM3M9f4PYy0RBxBZ/0xPZCZgG05p3590P2Uda4AQrB4P1ksQ2qxEJ9
ihYkV71RW0hwfh40Mjo/4KGNwPn2GNivvybMEPl82X4b4iolP7Muc1iSeasxg9bIc3Bd2yASHFAo
ZAVbSLBZLUlOcFpuGD115gkMKv70NA8OeLZn/TabYHxrYmdmW5SQaBRF+DX32QvwpcBf/83kiW4U
dKd5Xg60sx93uE7gGZb/q0LyFQ0qkq0MxU89e9ERCGM7VqVzq1LCgqYIiYED6V09om9kbdyVN+uJ
QcqoY9r9CK1jET40UjWEkgkm6/wVNpq4bPktYHFfckHzQe/VHnYp0z3ecZ4mQXvEU8XJwJSmCFLS
yx9z34hfmp1xlotgSlfgx57YTr55LfYeyZQHLrJDDQymH7VdJqZk2T6mVA3aKVcbEs5Dd75Hj7dz
OQeWVFHp5O70bkzBQNKogHvTm2cz5J8ApIZML5B3jdWFKt/HHLU8jn4GLhtW+S88h6lGNR7oxGHp
A2V2nzpQs8maPoxLzd/OvzHrM2p5mVUzC59AufbyQl31HB02to5i1HFG0RzppctU9ybaBNpAzI4g
6K8wPZXH4+uxg5BF3BnsFyCEQi/z2Mij5l+qhewEyGoOt6dM1iVh/H7wVIGqmJqrc7l0befM3RPC
rE5Jp3VDTtzws7eETNFRkLVHeu5iCn4MBmRa5RhXBkQUtroDsEcG0tJwXypPcenmMzT5HKHbU61m
Y25VJt5bDJhzNE69d6lZycvQryeKwYa1ajreUZwGdm0f2jh6VibIa4XplXwtwtpfs8xUvwlQKXFO
bt4NQDIjoMBzEFP1sYWNXG4pKaSSDndoMm5ashNQz7NE28KSyGKEqunSPbQW5Co6Q/PhQfkB/Tsr
BZ+5wLxhAQlo5IswqbBvPdGiPcA8AwIE2L+XQXX0rHcv13j78kUm/a7SkDgYA0pSC9k4nFRZq7Mx
ysjlJk4Do8CmUXDKf90oDXkVAuskAH4FJm+R+haLkUWnxR25YaZRkwBmoBcR8xaSQHKdItbR5zpk
EMS42g9iaealEzJ02HYiGygo1GbhCZWlQDFt8a1VuYUYxLPNRMrIwxAVp1ukFDOBewqxX3iPEYaS
q1h47l3xaWCyuncapF2OjyS6o59TEnihvUaOmQ7xv59J+1CTlWlH+lDpsAdajS07VQyoIYl0vsZF
dzTesEt+PIkH2FP5VRKQE2n3n4OzEpSFcsYRu2P4fLdL8nvrEtU4m1u+iB7yehj+L7WUlWhAJP1+
M12yfFx4T/uOdJcOENdiF2pO9OcOpKMKO0OCeFdslY9w39QugYO/QugPUEtVjIIkQ8ZN35J6ljJg
XDBBuM+Izqo1ver33nREtm03rH9+Xw81DOyHBbSCfBMnp/B6+c4DcXhDXpD2/i85Myz9i5gDCx6y
wMTsloUVnbg8KzzGwRmR3fVaPIkiz0X5uTly/kAYqDeYs3dDDwWh+QUFhpimS5bpCwBJ7ocnDsVS
6i1GpibbLiH/MJfjTTZKGReczBFbT8gv0dD/DIUoDLEosvh2MeyWZkawv1oDCJJNUKCCIvBg0etA
9djKLiiXiSq6V7xZch4XCQLHQbkv+Kv1PVCsO1WRQGpfeLk7/T7wFHYooJ2twXwkwmP5K+GUzqvs
hpckCtT5KvD7YYAJt55Xkeaf18ZJkFtAmz3NR6gVDNNIH69diXdqpREuZuZWQFpjoCaJPTHkpvaQ
P20Vd+aXYnolk2WLU0O8FSh1Kx4TVOXWmhhmTJy0KDq7LScTDRkb4v4rJXtQQmD9KXYp0CDV6ZwJ
gGMzgf2dKZ58C1r8qydsEhx0V+WdPExFbG/JgkFZNpueJvcr2uJFa9TpunZgdrNOuUuSFavcAuBc
o+xYhqfvDt8xmWxYSj7ilBqHqtj3DnZNhlRoDjVHv0jlXvDbB8j59AK/0B+kEiiceWkNRXt5w2Cb
Lrrpv/wOurNl6cZ6Jpz/pTpRYeDCx0xIVqMo7kzQ2dvmj76bkc/+c/As8n+KM9cKm6Xl0khbhqzB
ShUNSzAEC29gL6/9OnnIclzFk9xlrQ0dKnETffw4zbqQbNHuzJS1aQsH1cKiaz2QMRXuIIVJ4eEt
4EgqfyMTdXS09v+Y8dRj938cOM/+we5NOdUtdjI8K2XOW6YPmcZMqXdEwlrEcbumogaRl5lr+cS8
DealAPCd689HeXajI8lSzFpeDnL9cE46LQLvCzXLvWhtqtMPX6wzo6TzVJjv3ES4TTs056auS0+a
uAZEnrQciNoPhq/Da09DLyb7oDRxZPU21qO4HsMPGmp3lBEtRvH7gVyCf/cdOrokid7IXAkW7o1J
Ol0BjsIGo50SJ9hgFrxMoZlO/lyt22XTs++F2GTAGxyc9j2xn1YO56II4aLytIgPMBcJss4DvC+6
lMlRPSQGjFdUTcnkVWfjmFzk1W99URMHk8BgtjSHBTInB3q13Apah6KJ0oM3m2QUb2HiCm7GUNVL
XGvqrwSAvFV0XF3osHmMd8rw490o4LffRLGxzYpFH5F0fMN2mDb+unRS8/CRe7amMKE3Na8vCWq6
aVb8ubbFui+98CrupQbCgXizvvl4mbi4UUinXCPQ9gZ1oG8vM0dipClBlJoXmFSSdWIOd245zD2e
KF9b68gqD0AhoVrn5OmwZpCDWrfCHtJX4aPcMLMrSY0tzfBpzQ3jDAFm1n+/Sl4VHWLru289XM9N
xjMYorBt9eMViZO3dadzuKYkr+L1hqc+Qk3L30OXHccuXpQmNtQwaorqav9L/RIBsUMS+ZWta+ue
peJPlaofrpGKDduL4zeTmujiXk/RDLleLc5hpZR4csDFVNz57KavGhAFA6ATJa6eztJwWid+l3yx
PMO8+BzUHY62C/FgHNHUlAJoAKqjdyX2XPl5w3jlaG/O/diTMXQHS26c0vRPDcL5NjIXuneOvMPc
Cg0MfAgTL7kxkI1OnWjiLBf22URbb8vbmP6EsFAp8tlgRO+JDvm/b3mz0T8P3lzEkpQi6MNJutkF
+hktwcm0vAY6u+xhsaFQ+otQAt7WzAp96jONRFPxZcXkrX3dQQ3MzICXBJSEMzsm1XLzbj/oCcvA
ULrBO3GouLangAvDjKIdm63d5Lod3BA9I8WCD8IdBMB2dBmVZsMa6uvg6WOeeIG9wGWCAVZe1zgI
XSOr9YiGRLkTHqLjKAUI5poKWqc5KDAALkBcVz2efVQR0HYVV72+xoQeNC2kCE0uoWO8vNHQtS29
St7dinAEhAVT3XWf8dJi3Di8s+xXnLWiThKiKoKDtpwjvNPejE6eg2o1AjfpOiEzUzL/R/2gnoj/
dSKo3zO+m6qKM/eM0Q7ltkYtn/E3Khu/AKy4WrbWZsmhCGFHrqV9+BeKyjkiG9kb82PsxKxe1z8H
icbrfK0BJ94LP/B4Kc+XPnJh2PUDecnHfRWGl9XULNv4ChqB8lxX2J/RsWPJxzWdpLV5j79OYZBb
scZ0oFCNUy8oYUUXRCWjuNkvHmNK4j4H/+Da3FtmQeUwYduCXGbnsWqaPkhP2bpB9rJ9teRkxkZa
Uj0mfC2LwMdWuDNoTZFcyhakc9XEBsazhyCnj2JNBV8fogAHm67RRr4XNPGKWACizJrdMos9Rbef
Jil7YCj309cEkXZdNFKua6nEsauToPXfwfsN24fQT26dwgbpspc+wZqAx8+o+QhoMpt9TES3i/eb
Ab8/QPzZUECv9+YJeghi4VMtZpmr91wK+C14axw08kbBa80UvHxHUrwrplhszPZ3AuML7Qg8gctV
am3tlM8/NYoMj5fnPQ0HWR3ATU/9Jw6lHvS0fssmocPCfc1EeCTQfqcSC9TDeEoRE6kB7ArnbgiJ
EXyABOwbM1u09KsZ5tSKjVZ9ttE3auvCDJee1LnFjaRI/TPtTFJsv2QkBC0PipWGPoRKL3LdrcuR
eyVSCgUgbfjWJr3Co+oJHlRZE6yNz8IgdGGvo8amJ5NTXDUYeOGkJcrZxTjnNdKeQY/R81mXpC/q
/ZTMrjIazcU+0MvowghuI2Ru1ni7F0uX9sSzOJ5em5DExFLYubXJ2aFJjz/s3NTdfzfH/zKV+cg/
0dVPN8yTPsv+zvDBnH1oTZyN9tEuzno3QP39BOiSUVaFepLvKq+a5GqzGo3uoqR7tRn0XfLBiFoo
fwoPZKLzkAVePBfCU9veyb8nCBSACRUW1NDbvY5PZ9VQA3r/g/2Pd0/tiiw4CY3Xtp4siVLalVf8
ruZeVfKdmvQ6594DxRBOZzc4XNHdrn9kAZDe83sMY6M2VCm5qMmUAs9OoRjs3Z+HzuELBKHR5yNx
3v4byO8qAIqYn7I88VDr/c+46D9M9Md2W1dMcAy7DrxIhzEhKWvI/4fb+zBCS0yMfjFDFc7yPhc+
5wlSlcI+pH74/dUW6Mv+FiG19EAPIcOxJ02+lGPGE3asNKrobBhafEk5CzbF7BuHbvCUs18H/v1J
ON35/NG0DqtcDyiTF9Q47Tn8N0MqSiOS9WEBzM/fDqbii0CQzuQT4fdArqtXT5HvG0zV4ZjLtqpD
thlNQsl/7yFoWoGFH2AF1YUBct3buiXvrUAwBedHsV9Usm37mPSR1d+JuLEOocDkZt8yJNHnClDF
vO3NsJ+basPZ+sDrLdt3in5RlkojS75cVQK9PGd1XYhy7bydNOQILc/nJVE6LeSmYP/UHlyG8Jty
dq4ypaxvnsEtmoJsaBIIv3mnaY4UrhXkXeRjAL1eNp3ZV2nfCthYXogGWfJLNOI4D0gvAOLNKxx4
Rrkaw72fYBNlanSxpuV4jE7TbUibZd2XSSb1L1vj0xCA0U6YELb+bUPL9Klxzts9esFKpfLPOtDY
cCQMFO9yyCHkWhTu6a9nLKWkb3DDnZEOI4weDhI3uO0PNnS8MO0gCnlN8k4xzl3nf92f5uRzdADK
5sMQwH+dcul4A6QEIWxozEUgQtTqPLVmrdeFf2/WC9c0WRKpLuWJ7RP+vmvi+SCKDpGX2HNYRYpH
JVJQOGAHTgVSzhOyxVt16buspTncNEmB6eJYju2tNV/BB6KlZ1QmTOcxHBtzrtoW8E7YwX23wDqP
U8Fa1omigQwNAbHXi53O0d1/6XaIz7RwiFJ/PuYkA+WhhJRMSPoGNnyUgMj5/T7ZjWM4GjHlHd2b
LLuCJ5UnjE8/B8c4vLAKtJY57W+W22jQyKydORLtcmFAD1izROIAiGKCSTHIteXNJal3p6Yk22Hd
BpszmBacKSWUdLPTCzTGhU1x8NGl/doOTbsJvb7kX+GAoEtAKJog1kp199FQ/YG8RmUnI6nuFtpv
jcdjdAM5nQlXyf2jkfw2DjdaXmHWp0LZ9ANGFn+ktKa53iOTZ19K0DqBIyXsPEPQ+YE+9cyQcVqs
d/i+2xXUDVwy37JuftA9xFeA/luHg9MmRPuQC3dM1Q8sLI9rEeAs6zaONtQ3x9Qha8k0cqzaNR7k
AVFxI2EThJXO4u3C6dvEhKnUDIWHPlU1TMbb7BHp7ySGkpzrr7s4Rl2N7w3S3ncJlTyWxRAmhaUu
B6hnKW44IjnMgJ9p5LTGSy/x5FtHZMTwv6fKOB4Wh+7xkk4DbTJ59sJ1ljW0VZQQFpdJ6jeI3be+
J0E/4A131A8O8m2FZ4JP/70kq22f8IHaJ4BYhwGWcGg7AF1Io/pnGwQbA31IshW1gK2iDpDn9qJp
+n9Ubu2pusL463GSSmhEI/tKWy3U6AbHUZFz5kKinLC1auZ+jVhRkCoH2Mm++pVHV/R1fV5XjGoY
CiT+mvSE8eoPI8r5aG2CvBOYC/xycHfA0qQU0K2mmI2H7I2NkfViytTXtkwP1AS8CLaBsmzpF043
CqjZeVaD5zVNEGbpX7vsl+H7ly1A7XtvmNfi6jfaUlF8LamwJSaH0ZpYvw3nlggBEN/BQ/Wb4NPK
knFaouhFhmOEcKQjgijnT1suJwbU6m0aEgD0/D4JdLsvlF+ra2nvJ24GeKCIhhFMhbhNv9HSy+7r
+5EjvXvNyZjSHT8R/jvG2HawpGzyNKuRbne03JdHDcqnZjop94mhnz9B5TXhHjC1LADmNXuKt+NB
c7VeJiH6yjpuZu6cZRLm9zTDsRxbe34Vq25EYwhK1i4nt5/CC2ywoIIvA7KMG3V534asrn5BPBv4
ed5fc9mPLLf07HwWbqbvXqujOp4/duqLn9nv1bl3Tnm7m97ksPNkB+Ye0kaa3ATGcrEf02IMcYMv
VuiY574TXMaha8sS0RjOCunur0MfZA2/RWcTQmX1M8STKoZtORlfudDvQ7YOp8yO76SWTWj39pdD
8dWCcfut8Mk/tailsVTuVByXTCCCB28mRPSUcXVhxZV2zJ2aZb9WyNwp4UtzOkpvRVbtmp4tlJGg
rfE2B1djZfX3tNxY6kes3HdobIDx/kIc2xH5YxvOTMSeKaaTolLXeTolz5xQwACsgg8e4ScFZCAI
jGr6GkuTmTk6vEl8Sbz2vTl8M2gkQEtYoryJ0wK4ZaSuFpMYNue+obcjrjnNHcmHvl7l0r1/NEp8
D+yNuuHgDO5GndMpFVsAEI7v6iu3KV7ZpJqn0AMFmIE7w9ybezSiR7UxxZzjFZjnia9gwQmahF2e
PY2KRBnf3hVGWa0ApDJUGlpwvJqFdpEjMrVTywVAY35sz3bTlcSBl6LNAKDfizQrY4TrtHqEPLCR
1SSHvdXoLRbK444nCMD3QWlI5fjg6UJsEs+g/JJpOAb9WSG/QEEaJRPqW0DiM13lZv/wa+f5rXjH
dhJYUFkPI5G0U5lTmmhE9X6nrYcheTsOzS3WL68WTz/qev/lT5c8sOQnpJa2+gpOftclA+TBEnnX
/EeLyRPMm61eSeGT25els/PLKEVv2lKKteV8/+W/noBeXJcjCzOAMPQnqNRAuIhdQIuDkiHit/yF
SDGscoxc6xtUtyFKYpHfOFZOB1VRLiQSI2CQ/CgBi2oPGoeCam39bAIlGlGQVy/dd+DsDXiZX9fe
R6Y0SD+IAQX3/0SOLw4DdSHIzwuLr3A2IhXOt9aRM0bwzFymvnIg9VZOjvxVF7zyt7z1nh8oof7w
tQRtRALxDkbLd8z/xRb3hlwJDS3l/VRkWMmK9K74oYeAvMU+BpT2hjm4fjSg5I4vIF/sBnhiYxqP
VN4eRFIele0woqNy6hVf73hN9E7T3G8KyFVL5tu+9+g+wZzyxxCQnraR8TOdIS+NWT+r4Q7FWSSR
cvt3F45WavCIYZOmxiSH5JtYMeQ0n5tnIf1CxqHFDgGUbEqiCwcY8g5w4pKkIN35fjJlTbI6FQGr
csZjeoH+C0RkFIMvHyRJ0lZi8Fy3MZU8YR3+e6rlI/yfwyuw6EZG9tdEV2kAfHDyxaUiz1zYJauh
pHPVvvcnn1JigYxyMlqqmZO7OZ6pay+ZxO76/akK1FzfguiZSMvW4aX2Eb2ht24QalKxS4ato1Oy
+MFKTzLxce7lSGV6hTyeZgGcAig5yoY21dwSoIjNV9BWh9XWTGo9cybWHWYadgrJPkrN0sLpw1iU
Nana82PeBY/rUewsclf5+L6tW8IdeTjY/PjAQFVPSd8IXCq53K9Zb5lK2ppBN7cdodS9Jfp+LC1e
OH+SUWe3EsOG6SlO/Vu6HwmAx6Z32vvNDAd3TNkXo9kQSd8D4K5jlKfSHQ8n5wCO2NWzO1Gi1vwx
qcLGWTFNj/E/UmijtlUJ+eUPzx278wACrdh30CRoUoi4dPxIJnGnIbqt3pR6zFfpCORrkUz0ibnJ
pDGJdVkFHE1tgJ0IL5A4nUMdQuORsntKMJqtC5QEONrJcOF2iuOhTW6LNL7xm6tI4EZIn+gwJ+nv
4vjBlnfXTUYYsjTZe5ZTvg0WG32WNQKBzyNaKP7MScZGv7y+SDyqrWtvUc2XuGd4I7qJg54thIU7
fTVLUSTf7SIB5oy10faX3oLTZo8pFHqG9xSTy7RPIcZ91y11b/Zt6SeIvE4u9b2XQ9vtklvvOWYa
h8c9uoBaiGIoJqPGf11onVurOHPtAtlQEpL93PifxOeWcm0AB5WzS8VS7xc+jfAWWNUDG0gyDUWg
g0rWPwqOseNCQ0+CpBXs92T93+ML9wJ13nrALtPMnXQw53cEnsQb3LcS/93GAVMtWd/yu/qFxDkB
zjo0G2uWmBx+lZ2l241jaXI5pklN9sCCRNrHhmU9K8VpvIjiF0n88Itaz/Z2T1+wQaMrTL+4LvcX
LpVjgUUQU+2yq6ErADNHksJYytZLxLFviLcezf1hmdF/0sBvgMonWCzpAHn5yCIpP3UBhdMBRy76
rCFO2lemiZANa+jjMnUeEK9XrypjXROuf0y+xUqngiE2/V21kQc1nRngiYxnUxXj1JBbCWrWaAsb
klPQ6MXRgBs8g9sPzO3ayabv7F3A2a8LaBUbUflDc3CCFBPG1RUNhoMnXX7OJBuNDKH5cKKCh2mF
w2WVRZlN9wkx2VnIYQFk0wih8ypLeQ3RmwYJJMOVViljyBVc4Jq/Acjoz7SUJquo6GSt33FZ6EKB
Dam06x8kn/+zik2uuIFUh512T/nBknVYriB5Jd8T/d79F4xdcR9k76pa12QYLppgQyzuuNXyUFUa
uAvXgfiXfkm/QDfSm9L87bOUB+KOthrpsWKeOJENIsclTzC3vCbIU4oPBxhV0YP95nEN4ralpPcZ
dpYXdSA/MQS3NIOjRWlF8OAuaGHUC8QtLkOK12eeOAHsJOPsZZ9MI0GLp68ShppAyxUiZ+oZ3V+v
AZmi4gQT3ZcGqCWpNm/vJb2ughTW4L1mOww6AZzaMh9ReTgt9jF3LFTvCU3hgHwsfZbBs5ek3dLi
vtZ4zYjqQ73xlFgm7f6h4u7fN4sxgB2i6wa49d4th3gXyYjJbRtBGnjbUA1EmjMhlP7lBgwq4D9V
Qjozqy0teyC2AwInV7JJFAzbSSnL+REVAexegyex7EdFTx66JD199s4R05RQCyTLSt5RONHdvD/1
3odrptZ7K3FtLFQngyKui1FPyVt6BsEsAvUXDhkWxCyGnLSKFDZ8H+YhNx1pHnDJMBazknUj9hh3
F0XIMnWXw614EWaQimNoZ3/j90J7xaycsX/29MZHFgm7lROWwdqBLMqgL35qqlIcSMx6XP6ZkYXr
rvLfZ46NZa65c037BU0h+qmBxpfiQSTwpBMfMtDdnL0v6IiOaneZ9A6uYPUKcpU2N6BjgR+TcM76
iknNvK580StZGBPlcI6/F68NA83RDU9Ymi7l2oldgLNz8bXkWzZS5wqC2/bwY3ciFmD4GeFmT/qj
19f3rWOcKLTrwkcoEvIAcJckpp2kE5Bd0pj9ydLhx++4hNjG8QE6eH2cUe9HFlUQ239Tt0IMbYWH
zaJikyUfCtNDB+581U2NRLzwGgDdqFQQWYuM2Ubu/hoNIeUnR+hK/g+Ps/I997YRe+0U9L3OsK06
SvBYbIVICUYET4FL3UUMuFfnY2NQ2vJpqppMYQ6IWbvcZRjvkYi2zfEtvtDdKIBqcWGWBMgRcgF3
myHDi92X6btCZiLV/poZCM6amgl0USZTngb1v7HFo9PUBpdnqiOmXJmFSbGxZBM/92lCLAfjsG8g
zMXTBmfVN8Qu09+OV9xDbS2uk3Omx1IYC/4TpNiCt1xN9S3LVq/5qMQp+g6rcCeNYaZy63ox9dsa
9p8oYPwMkyqbuYu+WVVs7tX3PLhZtc7nX17d0mzdZ7WKOZejFXgh1/65+bnf67NwfR/8ZzzDCQjW
9HBT5K2U5PNRyJTaeeM/8Abf/YdAJ2gDIhnuZccZFgWxNLX15SEXwcCTXZ65w8GYBXhDizvZo8l+
g4eyqYJfuigJXV5JCiY3OFRsTU1VGiaqtAXbG5LssH+rfT/6TrtINabUOk1MmjMmmLifR5lKk2zi
ZnDFtFTXgBB6NNLjNdkeNEgmN/FXl/irIIIj7DtyyD+MuTHCX4o0KqQO6aeoagkClr7ee9Sav0Q+
caaby29O8JzqtLXBWMMBPozxyMKJ5xNYhQ/YObhNLNMF4qWRdGaW5wkaB4T2Iuovzik1VtXxc9vA
gslGPlKOSXPzbPf17efO/eHj3sc3tpieMaUfHsFcqq4g8KBwXIE3QLQHvuHtk6VfqSx+AV986Yxz
dpLbt+Khj5GD0WZr+RHO/jxqVoKklNEWl4uwGB79y6xy+18RCKZFh9MYQ3t+n2oHDP9SjGKF+9XP
KXPfXx8uExjrUIaZ766x4RWhHUEE7Yri8Fu+Tk/cAVYJrdsj7w8nEJ5jlXP5fJfi3rnhkHOAwU3E
Wz+uSvakC4cFgzdSNDTyrHX+TP7lSKL1Xh4vdAyQGq76HjZZmTXy/jcnHLGqGZ9X6VuGS9IumOJd
ixVMqRA1E3cXeXrhX7n5AegVMAeVCVxx9jhbqquyYjj8miOVOosMN7ghrOLrxpCMHmDFAJ39QXmS
cMa3sy7vaiTMvNFCslJAiSyNUWjcUCdCpt7cXHrp2HMJY+a3vRem8yRaRygLyZWya8ONhwCdJaqX
3wBY7kh1xyKa+LLzeeYP/2VnHsyq+WMWhl53ZBZ1Wl8crNu9OZDabMK7U2GMaA2YrLB/yN+Mki6G
XP0C4uq+U5YHjGuCxPk20fwSCf7FfVghsVxIi6JEoYwVQoQwW35ru8KPkaQUhPkFBG3sWQFoL3ys
qwnrBJp/Y5KXc67WwUEWcsB6ej5ydPDLmKkKkoGpqcTTupRikkk5CAlClLD98EsMoRkMHnFUsXfN
6APymVmVDL9ITW4WsUioSZp3Fe+0X8/JFsfAno9mVzW0buTBNZpke3qadRIGOwgIbbfTmHg+CIiv
TeKN3A2ehoXJS4fr5kYGuHPCPS4Vu923DwSeDpe/UuYxi+Pqie3V1tqyvUoeeLr4Odk0f+mJgDvs
z3gs8cXs0luxIYduSSfUQUsm2ocUiJVxy/tZNyedytqTKodBF7RsyYVRe/grFRhaXEPNCqw1bZxc
M6NxaNjAs/2p0dVbnqNKgYAwi37h6S4x+78C/MZPwlJBuKkWEvygpYwZS4ACKOoizLCjByNN6EOR
9bxPlEIleq5qcaM1j77Qr9KTKers700KGdit9Xhfh+QJCNKj9dJe0hyO5tQBAXCEfI6/nywl893A
3QS16th6HOXJACHE7BsqxkP1vLvAN5Ej3B9ZkISVOHdfhkfuspIpXqE+tnCGoaAi2n2NmepZCi+7
XMFskJWcTNDe6x8MiyfWDmTRCItXrAvDu4E9qAE9bhk2Vuz8gtK+pYZfrkTXVPdai5/6fWiPiC+l
p7LJvAOsdyMDrsctH7VmD6JZKMtLZXbEX+9PAtLmJjqPJk6kZDg8BoaYimToLuv8Y6Pu7DjKek7g
i2lvPTZrFLKMCw5DVGT9lQkfJsG2LQaBBgXINqjVaxT2ZZ6RuKWW99OEHj4mkDMJPXnzLWZf+1W4
lnAaRFpM1O36CxGfUeL9og7Tz6/evWGguEfh9+bDt76+ZEHl1AWGDCy4GPl9vhvIfIwXnTiaqWoG
sm3ajtCpRnWg4GenBL5/aT5axT1MIQgpgmoNFE12D93Baf73Qfmhj5aXqu45qIGcDn9KMJM4n6+M
e4Ob8vruzm7ZotHRKzyBd3LxVaGUS/fxVuaC8xXl/jS+iCQZqeE+2CT1vsAiPxbSVI8yJmRn0yyC
ct+oeVJgJ2wad2UiZCTrRPqjYC1Uz1TdFzTTMoBGdqVxpTHMC7Quj+TD4mYe4TnJxEpf8DDyAlyE
QASFwVLSNLS0Nhwyn3Q+NSkmGOzolcV85r6mP1zHrNkfhlrGobXgdagvGl1ux3W0SHMzLeC847RW
Mw67dHixJ170lDG6RdAsRvwhNA8pSV/x+jlviO3IZgG+QJYwQhLTeJHJ71SAecB+qqdJ3UfmYnux
OD3WyVZ2yr8DtEutdZtfxNj6n29iRIR4EX0cKkJHU+ucXMqFhLGsy1g5lb94jGQ5R0kcbdSP9hEt
3UJD61kabYBHZrmNsj64lXpYijpTxohW46r8gJHFr7uvj3ByH62HpVbVqfvdkYTgI+Hos+66yk8M
3m4usDmlakPup+pUjuXM/N70LGAUqSwlOVSvzYkAiN8tVsygGx/KNc3nU8aLjTJhiAxTygFMTkDs
omV+iWDK+dfW6WNYqZzdc9d9yPj8DaLscU2EvqQOHRtKqH13BxoCgwmHG6iY4DDnISDL1JwJ4F2h
l7kvMIXEEuFNzAWhqpTeGYrO4LWUyyNELBdkRbpa5ry9IbnghT3caLCx3ex09boFHPUbXvDNHo0f
3TNrQg5prNgQ2kKVPEc3IcHtknXqXTb6v0Ft0Fj8DU+K6QDgWtZ/305hFupArqYkx4iRmn/D+jQa
NBBNAJWRKIreIgWKeGU1M5nScJCx04Tsx4wbU2jkwU4GU0xLGufcA2N3p9yP88Ox9XIYkMHSjehp
wFOwaEpiDju5YqnQNxRBOeMgRtLFJATewGtWGB0O+jWxIIMMYTJbnDo3MIUZhMtes4oCeTJKdPmU
HF5nT7jd6DqtA/5A2ODRy8pzevAJuGECvyHCdzpOLIFHP9p0XXQcyvhgs8dRmxY8mh20eIOcYHIX
LRsNBp/5sTPeH5JqCeXctQhILS7WebmYQV/oHhxH2ZVVM0qe0KjTgHO0yS1+juFmKW3rtZx574Us
9W4DZDfHvQQVDSRGyMKMKMedo0VFBsf9xk8KfaUd45q+b2OJ8Lm0y/5Ssy9cdPF1JfWZY5qNvHS3
PiyspsLI4OxR/+ZIMpW3fhSoiVGY+jTCwlLnXnRuF5vYc4K5AB9NaQLm/1q63c85LPtOMsXs13aB
wbIEDzvOcCcs1bk5WvzvH3UVN33y3qagXZB3QVlSB9JAYq3BSNHCiMjSTv6ag1htulicpPZTJAMs
/XDQ/itfQlXxH3n1L5hVwYkmExUM2tSMHGMYiScA3BZo1HYY+bNjffH9yAfFLN68p+3pH+8p+1Od
nGnqRN+nwhTaAcebtXCFAX88Hk9B4J8ZL3Aq9Ed+8/deXCYVTP9hoPiuUkx31fdN/AA5tjk5EMee
trWRd0UcrXVddk3ue+1SLaaOgVlnmfqjlw/v+Abpkwq945LlIEn3BanKDPHcrG564AhUaKFDXHym
RmxOffXD+AuNrv/xpG+nqQd407Gvai7z9bAM1wbOaOXo/hcr7RZ+lyblUuwWZUTSQJiVTj56J4zE
imzPpjIyCItyQpMxGITEjc2Z4WMbdFlB4hr6WHh4wylOVvOm2KJsyM9sRYAaqP6UPZ2u3Rd/fsWb
Db+BOvfRl0/iaL5nH716FAOJ5iWLjak6KzkY+UNiUlNN/eqKD8LGObCWoRD9ZKKlPbWnv70tkokZ
iakQw84+0CmNOmo6wmeJTYkrDxv/zaHtcrtZdsj8tyJ65dNP+vdv+IfYAiGXRq9BIsRepOkBLnOq
eA5TlGkyNPuuH1yoA/pP0X8TlcFt3bqC+0Jh/RVsEmeBIrf1VUn1sSBMEVVkxO6jWUPsTEQ+81TY
ytVmVvvfpZ9A3MsDF+25YKCjk0DpJ0YkcOqIwZhR76IBXTzXoM0ErIXKOHCzXWSxgN0QvdI3bH15
YaGxo8bdSxjYP6OhiKw2oZggVWy1ZTe8iBuOesm3x29zTlcYWQ+FHxJBBcAW4R/J8gPqt/YZaqdJ
FppUZZMw5q353nRyhgWop9+mfiHUjP8Fmbpos3DcKkwpdlDUwLeZ+KUhwyQkyHgvkovMCdqf+ujr
nGnTVtZOwnbZ6Jbg0cuSC5kkEjvIz+eHEOWDW6/JGl8tl+iqIHKrZfwBvQn2YLt3px1+F7HpmVWy
5lNTvgY5Z/6FyILGw7BR6GfeMk0qWOkQcdDm1ClxbmucaV0XYQWXRaB7dF+Gt/MD5FMZ6FSWTJ7R
trJu51oLWTCIXZJgAR32cyDZaznzPaxcUB5DZmvvMZzS5xV3RY+1Dv7BIodDwSq+CIYef+jvccl3
Sfkb9U5q9/bOkJO9LutsqNy8f3k8oQ7BWj8QUzVy4kYCi8dgIlGiQ9XjJAJ1Otvs2UOol5Ik3Fil
JOxPdFBbVfWRYmQeWTJwWZXRRdjUhkuyYN8AQs3n8xTXbQ9fZEgnA7Gn8i2vg0mZogzPDhG2KrZr
AgIYdcwF13S0RjnfWss94H+VK2xG7c2LxG7LGjcw9BGubM0yhXQO54RrcFvfAe4+B+vT/GZ7mQsa
Qp/1DsivG+1CM8DnJAXaQhjaUhTKWoRwOAoL5Ymx00g8etKdE4DQj48ZwChfMPHaebydaSHG+iIy
Duo1WrSHvHKCePkvLCQcdKVlBotS1l6tCeO3j0Q/Fz1vAyHYj8Vww2B9DNeTwUvZEWHVXNCRElQd
FvDm5iC/3422zFmkWeyuDTkXyZHlpORsMb4C9wYA+uiJa1lG2O0fOgy1b4RmEL0Ppsd12BQuX7gY
SuxY0lxbjnPa5FhnzXlrMi4Y5Bdfyxv60Mjh9KzkX9rqc6nJQqt35c3WwwjU+RChPaZzzcDoYAO3
sB4o8ldVD4HxHwPu896kaSNTm2NAa6nPqoy/92hV0fR9au6V5GdX7K+glVbmI4US+tJD9c+TdUs1
srDB9pGumVP3W1dS0JXeGBUwsKre5c7i+FyVMJwot7ZGKp2xGuxW29rpqcEFeLCisqFif6ugkOl8
puhbQE0WegsEKAyNiNmTxKv1jGBjsYLbeYLFVj3j0m00BOwakiVmUW9P+3tMHJlMje0df9c+WAXH
PLcYnsHXrrYy/kj4yzqu05k/uqzqygVLwkf4/ZUi5Fn3zQKK5mOULhb+AhirN9yHg8O6NjJfe1PJ
YlGJZ40QFcyrHSTpJgcUeztNyNluhpSQmLFBBb08gvD9Xfl2ALTxKNk87bPNRuWfnUwN0XQf9Rfb
cJrXCjqAKEsTK/laElkPYu88T6cQPrAYyxtVU6A7X34O5QyMtKYmLxUR2ICYq8mdp/3jLQry11ee
nbTbDwwu8/nw7SdPxU+mcNc7GoISH/lD0ISQIRoj395RdNiDfe2VLqZUOSetWHMANBanJAui5VB0
7JU0Cicc6vV+bMApUfNBUL6IIpU8J3v5/IDnssoRbyHkNdsVFMhKd4YZGQmmjAwkcxeRl4IdPCUW
ZIPAbYu521jfNYrQCxGOMl8061d7jKh5kYAKyW6r0KYSD+X774jYfAoZVBo+GcoIerZiAFv7mlfm
x7LTx2juvd3cbGsBR3WYsnxNZ64b1pvAjcdyhENTC4V2b3Hae9LQwWfutibQD45fZDzGy9gBYu+J
4HeBQfHFVUPQG3G/U4EAoEoR+3MoWJlc9TQwCE9owJO6AgRf/EyFJLXQ9B9WO8+eeE8VrExXgJoz
91NS3I4LCwZ+g8GkISNrMREB9X8LWMBy7nReiCMICcCW+yze8QzutQ/flWS5B+zYPuNeXoNf+2tk
2dOgPpaYH6HzfQ/70xzdKEpQt7Ar76XNHawG/TQHnkRLKAavMmUdG6dpuoxwwhDa8e5rlz//xfks
u7hUwCJQR/w+97M7L2XsteWIxBd46WDSIwWn5ERuGmUyvSjLoJqgE9zzdbEv6wdh1qP5DpA5tAkX
J1d0RlVx6mU5AcUyc3D/rDZDvZMA6YyvW5OXyPlJwIU2YQoQPghXlieyzaND6RoB5EDJvlEZaJf5
Cf90P3rjmaJXSecYJCYbgPUn5ek2qqe3nEQpxtjdfydOtpb4wzmLxcy9p7HgO4PsO5dRnX8ob4tZ
du6PIJ4L24RJW7c3ZCrJp+C1FioknDPsh8w94cROCVXzGCmI2/oFy7Lw6FTGAFyQPljM3i70mWkF
jpFx5Hdzuoghi0hGfsbVThQ7Ok5epjI0k7wU1A+Rb+5DblvJlzK7OKDA8KCI0yOMRV4o4So8Etuz
L6miNzZR8fGiORrAJ5LCIaqIwfSTfeVXF6xMKsDWgt9vX8isckHhjaUQ1ReyGkF9RfW+TCZWTZ4F
dFzGXISotpPMWjAe4bpLHPL+/WeVO6TnTdEO5Dp/ouGHFF0rovWTs9NFRXEY8pJCaJ+0ZwDSzUT/
5JTzw0wsmeyr0vELz4k8ynQoEMBKG8kCRWuPnWTiyvmKjtuaBt08IrAVKP9IOXcG7nTB+sytqf6e
gXjb0mB2BN1uSqTVjdMovi2ecROe6F6L/7TKwV6c2P+r2ZhSnckXpQ8FwsQuNBzBtt/MMnqTHDU+
wlnOXXa3VJqtZ+6nAs9k2sRnJWzTA9y6qw7Culh4EDmhFm92dRzNBCwB2Zbo25KL5dXXQaGvEDsq
MS1HkgtDuQR8S0JLKDl42HMQmHD5iT8EbwxDV3LzWm3/3S2pxnWllfo65PZWst8LqBVxM0zchNvP
9YK/mQ8oazAKbii1cKMdeIR/Woc2vSYhK1+goWbuVuBc+1eVEAdSHZ3b1CiNXLqXxlUNJeV4oAs/
x4LooQ4ChIi3K5y+KSBg9C6gxU9ZRDN3aCZsBGXpLVY2/CqSif84JMR34WPKBCILHlgINiIs7Fd3
PE0sow/keryzaznS7gslpGdUXEE0TsBKdrV2xybozGWnkjG+YMSmsz6tp5c4wABggm7/mukGJukR
kafankdeMvj4ag9AXHoZfX0vg1SKNeiyTispPdgOGsCxGRzNJzfXHD2ldi8mtTdlPkWrSP4NC33c
CZ7SS+gFoPICtnnfs1TBjSjfic8MthT3q/3TGBAERN7FW4YP2SsMaUq9S0SX4zXBMdH0uVOMc6n5
GOpuBw2+wApX+YspJqEAfb+tLbo56202fo/uk5v3mFwJ8A9mSAHPLyC/7hc7WqdIhKvDkmVsk0xZ
Ca46GKf1KHd2jVc3ipsqoBTpsuXVzpHm2hVsjhoswX37V39uAxOthLKSkG1GRc/jlTBACtpqRLXL
ANbXCI3nWDHDA2nABE0NItgoXLi3JKkTY++e8Q/RZfJM8ZOZCxlJBtNPMW62KtwYOKy3zsYdtric
UgLHjR6uculmYVFwe/5IH5etVqHac7BzzJQA2n9Ak16OHWRrEz8u5MXlxpJf3TcfgZL3zVZvvg7V
aa+Jq0PCJqGIAsAsYKJNovUn55TlS7gvn98TttjvarLurIdd0h62pZsQhz51Un1B0LagNuTbuWdi
H08zuRVOBgxDZuj13Nec8qzkOctZCZ7wB++RynL0tGbPKVuspY8Y/YkR9TJeSZpKHOrAFmZWq0j7
UN1Ke5qyem/SDXYbYQ15vJ31i7lbKtLBmRM2ifzHr+e0jtsNutv9OcmSTDHO+xR0YhfSxB4zDWuA
DlifTf/RVCurwJf5NpvD16ypVsvpFzQl6TTMqHFCKhqXA7O1IWG2gZSvV1IdE0smjrvE6ZHKlT5z
PM6JBOr3g78q/S95iYpeo3iMsn4/CnVk8i7wZc6fAyg14CpY+uQjN8PBSDTjD9WNGNyK4vc5MXEe
SqOIIYc22mXrxmd05LMyfs+PkaXtDrOTOIMfbFTKFlqlU9jZlgSvK13bfmiTzzJME/SRl9Mg+Tqo
oCC7+Qjj1vNw7p/MkOv2vUHNBFHLcbc5qsBZktp2GjLvdJ/0rBhv+4rBfWsbBKBHYeISyDy4CeC1
LGud8eoX2YsZ4Pl1zBfzlCYiZIxyd/ELFosVX0imD5KXY73eEMrf8jmop5zP9Oq0WoeOvrxXV+Ke
iao4QAIpXcseyHAdgUY8nj3kWY6C3qWGE/aj5jk1xreiDQBrC+8zLQGrAbYJRB8AwyTZobW1D06J
X3QHz8vXG6kZNtakVkCjBLymin4OL9POTM6cJTiUtGyA41/+KB8tqoGaFhDby/l8JtL6/Ktjzsp/
oHxCll0QZY902tVT37bnnC0wXEd4976ASHobKSthAYPn4UbRa1Wcf2xBW5V85hFekB9JFW9hkrKZ
QMW4Ap+6D6yDKme2h+kxrDzD3MxWF3WmbTpcOJDEjY6Xgi7ypD77Vhbnu8UhasaY9e/2TjOJQl7k
Ck6BxPuZ7qSqEy/XzPJXNOpQ0IZAB1Kpfa2Wunh0crCULnnX1L0jBc38IMmiuPI54L6LQkMmtYWs
l6fnTNshO3l2vmhjgPSDrFen8cYgmEkR3raAR8sLoc8Joj9rzcVBset76J8lrzbrt6w8eBXmFRPP
mMgTrmJkmT8yQF1nPI4CwWZzrWdvtK6fcfyR00iPCHuxFuwJIHRN0IPVUxqY9fO0cc5Ad8LZto1l
uACiPQKHOpWdeWWkRCdZBgM72270k9FI2ahMAXC72iErycujBLEBlQRNmuZyPpfQ0Ut2U+o4+zIx
uz/i8RdB5yfm8/Be2nLFzQpWlguYHWrMdqOykQLepSRdyCQUEU0Llhdc4hdIRIw3BNaCQnEyRM/n
0rpUnhStKLY/hk7b3jskp9eTwKTxprJoMwPCGVzvz2LT3jtJLRWp/GV4csrItTbGhC74WGI4No4g
YMu1u6YXObuQyxkDawifvhvGaSL3snT4Sy7xkfNp1HwOr/beeQbptS44S26WtGNdyqiHyt86hUCp
Nd3frrBWUbFSHl4l3QYnzT0ll5qyuAc42Basrft+CtFgGybTalVqExsGmp5UsrvOZ1B+lRINXnqf
Ng7u3maZ8H/lFK8/O3Bw54pVTNUbCmBxe+ik0CaYbbu2bScSUfPAx+OK4nsdpndRLLqqsBkVvPds
Vqd6v0BmO84FwtmY9naKrwXbXLralwAa7vrxy+fAev4t5PxDN6Kqqz/oBcMqUx8jo8QIL+NV5aeI
Gf952GaqlFRhJh6j+6E7lQedI0ngOOqm3ULg2zw6qEwjfa+LmGHZ/nVIIiKaEYRRX1f5uOHuSxEM
KMPvrnvg9jfHqvyZBuzwnarYFUaibiC14Jf1BUrGb/QbLKkViAgs/n9PBjRaSSXQ7FutOFPG37gy
b24xuPq3u9YGd08NG9vl7P0k9LLT5l56GF6L3krtF+FdL8Jnjs/gVNgPsHyqE+CdJIW0FvoxoMaI
uDg+ZQ39XDPjBwPF5YyXwCEqaia1HUzAnqKVz3hnR/BVcj7cBSNkbtxAdRtCaSYoLqT+YDPCfxah
hirXMe1/NmggfoMRw8yqsxyPi088nuRyYwzbJ3t8IZFUvkhBy6e13yIvpoAPyW+MBqw4hzVh6XU7
HS/fMvyqfnL/skL9UWueJdzYirrRhhAQ/4VAUzgT7ewj6EI2WZBgWUcnOpGv6uL34yKcaZLLsYqO
Ch5e4Ta1DmXfcRiNDND3lXZRYcYVAuHyKafwh2tT5efYG88SWr3NwuxesraAebudxE+Qqe8LF0RZ
Vdc+LW3oyOaVoqkYoi8ZCE94eoQfycgZGUemw+aqDItFruO6Nf8W8o+oi9YdtYcLfy+RUKP35LKs
frl3j0rAuPB2QzMCTdpd/XUqYpP6Lhbh9yu7oaa0K7s9Mb68E3sb8sloqaB3fmYBLisP9UWOhc9G
Fj3b0gLmZUybFZLe2ZAALzV3kRpYpT7lKA7D3fKPXJqhI2WkRZUm3O3PkL7T9GelTb6IdmY5COIU
s77MzhLkFEmczBONVy9tVUiRXVjLzz+YOOwzkfKjnHRRivhmQcxjDeeVt0qMI8bihRHQ+9gsx+H2
CDIdAabSeXyq905RqiUkJmtkOoyuvH+snSzrePg1RsdpnwClTh1jk3NGI4G6GrL5BTgsCzjVOBb0
vFeEaf4HEcTwjJbO2YLS6AMdx3QkNWisaw01jCVE13E7FcxXj828qWNK4hnat9z/GYp5hyt/nFgT
BWgxn4borAnCUvViJYO/orbTKY3Qb3R8jZvxZbU7ljvjlLy/XYnZ7ylyDmVj2C93GRDOll59rShx
+P0MANxGScjq/eOSM/IpYVebV/qdcwWglnFcclNSteipWHmaeU1aVaqZwVSatVp3yeXLEP3REXlx
2Oxb5EO6bB5YO2VjAoSTNua169GyzlHk13Bx6q18ULNafGaMpEUm9yCidZ+onZPDtfRTARCoP4yV
SXYD3KvJjR2K8WO1TZwlEqP0LVvzxBrNSRkDpW1SsoraML1yoEuKcMdJIx55rO49Eih5ovGD62Sf
K92StxZwQJwU4UFdp847GUYAajnmcGGwOmoLvYY7KvtV1wkwbElgGNIlWL+PvEv9ZBS//JF7D//P
/sm5g9q7HYntxWK5OJRHJC5RRr28JiQHJMY+xEd+c8vk0YPM/7e/sU1OPJqqCyXSsQh0jflEUP+l
qDX+vMwy6brMySnPNSEBZ9GCOw+L8zqbc0O+u+dstF2jNClNChvs3fJcJnBfhEEOFkam4Y0l9RIh
i2suDhqYkDH+2KycjAnU45hOGxe0tGU8AtAV1WjgxklEfEbpvCSCZiIKPwTRBGNOtcTkZQvDLmxM
zpxBmpjdXF3gAgIfXKB5xRVzE4jS7vgN8ovI6+GjChdcMONXVXtqREXBSs+lI7DuSPWsMjC5cTgv
VRzcjuAhO6T+0OZ086fXhAgPBm2XQgFyBhrzvHjekiKaVEJFe/FzD2JrjRm019cZvWey4NrwUdhD
E+3sU1mBvaccAySoc5BUfoRdv81TBgRFdPfBDCzqSWSsgLMnMwtmGXLH465gpp91h/tJphJ+gui9
BxShIfyE50umHDMXxBwMtUsyJSkjfUD3U3zPJskh2xBJf2MIpxfYnrhQ4vdl4fxYJDjDBDZimvoF
qgAmF/C3UgNvFEzTN/qNa4WEt1Z2bVtWRKj6IEibdnStrXXFAXGRUR21q30S2g+m1gNkCNhR0sQb
FE44bT4axa6ddwB7DNqbMX0u/KVn1w8bOHERYhoeqUM2+NUuNT7xDPHtll5BqLMtJtPajJseXaa6
vBdSeSjvRs7Ti98Jm6wdwzg5S2A2xTzCJhQtX6ia3tm5qIEtmBVTiPio6dG9RM5NqgPhoBKAj5ag
GNun4HO8aSaTR7ZDArqYHHAXhAvn4Dgax8F64XPJxB1c1wgEkQ5qm9D1y21QHizw7QsSJoKLW9tE
TsOklVMctcbp+ejvMmTFL4BoZnzqjHqF0EJpP4aSTDWi/Y2L+743Pa7UX8wFLw5PtYPss95sDUgj
OSdhZFmXLXTZEDfwvmpFfIVxbf3WiKs0E+VoF9EUlqjElZ7XlDrgWx3Y/vw44bUBl116UU732CBY
e5ncZlg592dPPe0w/c8uld6IkCnKQjsMy8IqsiMxhGFlVOpg+HtW7WFc81b3fqn43PJGBlzSlgL7
GY/A1ZnEgvLt8elrcwcbFlYMjaTZpzZsfoDElwloMDQsx/UwBZQCKSWZzDAX+vJYGNWe1nseIXw6
vKmpAuIPYOXprGHwSiuvdzsatvbdNcwmVadM5MgCmw+vxKtCfXPJqxzb5OGtHmQrY7kKXwhYqmee
JjIf+TCtapiCWB/Ss+V6KnEbgoFkhzzO9XIAMSbbcwrZCtRhEwggS3UDeVXjvCA9OEsjkR1Ce/DK
jLViiRmO2oEhATOCs1qVQMo0I0S8Ot9mquJBapO6/pBH20na7WRz8IWklxWgTSEM8aEacn1FYI3g
UVPu1yEEe0awBQ6XdGciIeZXWU70d1LVsZCLJKDgqI0xt1ljteHrbwdLQyfDWp9otzYXY9QmbGDO
4qkmv7K0FvzFIsdlvF0Ep12BVRmyVLzp5/6eHpwLy0iCf670ei3ompLr8G74IPJirWW7B3YTkwZV
1dFBw09b33bkByvV69ZDuqlTigEB/zosvMPnTnvMgwBGqB7D8im8JzQQL/5WA+uIzD5rY3on5ZLS
jIUcDfNPE2XZ8Aumwg1+AUV7B2ap6hqR/OyUmH1J1hHI+4zXq898FOYtkv3toB6atW5mRWxaJCbd
CecLSmuaei0o8rrcRG2sPLSZD2Ebmi9cg97gCbzwkS1OEb8PAPTmZ7TIgsnvrsz/WdsqXeflc04t
iz2679PMLZbVpri0T92p6eKRVwrNsRiH7EhE3Nfjiu0Vie/jFnrzNBaWqXnmAXAmGS5yKkP/vHYb
tt/ITsboLlUtf1EbxKq+NONQ2P37CBc2xqq1a6cFSVS+e64+UggeMCj17n9UbbSYv+aJ/UfdqaCD
1mOJ6V0J6bO8pSq0znAgeFQW21eBO2lUpuGQ8aOi3Fd03e0AlgYjLD9NxC8yEqCkPJVowVXwl4RO
cWzf6xYV0cdCapSL3v7k7xCRQcfST1bWiolnsHsIG4lkv8pSae4vA8HEL2agAWAdy2vkDLW82rCm
zb65tAoho1877Is6KfkPW99h43Gdz3qak40bjrdSPOiRWi6MXQNuvQi/FRKxXOtQJQ1K1rfTXAWs
yRlV2wzgy4eSjOvTWDnExkxu+qPoiKjA1UYepvY/Q4GfYRqmLC4INrut5rss2q6PkkvgV6NgxksI
tsptPBMgreUaaQlPWdZMBZ53PHz9eImPZFku1+gZOqTe2m1sTaoeWiahPzk71ycnToTRwNs9yQdp
5WbdycKcDhp0+MSt29HlQeSNE5V1xFDbqO2puJxBlHeRIyR0V22Ej/yifVcrjVmVpakBC0OStY9w
KiN85rJx8rWhSr6YGYf5m6CQr5jVHAIutYV/ny/DrBtlVqFmo7hr1Qpy7OpF0Vp3x554BiuDedF7
LBQMDS8sHBj5okj2SQeduMAWYJ6rjiuRUqhNYnFUlnmbR9tkwf8fq+is3jYsfUlohIugkgq5oE3L
/+zCyMiEkiOYJzdGEowgC8P1MdUm+HgjEPXh7buJGzU1ScrGXkrAlrAlI+JV2SCMtpJH3o/U7/H/
Iv+FnsonCTwNufUkC3OJV2CRC/qmnMRIbGCZb0CzwBrtmmvN7VMar8nWZwSrvneynaNso6YyEQ/n
zN/2qgmTOQFK/Vr8EoOjSRV7i//RIWBu8Li+bO/JGd+cIMhmDlFV3AqbAhniZFHuyeIsxfA0XxQQ
wbMrJmVq4RwBmAEYLIFzf22F7Gr9uydFxq24AIMaHyKgW7CFIW6Yf2HfU+D0KymnvqroU2MGB92u
ZuyzxTKp/xNDXd3mGdp9PHBg/IRKrl8A2XTgzRlia8k+/iG1I78lIgRN+SGEopYIrfUf79HXCSDP
krME3mGJNpQzalnglkYBu+H+WMEJdY3mNOY/kPpZ3QUd5uhNE5wRgqCV6yR0ROPjgpR7kbZCVRvL
FwMGinmw/ptbJpDOuFplqG8fNj31BAQn/2YmjgT0OFNxYJ4QwbF2SmJqJoCVVJqIHtj0EKe6DqM1
1SCWEe0ItvqulNwR3dixu/H6KTrKFa2P4f39624IYJf1b02qBbB41xuBTWb+b+ARn7N9lPDPz/G5
SG+K/WN9NUVsJSjmX3HSHtA0k6ynG4UdjpeDiVuA5fMhxtSaxXnT8TkfSgl/+7ivdPGE5qxKff2z
5G8LXa7XabFxOLkLFGZHssjfhI1ty++zsuuYKicFOLfnwKxET+Avui5lcYrcL/ne96L4+DpsY/1t
a5ssXMcpqEXNnoqk+oiPI4gcXGSJLCVSla7jKCQuun+j3LwQM1bLzC9TEEj5vAwosv+Ie0Q1FuFE
4l9RGya30hyEq2DNKIwLE2Uz5CsvaN+NeSq0RP97aNyPVe1hwu3dq2p4xRCbWSl1FbRhvo5iSC8e
cxMwhsU+27dnFxGQVgMu1uB0SfWfhmnNUQGs9FAW4/hxitsXJFJ3d+61dn5zopbyz3MKj2YzGKQQ
b9+spnzKoWgtujUNixcoJd/QjpNIQpEXiLc1C9sGvF5eqsMyGAH6mIZEZvSyu+QkZAl7727ILyuq
IovyjGqmlcjhEVGg6Y8eIzai3TsdHZWG/6iXZpb3FiseI/lroBR40WoMqKdzDUKCVshZTRmJpqyK
D9JRaYk2eW3HxnIKFVzxcB4kp2HyybHzhkDXG/N1UQtS83SOoJpA5DvM2tdVuIdNUHMzYkWP78l8
R/gTx41G49czsDQEJ8KmT7t8E9UAuSTucvdqazHjRKhW0uq0ml7fCEaluFY8dYgYaqNGUZ5CkeoL
2grv3OIeVOAbKomEM5Q4w4Mxa9haQREb8Kl0vwnZY1oEEG3Pn+y39Pj84AobdN2o8r9VTHuV5xd5
lN2uTIPjyCYbXTOj7x/5+43zzkGrHL8naVTBDKpuiFTDNP7268/OUtMxK1pGINryl6djBbLmJoJW
y5HK0He7vxCzNwwXGkGRCr6qJZKF6O9juCFmVjoH3gLRoNRw+8TpxXMKLsm01/b/wpSYbv6hJPoL
8fpGeauKIHVdgoNI2ogYMbbp+bX2/jSBohdGVrKOAnIJysDUX0sNnPZ5nG75fkRPkNT4XmRpCx+X
9esLvQinuiLfHCOWH63KPqNFfRTp2mubEPvASvUo5ZKNfRzcWXcrim+KnpdKqJ8MRme+Db9ccglx
Eb2Q3xqP7LMFz3nXf79cZgQ6W2VKFTHLUlc1Qlc+aKQrzpotUugzqkddiYhfz3OD8cR1BPgHwqqQ
J8chw+QBt7JaEESq3VaKZtC1fasTxL+zs/Qmq9fHayQC4Nc0p9zgCfEVoRB2kDddnH/05J7f4Wqj
9aCM31HYNzy55V3RiSffUJy248oDWX1s1zXcOMxHOPMnqZcRJqiD7MM8i0hzE95fEqWjikWctD1X
wVaMnals/dNc5e8GZ2WQtSCpf4+1g0F3tqEsLg9qj27wUWOjDbySyAVChMNU2jF5F7/3oaSoEYCj
ts/t8KJBU8A6jstugpcIJPtIqaVtQw75N73s6sUuiHt8wIhxQ8hNpkjffeClYc4WR20vgSUWf34l
CgPj3EqrYnOe+YVUZg1kyISS1NKnDdDuuk5BhpPENxrNnDk9nNYokUxCTHK93vnBDiCFY+TdoJBC
MRjW4ctU3HCdl6F94PAX1dzjhN+DshGIBzMFN9LR/YgfOIzR+eDJSxBqLRAv8YDiaf4C4/zyYEPU
u/CKEvVW2MHey1+ffTbz5ziaUxBCUAYpskvo+1sVyAl15M8AKn+RdJhYbNoAGCkFgiLW0IJcwliZ
w6P9vHe3MPGoVMliHmN6psfqldry75cqN8An9GKCx52b6tOSaKragsoecldVv+9tZCMxUNCxx/PS
arCPGHu8R0z4F1MwQEWjAbHKveo/J0owRrVESA5f//td1sT1tuQeliyzvTkR1W0WOXY2g+/H/SOX
cNz5bDy3K1gyNAnfnOmv49dAH5ZBqyffUlTMAI38SNIg3j5ztTegInuJZl37LTiKi7/A2ss0Nl41
7o/ckcw4hkgoaeMb0J3Xh+r+SqpjXwo1avyCm024sO5e3AahGmwHkWSkcrhRQp7ajFqEB2zPlIEz
0q76WY8FmSaL8VJZ0UhyYdszhIjlqH221clL9MjrlB3mZr/ylqqG0+wkANaNgJicaMueyIn1TSD8
KdlyjYLZqyPfXEek0Jcaxy7fk/uzrD+y/OKTXLnYNA1Nf0jLBp+eJ+FZ5AWd/hlsONt6HcloHKTM
f5FBzWrGKvtJu9f0k6tZWCo0BLXFvnd/xXWphtJEWpWWskpK4P/3jtRO8wTLKf2n+wq7mgDx+8Qz
gbKRMxRmzhiVgepOTy0k5DPs1smBdhob4N1PmWdAf+OvLRndl9IzM3cxcvmrixbkQW+OekP4Ijzo
C/ugTuvkFT3PR+SsGCmmX4B1ECfGpZpz1RHWxn2lFZBBAPYSqHB5DuaIwadwxKcrGLz8J9gs3Fl9
1wc7pWZAI91ll6QmHw25dJ6Tf0pRz8bzlwHoZ9+2ZMt1urweMs2ZVb6qE2oB5MLHmlYWkabuHZ/c
KMRXncLFDMQuBciauDc9CvbwPvHOpo9MgDHkRI2qbUv1MGdpWLp2ryZzOzI/9P0tM72H8hxj4CDt
RZoLfBhKxvBu71eKCV2wqyPK3eSuANaHRHrKsHqQ0rk9XBSaaJz/ja/0Z2CAU/qkTkN7eb7l9hEN
nrgJfuy/RScw9BOAmyZGH0LaEfIUUl4Knj/aBPDfs26yqAnDZ+kyzV3DUPyS33zTHtjxuzwsZaKg
XxZSmQbJM9SaWE3AXGZo5IFhXw3r5xkKOSbmyhGqjerMQDDWDB0dN/MPqJmckXpM14IOOH5GaZiW
+yQFAi5xS3ZqmLOXquOAGO5fwKVtyyyzJwKePk53EenLpeOLNAg9SOvU5CeZarhxmTornWgTYl2Y
Ob8f0EEXCu3CK3tk5fEp9XcVLg6hSA0t0btNByeDBMhUwAfbVwql2M29J7UAOekA6LtxXBpKw3rC
bTSykLd47z4sc0vGvPjEIlgl74blw7oUB6L7BkENeMjj1+S6XsYQ6e2XNY5CBHm9UeBtwwp+ITJB
RfLDhBJwvSi1jTQBKtMw52JhGwdeRgHTsLk7ItoY9tZSx6U0Emunqd5AzhsBCWQqbfaFbIKR4DbW
yn0/LP8jab7Y70NsIklCCl9x4TD/GaadXGqvspPYe7GAMD3dmoulikTERKQwq9ffVNoVHTQ62+fB
/XtHRYpZ9FG0mb+sw0sW2MwpxSr9PcXDkbx8r0WwcYXoh7GLMummFzHONsyfJwuykv8y8NXMkpZ2
2wqfb7qutvez6JhIEStNiO+rGXE/aitXP75QqtGmvalkwlXCnS7FuCxr+dcM2zW+HbZac3atgK8L
/vDTSkZD9ybKp7+OS2MoujGvJr/Ge2E0h/MoBHMyBQ3/CYR/TrxlS16qZ3qTludZlp6QuWBNA/nq
CCWBcyM20FM9mJq5O8+azWBK0NoRKIt7wW032w0MjuCiPO08Gsgp35o8uoPAns+UOLKPbygSs4RE
AKwhZcW8V+9YDJVKBxZ0Pwd976ASGG6ZPaXhfR8JlI3NK7BGAHykHRU2J7q/LDs6nhO5l07OJBO2
538j8FJlu7PSw3tVKfY6/qAqETxQCGa3PZLBk/INUAwOey9BJZi+s8S7DLUjeXTmhT2E99mzPZMs
7P0uzGK2f+/I0pdfSwnD8NW0zwGkPUNgvbQaUcJm4jk23RzEfFjl7ICt4bLHqU+LIsNg4GJkRpfD
4HSl9Sp4JhJvJyal4kukkRohJOjkxreJYgCa0eN1uBZZgiNf1ijdYKyxWsXTmCWlrxyDAS9GBjvF
w5r3yGgEMh0BbDYFU/Ckn7b8VLxcoPj6dz0U/r6n1KZPDCw3hiq18yl/2DiFrzuIaKX3VgV8IChB
6p7V3RlVDh0wxgaXdCJn59UdZoNG88pNewqIwfVmCdusu8mlbvc1XzF9+wdM1E1jD/5YRMsAYUj5
Voa8J7XPnZVt2rL6b37szvf5wHO5tEMAP1TussCmRHcQy7BJDH93HQxxhJd+TIbYBsDPo1ofogNu
tt9XL7sxzBcPKZp/WQUvzkIBoNfOKudP5udleFTCpbaNEgVbn798wE4THgFe2Vi64eiCRVaumZTW
9oQdR7xGFHoxZvwOcJFhjWhspngGKncNbhMfG8YLRryWLczBcooEnmMFpzPBsmyzYfiSUwQtvn9a
BN+k1Oa1YgqLEf95rKiG25E7bKbnCzXVkj1D4tDf3KK80KdNu83mMgAkzXY44iHWilz+lefBCxG9
3oARzBpKqqKjmxox4wuZtCTaD32TUBQ896DNgOwYp/VzegtfVVZ4nDR5rKZ2iLXpyGdZWJ6dB+j6
mr+RfwLNyvd1O2Y6uPr2V/wNjFBPbGFqYQYCwjmh4q6T37ecILSLOHp3+WoU/e9S/GYbxq1BYGoB
FPWTswA9MTwlfULv/E63x7E5K9MAUsTmDXUkEYBAim6NJ6mpXx2tHmq41RONfBOsryZdUIKeqyxc
0RSvkhSYzzoybeRksI75AhwPeyboTPCzvcUBkSDFoumuN4xhLCopOHaCc3oF8v8CuJEY9SO95oKU
hNz3VwIAtaWGLUyqoPBXLn3yLhTafEcWgMMWyEqA+12mHpC6WaUkQTURBqz/lPJwIlUoNbR7Meq4
OUfcgoDo3VaIsmU2wIbQ7edcqR0KXKs/uwM8QRIK4xG+RhAeebrr1HC3MKXBgOu7CC2uKJE/7tR+
119GIdTgm9Sh7AI8CXNxZt6uWliruYwtKQSutbXKHPkN/x/xBEbcx0BFGjYqTGIXp5CFQMxQixGk
rUsqZhl57hkWoEX70ONQRKZ6vwRo4tI44N278QiioeyANbU65UBt41K0pjxuYH51Fh0uCyhOJUqS
qaFLkFEAbBQCygRgYiHwWs5FNdZ6O44jt4i2+0h/X0KM9j02bvQ8Ig3bxto/9zBIY2D2w6m1kAAl
8UlGd23+CUua/6EjIszOQEdevrXT/g/jSuJ6Yjw8OSHMCMVUFtu8w3//inoFw7AVA4O5tf//XaIf
FH/lMjRI929Vlh0bEDEX8oogkZVso2V37f46eWOJBENo0NcVhPvYg7hczcfCioZ0RFLE3nEY88J5
pvHoPG3dHu/wOdJrnJ45nVwUUYKYGgjskG/G6b0DDeLTrjWjICYccyBAXz6IYkycyUJ8eH0VdUHE
VojRiSb+33BaDL3yGxC/+gaglA/7rxTuO5cd9fhVST4QP9ifrIL58DDGqO4oh8MUM6KcM4p5S3/H
FItu+NLUs2t4hse27OIQTdM2XlMQ4K0O7mseTWDB/QROoPUdzNI0wb1v4OsM3VlFNwvuoZY4W21i
UafdSQOjqJdtw3jkhD/pMumusR10Eyx06nLh112UP5OOc473vqAKWrFInYEV/dsJHpoGwilLW1bd
+eC75QGk8Kink0odgRk+ZXpPIVvlbSrjWqnXLjXjkheWPkiY1R/tZxLei5H3bOR01HX3otf7tG79
ltD4ZVmXrQQI6n9jkpKnY+d5TAAj28CtfBBLG69dzc3pVotyNbAzGva78lc3n+KQ8ZPfXq/fO9YI
+EF4ZtPkjIXgGJp89C3yznWgSn1C5VfTLLIGoENCwDrUZmFhs33rc1C6sy9pwUVO1ZXAVTA7z34M
3wxViK8cczLtGvM9qvbvr+R+uaRem0IaGwYruXZTBz6w8A3Z4wvXYGrzsOW7UFccw6BWSbMVPfVM
AiJOIlMwmX/YekMsvgnhnldIj0p2jhumxNTEt5VUKw/LMUebpbBx8XNTZSaeq7CYw0dTqJEGBTJv
IqNAVwRh43ziN+MDofFMRJ0iKrpyeWhuKv0Zijh7oU8yyhY0SKiIxXDpmbpwQfoRJHuA2Bv8vfjh
Vnqs4PLaETA14RpeYXc/TH6a8/AhgotB9kti2ZR5GuHoph69WcsYl1dNWOHxNN68pnhDqEtgIIbX
zvnzndhG4gyWlSOH/Wa4BKLRQcJbS9WoTGSBMrABZrYamATLOWSdNBLjFfmOJkRY2J/vkaNfqlEx
yKWGJOXF9SAWDQ5gpC2fBO+WcZJ/U2IEgRycnfLzrRaOtJutCrvQe3SyYDENTu8DRimVU8a8VUUZ
thSbxeDhtg57KKw0dbs4iSXAo1c58lqccqdVLtHrja4UogihH/NhT7SvsJT8fztDdWxjxnq9tJmW
B6D5eSopDy9wyRVuufRq0WiZsASFmr4pNoEnD5zi8xEjS1URLdIPeQ3z0/TRqpehVD/DIbTlnP70
5FwTxgiijFL+OMiZTGmpkEuac+Qbu1uIbGdKTVSm+tT495z+MDpUJ986CoXRd7P4GaHyM+XqK03H
sgzOwn/yEbpWWzzPvACndpLF3frljoPKv2medueiYm5/5miLyQzOCTaC9H8oRuloMgBU6fUvO7mA
eM2wXyMjTSQ+aa5su8PKMe1kaoRgtSuhsJTS7b9T8FxHiwh4Z1fYMtodSMQPae4x/JfFVEA18WIe
ERr63KhH8vx4kT9tTq2Jv6nefqqybU7FlieG2xSshGOkD1Dpcd/N3iyHziS8wkDFUoc7KhHzV4qx
bDAT3MBjcPNBW/kMfLBBsMVVuGIuK4W9cKAVHOXdPk7FC4oz5KEhEw2f3GAjgJN72AIqwkSRe5+z
o574LhXUtDwMrfnILfAnPF7Kw+962ooqCBsptUEKk8TG4/HdnJ0IQug1LHt34rYJiv32hngKkQDl
awgdGPR1MR+1EOQyc8qJAOy56FxYBj2HBZsXNXFtRqBFCf1gTVdCUALpa9Z2Zty8qWdAF5r5vII4
YaNhStSutyXyCU03aQXv49HGu0Id6Xf5vD3Dw/z56Ly03qV7Qp1K2f3WzFsoueUYF/v9YFuRWTzb
eP6BWTmL55AuOnu3/eCEk1qF4wYqLAFyLUPlAoocN3VWW0S8CRDcKT7CIz4RmmQ9KckhtiHiy7Xg
nIuWqqp7CTgfZudsvK2lvQsfQp7ckFw/vf2WTCdb9IHZSpkVEXsc/Q4+5uQ89x8IHWiWutkPMzSA
Ku8iSVL7v6tvyPNYe7jk6RVtxKOSfDd03w3rUS4cCCJjcn1mj9jYB07ZDKadOlYTUUBA3BO5daW/
02H3mBAZi+Cj9nN0c0dCVLyhP01i0xe8K2daoq1iUQlJBjNeadGm4901XNFiEsJ0gaiVkuSWax8x
aExOYHBQKSDBHoA4hE8y/qqulsvNGV3bx6+ZZnujex0F3600ri4/KTdw7QdwwkKtviKTza0TxC5d
1p/MSALSQRLy5LxnPwYziUQdAKFaVhPzN5fH2oDN2s07adzdC3v9RjpNIp252eRyuU8nqSnTJ3vs
Uo1iQxWcoglttWH1QOOUhTpapX6orWrZEF2q3hKIqN05pvoxIo9bottZuDKIEveI8lt/8Xl+LdI2
NKFyUDFE0mEPKvB+0ldD5aaWF/PeSJM518IuvtOlS9fuBOpl03syRUXciS2dg4mVVYfY7+Ixn/ta
Q9RQWuQW8oBZ1LAQqbYH9LfgIRq16C2SNZn0DCkzqRvuoNY+vsbtxubnFDXYK6+pEGWesUT5jpfH
iF97RnOgjq2Ed+FB6Bk6Enp9AgAdQJX+taCgAkdOcmNt0eI+i79CBu2Gy8jlCvIPFrd1LgffuFik
n7vSyV+QTUKzHNqUmfY+wfb9no7dqNT9UFnGi91uP3zz2GL+tgBckbLZ3oZb2IXs1RCLfE2EiQkK
8+NZgIekP5cLhlXyugs0yzKzoMRXMsob2Ak/TwT0u9I/ml3h8a+n8wkniCFKuWhNdt2iYsE/Qb+R
56GGzM7LIzth6bMX86BVuNLAMe0Qk9aierxzAe7k7qinEymG6tLeywXS0ihQgxM2XB/+GKeKbSIP
im7gkYscE1XakvgtCcr7Defsg6/0ElPrzdaf9DStolHIUs/23ZYVO596TM0eImmDs81Of5Ea1NqS
X1w9a0gmgFvGPI0eqX/jEW9d+az6t/e4xVSukGgK/2qrEcmrOy7blQrmi+Hw+NvEHzXY7QJiF/Da
sa3lA2crlH/nmYiw/RP8YE0C6l+A7Br27Fd7cMqWjSZZ4OnX9gcECKgFK6EA2V5WfK10vhgMLsxp
sW3zNQx4VaArIc1ysCkIx7dlq0Kvv58VIS7LNHQ75VoFtHHrxWIPMZnvxaJuXVmhM1iQ/INfSVQf
65C2rwndo2f9b9I+j+9BkUbAabY6lp2YioYnJu9e+S/L8uJ9mabAa99r+NPF/jdH3ZqVWL6d49vy
bXJig9COdm5wwDVfyOx0Xjc1WVX2TmoaFP/QIVfZ5J4C9oaUH9oRrx7aYNyqVtk27BCHZZFWd35l
XdeDNlE/zEwo6lUdEidGTOQRgIp+UOq7w/se81ZinYb5O5mhTOh4VMR5TywMra9sZiTQwESD72nE
t7wFTWlJdzdXaWWIC+Bilcd59gdItd97WUoU3Je6SK9LrfPcrm5nhkIsRG43AWHdAIaxvsDqK1VT
vqaPahni12x459cc+YFUHwxwEhNUwQ9OTJTm08B0CL8h9Tu937sYo/C0iQnBmm2iSalHuGUd99vf
gRZ1NJll+1cZkAJm1j3vyiyaw5kRUzyc/lJkDe+/fQhqs54Zf5D3EkWXyjuVbRrn6wfKZiX76OB8
Hr2DW6gj9Y/H935et3Tt7Syt9l3c5Sxr28Ulls+JcT1AGhH5q1yKF94gurqgszwPoDZSdoOrUCNK
0WZmBXyexBwHMiZRuQJx/PE0gj+L/v7zfycnsgErs89KpxUM7Z09YC9Eqq/LQj9dtyIVk61xpPZ9
CN0+U638E1Dq+UVGEMjlCeSmoa1GOEuNQ4sl6K0CTR/4fCOJtRqzhz6drQ+vsmClx63m2FI/JcJv
J3oyoLFEDEQcMctN3X4UCqZVD65hAX12fwo1uSEoRCnb3bpsdg10LkerwzR5itHzKVWBxkQ5m3u0
58wuRTwPWiyonsegGQ29RxoAoaorJX/djhRksS/DQuQ/SG5WKDBiypzVJrHu7xAYntAh7nV2o+2j
x6eMxpBPk+aJCDYcCTn8SbsBGnjwxly2JEo74DDKSRLKdlG0bGVLmoh+B/4cGt9RJNAVQgNXQV3x
yc7jp1iC7N+jXtI93WfyMXhNUyjVCwk9Orc2y9M1UsYep2nT/bKndc4en4gb9T43DJljIEV+8rNc
Wgg5HjgX56WviYRof6Y7IdECSAUZg0zQ974yrXHvCiJ8crkjvo2rWaB6anHyYx9wPvy/F47dSlES
AS5KIIWWczZNfbIiC+k98ce2l6o4F4yGM8bPU9VeplxdeHMJSlHJb+nAlqJFO6ZElYUJCfhojdfV
lj6rePzqMROuSNDMyRD45Plyx9+pGNwxofD+Z/XlTnG+7Jp4xzKup7rDgXZRewk/FtV3ApyFvwj0
jqhO/2iqsd+gcKUovVTLlA6EmOOAYJxmlxSuwhnyqWTPhDkN/YQEICO0VN+9uEES2cmCUmUlReqc
mxgoZigdEYENgI8xFhUBmmCIBovoI/wpZdgWkMWsXXGO5naYG7YNT/5CChr/9IohPfobGyD+YDmJ
NCTA0t7LjOvXoQJdGqgwCG8buXKHBBFGLhXybEGIepzCsTPuP5FWwHqoeY4jG958VGNDiXxC+ONh
6BM23JVpN0ZLjN0XDR75BMr+Z8u9RCB2VnAV1IyLoY2jGnBmcG2mYEkva0ASNTg3DCh0mgsLAr2x
5IG2nNyG78ZT8HBMdD4N4MXD3o3V3hQ8iwiLftuBFuzwB58slc2uYqJuOveb7bCL4nPd+bt1YEqp
axYzzNRstcGaXeq8b9r+FK5TIcTS+T3zkcmrXURhbB85HODWzKPd/M8wcMWp8ErahDJh3MqEfVOE
5L6QALMWr1eievXSr3y/qc3ZT3OaPXHnim1zDFCCknbMXfXMp70dz8TxotpBYl/a7otU/9zODypV
6O/Bi0rjRHLNXMu1bIMnF5KqncaYOagE77pJb7UKFjBawssyT+HIPbw46i9xdUFbnXn6x2rlunPW
4UFcLii6byW2bLcT8Jh7YjE1uaAY1/xrRqMLHpPDCkajmimM2YWjNeLywUTM+RXYxQiMQoHokxVR
q2GLlvLsHlVThsf+uJx+CQfAEHdEWyh4yk6Lrua7hR6P799DD8qhjdpvtCytMwP0B5j+8j8g6vMF
eHAfafG7x5Y+V1gN2r/YXmYZy+9wsk/+6mvezxF8esPRUenvz0kpyOjAZJWxfn1feOHV7H9YY/ox
b8CArqYQ7PGV/xEzzB+3nNmEKqPOf6nOZiWcLClfXW/VRXgXkeWCb6kw5Wc1weAWwSyg3/Qa6x/B
bpb8lfPrTICtAS63MGAWUPdtLR4vyQ4WakxP8gJT5Cs3zqnnRkgqKjlg0tYPlGmVJKUbRKekpB8V
u17TSIPfQnzt9jEN+XZoXJ2N2e62xRFAdcjDw3XgOX18+Rvb3+8f24AKGjlroPtHCFwpaUFDFKWq
6G5jgJywLu2/aDLE/g/GiByJDkh+Zlz7r2aG2W1ygkPGsjDxEVwjl0GjblqJRkNDB6zxMKzSDH7E
t3/iq9jM2mbAelki40yGpmFDU6GhUJ7LBMtjMCWOWhZbP2W6Uawthn/ffKPNI/0Plhnz7G4KdZez
SXbiiLoK45jB3bldkOdxqa8ADW50CpZ3B/6EQomTduHWNPy2ONn+DIbXMhvw/WzH3ivbQYKzm+k3
skj4dhtaSkw0+ooQebOM9aIt6P9p4iHQVvYzl8I+jll/wW1VxtZZH1IVf9aMnhD/OCdpK/hlLGKy
nYz86U/v0lc4lNjGFqMzabPH41D24o3dc1+Hr88xpnn8e29ZwO7QctXQLRWmwSoePVanHzRzN3pm
K6kjU/1iSSbjzkaqZnCb0r+lS5oByxsPbA6QPkSBOLMmfWkmgDCfUdFvJi83FO3J3ss6n8VOM6bN
XEXJ3ha+PY/RvFwWzPf7cfD4TcvCGZHhcP25HfEupg1H9rdVfJE4PwEz1thpe4UCFQUw9xAUIIr4
As7Ad+oY2QV0VMKqkL0ZEo88EfC6Xy+SHeBAElrKPaV6qwCdKWI2nZuD0Ugx+H1xZxlJSvt0+64n
tWqyWd5/RwN2/8uoU4aY5qhohVPPW6D6kz2q2YLCFjUQM96xcHgFJtEx2Wpd1UW/ihuh1QZZBXPp
vMNPfyV3Klh3/PWBdeIj8hmGwDt2W5t1Wn3AJjowpH4B/qWIo/mBRutXAtowJ0sn9eNlB4HVJSI1
Lf/1OddehwuyOjtWVgjg2DNJyngHuuPXzsTXOrv+mRKXfGS80rYJysVKRxQLhpbXUy+0fknRKmLE
cVCRxAYl9uWr1T3BpYffPdULGnHZEOF63rz0wuD9lnIzmbKBhPxL++vXjeq4Q69Rn9OKg9W3Ggh/
xCteX11dDKgMqLEYBLKXWruPP1h2waRfH5k64Cr0Gipk6BA6Zn2TG1BwKHshFVKPQRm9Go1H+z8V
r4llqeu+ElNUT6Zc2Khm8fscaaKNAQA0vlCbs5OFFbwejOzBX6fr2eGZZRw8Hul8T6NExNc+DzeR
eMhSCml9x1eQXvlvjpEqc6iFSJ28ZLhtguR3XK5+D9IwgLBZqC6NQU5/p5RKn78HC3Z70YMi2uKi
IZCuE85wHv8OSbQ+hnR3zm7YqnfVZmiYwuhtVvl7YBQHf2SoGe/CRED4i8F18CE41wWXvxLIZ/io
hEACXpplNbFyQmgmldMQug9h7NLGpa8njbq7Z74coHKW5IL1RYCVXO60kqp694m4gW8maNg9Ww6z
MEZGxVJ48MN7xi8o0XovgmQjfeOECLJ3/fi/NugtaT5Zm2PgAe2iCUNZj2kdq0yADYy98DPkveFl
/oyqB3pQqzNc9bZK8lzD76DmxCBIJtrkZHYqb3gKAlCQeIsM66MWaVePKGtN1zY4Mg1xpa1SGCB/
LDpdqw2koaD9NurTGGlz6v0PU/5IVX4YtreFNtC31ZYWWGdi4y5aIfY0EDYAZv+9IHBqGvPTC0Ip
tlJQFHX0TeLcx3+goINEcL5z1Zb2OmviVoEimSnjM+NzHYkLEoj8LFU6LDrp3fSTzq9LGq32GQSS
gEMmsQvfg1SiMbPEwz5xMOa9UtpVAnsJGFraCXcM0emKlzS9GDXDjbb18OOmJe0LAFuUX+TSlUR0
A/seI+/tTiHf9r0S+MyZQmGumnJVWQQbQ9NFQNv9KbBl4YthEBzzEFLnwZDdM7jxqz6h9WU15TNL
sEPkoh4sJbsesJOpmvAn7SqFOTge//hZ6ZvcClxLUN8jYPUCVS3Md9vjlAL0kMwMq8JX49EtHzbc
ICfgBbE+PQ+Yl11qdIirpy5zmHsLc8GHm/4L64eOnwM0mxlIgxGiI283NUqPPeZE3uYxinB8f+8L
g1F/76yjapGz4emCLOENGxKTrCqgT5kjRs8wdSnJkFMpJjyfTn3izeatKcbEb7bUpyeVB7Y5fQlS
4LpgVMG94Je/SWArNDsEr7+/gAtJBgGrkBv0khICPD9dj4Tr9PCC7ZK/2g36BAzeTkEgwtDKKkgf
uBzztwXAxoDxqpgV1eOddjLKHM3CuEOQHoCDFHLlQa4H1CYuV/jZMj3jdm1MdKI3fR78VFSRXZ/0
7Q9MH73o0OqHFIt63BVAWd/UDqIFgZ+AEAp2cY6/DirJnCTz51gkStWvaNSBvRDsN3Wf3DF/f8hW
yyJvQEyCFX1gp6JxVrk2KlUbChJny+b+Gp8zDX27ywX6iQhkjFIDK1/pUYPZtdqA8Fvskho+Cm7G
qJMXeNM7DmC01hppzXXawfTsohRUBsrlgE2/BjCU0O2syL9yc6/C4992VGN7fLhJl4vpCl0we6l1
rnLjxD1OX2Y4QPcWWkbAsRT2vpLQZSDhJZOkk/exmQnVvQ8hAmvID3h4qP9sHQqp3KF96GavNqc4
/2DKy4jxF9d16uYWg2BNM84lG+hnD5EwXCc4LdCvMAwBIUWJQSFfxwaR3so3GIyNKipoNfJ/Kno8
+eXo3TOfHwoszFjsLgG5a1IVumNE7meqSYSHLQ2J1zwfGkJg46EibmSmnSH+ADfcW3TBniygoXPo
q8kz2V1BjBdCQVyTDZMhdVcUpvh2TE6GLXZ6A9+8tHnmFLQYFs5qu+oGmdYjLqTogPDsuihuDQhn
7zH0vqOjOk50eXBdSzGXEpPN/rNKayLoBKdyvepAze0WZuIDEtHWXPk2RB2h0nh2tmwP8SldTk5a
0nT3Y4a17kXrqe6oE6bKvEBj04ncJZO2glxeP2IAG/wuveQfs7D10bjEENMj8Q02HoffLylZmZ5Q
D4HnUOLuPqyzO76dcSUgZqPAU2G0ULjuGNqNwC3dO9EoZXxPplOmjyuXJgNlTVX3MGyJj5xUz8rm
s8tKnqZYdarkf78jBin/r3gme6UUWbgp2F15obsLCPwK3povxp1cGyCMETd2rsgbZG4ottTMhKFL
MBBkB72vQNA+f1FRpcSqnd9+/gf9+CnTAgB3hnf7altBXwe532xli0Gbd7oHjRYO7yh/lgo5sMHY
Cq4j56WzfuTKjdZgVfqZ5ROduZPZYsVv3+j7ROSSQ+ywVFiFkifD6+wZCpV1QvD4IfqepwBhDyAM
QHYmRuASArDBRH6AK4xA4Upm2zLKnervcQUGn9kum8m9ErQfCKZHCoLdEvLJJR2EqfbTaguxqHay
l6chTyjdlrlSgsDlYjZpFQoAL49Xn3AfZqVihaNacylNGvalNXDjtUf4kPOUA3SNbrTFeMei6VdH
LT/bMz8NPmCKDR4syqCw/2fSqAuPE0WxOwAySFvqj4KS6UCdQnp/dZhNd7Jv9eDEGsp2ZwZkO40m
PcAL0u2sJv3leXuBMFvfdgIk3TVh1Thl9a1RmOwXJlM2SAV9/XmAJPnKRre5rrn+dmhZUFC9VIPO
LGxGLEDMKBms9dG59vk1WSc+DEkXYLyLnSSFqZ/uryZnxbZiPzD6+ygWl60TINJgP31wvTShw9HX
LbUz8ZPzoMS3pIlAb+I8+WD9NzBS+GxiBHZ1AL3WypCuVN7eKgEKAjHks35b6YYLgtiUEwFwDGjy
RDilo3KF/v6IjfxOFnOo/wq2cvBq8639aXwz7K1UqgOY5LFa/Uuzyc8+ISYZLxKSlLb4wZxmg9Fl
AFjSVWlGJjwKzga96w75Q52c7knmcVmTkbOcm+/4+tSaD5UCshM6kf4kV4Ob3qBjB13pDfCqaG35
YsFBMXIER5Rt/a/kdWZhGGW85KKgUKF5CLnxKBWK3AxG5rlXxD8JBJq8xCcjLXNiGYN280LMsJch
NVEA6BvZ/MM+WDDXBpyrk1luSIUXVYs0HmsYXdsE5MKGMYq4ANJdQ00hnBo3RB3cIicU5gTrmAW2
aq0mkgfPh43T9VpLPly2OAE477rAWvQ+NBlslJaEYzFA7pfJ4s26VahNnFF9EhyLIDy0e+blstvp
14QBUDj09RiUK8IA0w3LkWVxPj2bx2Bu4V49VAGuqEFj3V6bI/w1z4jREgvEF5L/bWWx2f79y0nW
7qrCYk8oV34QIY4+5rWGiYQmLyZ2i29CRjqWQU/F6pkSUTUcLoKY/D5sHeUYcsY7WhIP94AibRuR
zf8nNh1DTpNynq7rsS4gJwWvi1A/8+xzxhm6bKKS/aKahRyrO3Q8uSptGflFcFLlv97idjwJP0rN
kx8+eKoPEsiE1OdRirORG4d4+YIhrD7HW2G43LABbvK9c4IXIlrj90BIWCI88XwkVKD0S5z/ZAYF
ixIAZ/2cbRrfpWxRGckw0hHfjcGrjGqT3/dXXoooh1zigXE+6r/dJ/1Zj9EWtyL/O4RGEeMKtM8E
2IgIYZFw+CIAopIUvvX6JNvALycJffucXpFYjZaWVdykWVIlvrGurU05ohUgCm9gGNabXilUyQA9
6zYWZtKjIYpTU+jlv6/RjdnSs7YIuVMU4I/mDlIh78oZUVL9Dr4a8MODdSh78wVHyjXXtkgKkVAP
8DuL/4YvOiSKbWkS4f/wOhYlH7HfcCMwvTxq2PcfM9Z0oagwXONAHQ5NYFgblgUWHj9ePZMXWB49
qEo4s6G4x1Gw/blZn/lmv1INWW37elGWHaQtC9BsRrb8YATsWuDowaEtNUK8jErvhO5hPsVtMXHl
bgAqqYVvELleqU/SOnLgu20GUvGiQzM5SDYtvSL5qM2qhur6fjJx5np5lWmCK6rxxla5Oxm57kvc
9uRaq/5IeXBu8RDz07hSUwdGbHGvmr1cFdKKphvPT25tfXaAu9Yu+vzH1KvbBevV3lVjqn7zaFv4
EKGNfI8+S9KD8VD21xCKzAsey+rU92N2CAc/fnBBPBzKuou3CuZYdmcz/olwrEQGRJueuoMbNsYi
EPKYGgsLmyJE9JnPbVv719NRyyQRZtQ9wwJKLqGzvfOhvXxvsMwu1p60MbV1ZW+MTWdALQcgZb5r
uy/S2o1wQC2mHe0sTFhh5QyivbygonS26LkmqQjW9Qyj5HuCy3IfnLbeixTF/P6CwO4L+0SkId6m
uUyNsQ2jmAqOCkw2CkV/fEQzgRTLqmtss6xS20Jl0sbE2BiLnY5Mtfz88HGSWfTYj7ZIFTT8u25r
TTzefECkFFK6AZeFqyymL69OEcbVS0gwCXjupVdAer8/A0gIgNsjxvCd2jwQrmbQEL3Xv20TF9hU
kyhPL/FXyXxMVqKgwttx6xG8Ah1jffOfNNlp3X79TUBfK9NXePuFPN0829kg4E0g/KTZJQhrutqw
kacDyX9tmXoxk5rBwdidYi6qYq1V4jnJ0RAHwRatKxOlnXxATA/6qonmPoUk3jJ6cwATHquCz9Ed
lSN8TMfkjP2PJZkxGhNhY5I+9VOKQgZKfRCaDEnlxiA5iWVnE93yomHh3hg5Vmzn9XykOgDno/oL
DiHzRyxIcblTEa8neDNnDeQ8H4XV8eJ5uUsKBVP+kw2+OMM/ctCaGNJRe0ZHVotzdnX0JiCHE+WD
m1qVS0JwKnvQBUQKKxvsocAT0aUdt/VQo5wqdxqy8GLgu4fgYZKZkE4rBaEFdZ9+g+jwhsGjaePC
rZM1XLEQ0lABII4LyONMmSxvW4c2zEjwyanhgpg3HYWRmYMOPUN0LaG2DoQQY7DCgKXOwQA1ytRk
bWTkVzNFsQSwAweC+QtGOE0cbyashhScHeG63Y9I5a7MJVY0IsTSQBei6QkSuu5oMyZ7+f/nVszp
l/d0r5VuO03R1QJ8AEiG8AV3o/xr02AXpqSZeWXQez1PxxjOtOGuSuwR9erSOa4WMlVbSKd+MYwi
hcAIlpBKugZVz97oPdiF0mYUyIQdHPqs9mmRkwGnUrJniVBNbU2uts3AZnU2q3532NHzjen5zlIC
r4LMDBZQxND4c0dLINM2IXPTD9cnYtivsaeXdKCkjyykqYHoVl6M85IW8Pi+34qSrVvQTWIhPiSu
gEaotRBPoV7ah2P++79IZ+nl6fmU9cUXYbDP+Cmnl2mRxzJoJ6nIv6CeV2nFA+39N1/0HYyf5HNY
MsPWhrzTYV2lNB10/9GyTQY+Kz8FUHuugofGy1KPRlykgDyK0mJyiurQaF/B0WLiYiBLmq1PQO/x
mZ6Y0HTxKz8KG8tGCElye56WI7uyhhTYLaAy1U+hF1uUlpo9ROSPqskZ0UNbnhomwPRxH8jaVU/H
msQCcvds9P8JtpaucLHUessvkFV1EvdlRW2pUv0MgMyxURw/bNptMRCmwwFoQ/Szh7Quem+lQzxc
gZCs/UZMHCBabv0mBSsiuW00JxQnSW9MjY8l1M25Wjp/pYswfD70F0a6nYwqTqlIK7VoZ0Fwtabq
z+Wd+01Uhj3h5GRb91rT4vyzr0tOzDsgIiQFVcc+zndKfPxeb3QiZiIFh31SyIa+V+UgSeF+b2Wl
VX4+J53L7lwdSS/dfT8KTpQ1u0n290s/YdrLPlYcoy6VhRJuFVjtlHF7kI3OGH0lO0rb1I+0M1ka
em0la1x4vfT18OAUbVDC7ck3bIz9vkcpBmdz5pPazSCVhPqBajJ73+6UBKlb5FOWk2tY+IdhZg+Q
WdbodDc4jS/arfi/Bez3bULRm1bnIMswyJlJMg0IpojNpbFDp1lci5zdtrccZrQyGxhOlrRTlfQz
RoVuxYfz0dY1ljkMHk25BAvTeQ8/4MqYT3Kiwk6vCyRKz0Q/INJoImgbMaiQ3yD1Ae+u1+7BbezL
KwBvG2sbGOttrt261k1Botx/sE6+21GZz0U0IkVqM/0nYqvLWPvfl9UdnIG66DjIA2nZ3jp2S9Gi
iv3tCAjCXiCXpq1KTQ6f8xMEejKS/ZqXuAO/41I2iDG4Nhq/EmASrBzNOmzkRuZIeXb/K4YMOnPu
hJo/7mdahWHQLw0nkA7hHfoon1X0kNQL2Q4pnWcezD1lnkufb/WYMIskrN9E89IrA8KOuFuch4eW
gyBXtsWZs+VTHJuy1IdrVT4okglC7BQoyJXZEsiRmZBrIBTV8qAxy06fyJ7ZJAQT2KCuxmHA55In
Nj1i50vXEuXa5cQCJHNYKSjuwOw1TvlrKy4VXxlkEXt5o/Ya3AiME16zuqkXXCNEqPhTNdjgrXkB
BY84LToUjNzFyTXFJO6C3fwk2QSauj0IMwdBS2mbi1nPOWSg9Yq1HWrXQpqSg2aHH4469ldf+PTO
T8Umc7OCS1sh/hm0/8a0G3Bmx6m3pKxUPI7Wx5Xx3QI53ziWRMcbhGTYG/5dZQITqhrqSlWQkDYK
O4jx502RznxJ8onURqBklzcOP6CGkXi17qXi2Pv0jaNDnuOxGak3vZLSW/RRCGDoxyhrEFF1yMY6
0Fv6qAQIxWSVYYTiD1ZCActNu+hBSBTd4l+6MWRTmPa+17oXNPH9PDHRpMCUhoa+xHNfvW7Usg3j
R9S5iSKoxYnp90omWBiaDw3gBNmdfR73/kp58irYxiH0NR2Htkk/o85diNzwbUyL5pNlVLYiVMo5
NO5njNN0U7OM5Cp5ryEx967dqR1bhHLNV9zdZkVL1IE5EpLMPej6SJ7b8CH8I8HprKUinkFW4hw2
Ot3r2TUNj4UUGEtzfFZDCg2RpmoXHf9Rqs5uwvxb3fbPzfwdRJXxergcDvlpjDP1Pu35Lgs+m4cS
U+TDTw2LMzOnya0bQcCOVcJbOqs/xI/bwMAVGe0SkzUoK1DWxdJwWOhzSSsvbSWn0eunv1vMKo+L
vyovY/zGQl6kPitmKvQKsGkXR+mH/YUqnJMOTlDiaqw3KgktFdPOua23Gf4RrSENnNNfxJ08RKNM
tyMfXW+WITkOnjOcbGaSlwxkab3EKTIKwhycr+rn7zKW51j2lZCiUeoO/RzPSqI3WSnNIYe10uiC
atFqBwTcBmJZKwCqpWmnSI0KNw4P7bw+/i4w285n6iP9OMNgle+lO+UFSsJXYY8rAkBrtqXIb97N
NpWKn8OYdXkGUdc1Owq4v9HliDrhZbfRpLUgTDYXhUc0cYv1eqHJ+k2mFXXWeabq4ZI5uPuv/6cj
ktqbsEfHMBoyqh1g6PiZxroSiygG0LPJ8eY3zXyBqLw3mUaIIxh/Gomkb0SWx5f0HibbXFpJ2CUk
Pxp96ulUShih5+gb9b5aMrrVajM1pagrhPXzz9XKz3iC0sH+y0YDyseKcWvfvbeUtG+ftPw/y+tU
gTKyvBL3CKi4V4qNeZGjihiylgbC14pediCf+ntIDMd8SMVjGqCGg9tdlN/44cThONfnfOMJaZ0w
b/R8JqvjSCyygtk6UaBFQhCSbJR+n+KJI6SNbVDRtpLv/4Hid9Gq4bbwVZdyvRpo+SjC1tWmwpo5
h/xsos7E7S2mmLNoFI2KApVyQJ+sQ6t3aPBXtG5MRfU5pClaTzVWdRmGSzuOp9NGwDvuyesKQCon
xvdyB4194qa181qsceU2JePBQCLQH+eHP0S+Ay5Qzs4RF/JzF3p9Ie+yELYYb+iRevZjlJzBStm0
HvtDC0lnPkLj1DOEFnbQqcY46DRa5e+QcB4qcwMDgSPY1+OqMli98mX3AGibh/0czJeKBBCjBRDX
YmTTNPdvha6UZtK0EQ4y9MpOij5f2H4Efgu+28PIWoTjvthUStlHAlXl4K+aDUMQd5JL6YWgovQn
UrvXVDIWlLOXbpcVuDxoLKf4iUIOstFPkSnG0234e9gUnusjTRFL+m8jUPWnr26ejEt74uTxzzS/
rnrPn9Z4R05EXYr7qZr2jDwn/pH1whfM0cHcYA7T9NJZBH91cG8qwe1my546J50FHynMfrwYwleU
5Xxu5QlkFhX/lXAgM1zMWTvEZD2ovW6S1XueSBmqhKgXWcJShdh+oBXYtvAT+5jkjHTcCg4A3Fps
nmZkiUr7GOBf0Svn/n+JeYodzAi1tODZqnwjpC7JqO5fE64JqYAFgI6E/PYBOm1mkQEPZawumtFD
hpvyPHX6RBndp1dTMLw9ioMGvogGsIv0e61VbyiJYiKQxeU8iW0+JZIeKJFhM6ALRahTpFnPjDkc
8NaR2ilAg4PUfHR1hwDbjbhcPaiLX3xWWa9bTI0V7590tGyCHPQ32RqJimJOnfZanqJo29gE65FM
wh1fla2EPiubFvTWXOSbNi5+gKxixmLYOPg6v5+UGIS3oCiVOCS5peZUB4ph3KnOuy3wlJQtpAE/
7/unVzR1iFoO/esqyodDjGP/KDZFmgkd3rmYO6UBhO+YcJvcRD8VoPlesXhNNAaBtrbCrKoMuUCI
Yy6wbur+SJmG1gWowHxVDvo4G8YI4ED6CMt8pNrOt8/Aqakf02IZcMyPEMVN5AM2nzJitMG0t/K2
cGUV0Rysi4VXWzH3R3zPbboMAV1yUwnpf+LFZCCVjcDMLE71S+/AykcG0GZmKul7XIZfxxYChs9q
t36Eu2p3IWyryfV3Cdd24ioqUdgseUr0lpta8CTzjIw0zUrMopltzsiikYF07gnJuqy5XHdA49rJ
tdCz8xZjlNNiADEplpD3aUVFlPayk+KLJffm796bVF4QCsXJGVE/Q8iVGIH9VtbgbGnZ0Oa0KR9z
tltPzx8+UkIUPqjoBjIeCpoVoFoHs06ORL4TuDssAKFevpnuFJHZlLZ4Kku8JDdfSDmGW7a22R9V
QWcqbbc/cfPMQBFRWBFNQ4zqj+VPE4/9h6ba0tXkgSFvAjtguM8ELL8jXjGFC9qsCJRWh4qY2Qe3
BZHLm/vLI1jP9KUI4Htx9PBUnYgbTuQjBe9dpoBaH0UqWKvQ3azLusr8VvjM78ohjFPc7fpD8/xW
BAu+6BJIJ6vY+XbALbI15Faui+HNxQyU3tBC8Q9TW2ZtDf4grfyKjzu4iBohrbJ5p0UhHJ5zs9K9
2VrjYrW66SZnOsPZZmm/quWZOSyKNzJ1JfrgMZ5MzIYkVAI3RiA3IQZWixVekJRW2tGJaCAbLUKm
iLiY0mlKRfcwZifjc+FEc0pL+/oyv/7AgEjDnVYknYVOuBKOprdXbAtZ4F+M8SBhCv5WtVTliXkc
GzBVMlQe9co0oGUUf0SBYTGkZ5eyorMVyNGOj/nlMr/QvJsK9SmgPrbvnYs6RNme0s+D/jhDQ9Vc
j1tCJ9AWkf6j+4UZvWLJh5ivvVb7BkG0JgqJYKRm/vCW83Yi5D1xvEKkjrDUqm43ASA/4+ecrVbn
u45SXdHufOTKunAQ7mjrr1mm4Eb/2/Ptr4B1dByUV5PzGoKCtGPc5/GUxJbb+a6DsNSMUqLdIuUj
HaQMP+bskI5zwEJeI8YQVjtJWWuL2v7lnHLYvYTi//cLcZBUGUQ01V0ibXPUa8t6EmJ/eDjKYl9Z
h07vDj3Houk/Ru0t6mh7qPND3gc21y+nL4rLZqRV4zXYHyy9e8DjLCwtYnnzQl5jRmHo2oQQYGrT
4BF6ClEckYh4/GD5WckYHqeYG7S0XyjGo9OwQ6CzVNXDgRdLAkzk4iy9y8Z6sIO9e8Z+8bwKg0ip
KFE/srbZt7PKG5/phl7tL342BjfbjpBxLclN2HaGITNRHv6AEEy2BHxZdLrI2wLG6gNRo1Ln/OTe
GJdwE43OsyrSBo/qrKdvAayTHwdzEZ9sytraCQlbDlnZvV9QA8SAJq+UPrEu4gv0fPtnhIh5o+rk
orYLsFjJ54Tn+3pH2x5lhmmmpjWziZWn3UNID1QY5uZ/lH8u83G1/9FaRyErYAGeBZPia7CWvnOO
SsUJiU9E3H+5Jk+GIsP67Fc6Pvy6pqpOoFuOjOj3O2H7UNUfEFH8I6KnwIWpINg7SXB9iOXUccx1
VlSAvKbY7IU2ifU2Jv8SB6yWroKWF8VLP6d5f7dje6ylp+JijppTwahex0JbuMAiIQtfXZO2h6Pl
x84h09y/GNpVKmpAwpkHFXOlgtbMUiOuWXzpZt3Et+BHCNJo+Uj/Ro2k95HkJoymqA6Pmv2Yu5kz
EMAYIQSCyC0cRs1OsO851Xe/HAoWEtB5O2hfDp2AsLYpCT/PXnZjvoJ402J/zswKhOk9kqflpCMO
nxVXEzqI6r3lXZvrwKVDTYKopa0FP3CSTYkhSKmVirO3KrPWrnldugHwQrdTTfYKX2k5BwWub5Ap
Q1+Ec6sAKEKYb984mUzVvv3/j2GOBzV6FCWwytDhtVoAWGjswsNbDRh5+Q5KCW0DV0glozk01eRt
TJMr0xBjGAiaarjCIrgjaWJ8h+GivL4WpBOrWxR9lnOEURKN0fIwNw9szCLnMeNKBJE3n7tz6OLj
crLaTiHRvjknsw+jFj5pzSFNFb5PlFk9Xo43yeKz0JrDqmUtQVAaPs527nOMFMRaSNhNNlyMec0d
s3AdObLI20g3K0x7YyRmE7VVVg+Eoqeit3i0Kfpyz3BPrOzfd2JBwmg/onVpahnJd1c3gQoVNEYv
RKem7zl2crrcBaPpBMJLwHWk96W13beztev0gV6TPbAitMOR3S872RPYmoszPhCNNECfrc4atjh8
VmC+8GGZE4NixxRzURNkh6jAuZD8pCuoSCFJOOZLdtQBQO+CzH58HuWVv276v1kpNlgHKnYITUoX
0uga4DEQ+0noN52QTYGyV4+luFR4DEvPYMA93wSmT8KmLv5S22/AZG9T61bW+aCfXsqDJe9TAMG8
fRIU/OG08ykjU29E8j29Z+ayygEDtYGpbRQVR4NSeDzNY5uXJxChz+fDEyQwIVKbKvpvipp16Yhp
2vUCvujUpzE8kfTdBpbe0pMtvNGBbelfQr7/nbSZs1DcfautqgyMTeO+i0ALKjTS1uIwoRwFqxBz
BDD49471AUB244veH7u85NSyjsOhqAFAJp3Oh9LBhuNCZ71qJy8oAShK37MGPS0KEU6SnOPbL4Yw
xovX1689rNmzdbKSDTylU3YhnjwdjCCawwiLpTWTHBf80WMkXMMshPVRAZ1NyB5l8lRxB63mo+ho
5HknXVF2oci22b1BLbdxDw0sowszBlICy4vYTNPhnGoALRP8pwkwuxWV/MuF8EOPgFWOGnN1s7Ih
tK8qEbhLGsqlVZsEogHGHjEdjhwzry7/Sd6nEwXw/SEKT2wp+Fl1DLhWW90jz6p8N84jl+De6k/A
LRYFyauaXpM2V8+uaLhQe/lnKTSAB7giI11dknuMkoZ9QqzSreuTQRCcLaHN5yBtpytpe5L69dxx
5YeJCvICfng3/T57GWZ26DdvuhNuuKzrz7ML0bP9mYJSA3EZuTWqDPbE94eeBz+5xEHDG332P05S
rJr8OGRTE6R+pGVBSaAB7iudE+B1Ht7FZUvzeGvEyW54KDKEzVc9BEx1ZlHJ66NcNNtKF7dYQzcC
0n4RyA25EOm3Y16aYM2pYKJ4sDniEDZTXxi7VILaXGwm6rqXQGK37juKA9Iyj2nyi5dvVnYebIE4
AIS54kxOazNF8y5YC6nnhCZ9zZX3unT+dpRbOkAQUkSL2qz092nrdvyqbE/rqDVAr/gpni1usD07
vfjn/czC2L1HRkxOrPBObWQsQ8IAugn4mjHjRpdMVcImkPnScfq0Pa1KPh2tVJje+ETKuVzWT4wf
AE6Ij8jbHYBeoPQkhF2CbkYueZikB0g5f696nzW1ZAZVUN/juUananVNzYeTAUlobp0OMt0YEjrw
QKtc8Eu65siHxK9Z/0BqROmnQZboY60z4+wgHP/XVRjb/Feoj9W3e7O3VoZ2QA1pWBXVESaO0SJR
U/IujDJgq7AiAU148vZo01BimSO7xB3sJbttXFLLhBi/0S22WiPa5YuPBk4Rkyu0/PzKP5ycsGAe
It9PMZkB5wZdQWJh/PadBn/f0jUbDoFJCD1OBkcQAzcApFU+5UA2YBERrUue80hnsjIiX4cZQAOD
cRkg1E13p3EVCV0qFLdlbN5XawGZHZooMWvBDQFIGTyV80PrCiIPEZV1h04PtE02TTL2phwk78Au
yEnWpsjrlhyDVsa2l1ku9LzG6+j/mjOgxsi2O04qYX35VgdNdaRHwsrW/LuULZw5JNnrVwUC3y7+
W8be/7kD2bUajwuvhmUx82HBZkzh7JkrHsj1Mvb1LXWupEZPIWhBRqEC2cMMd89KZBD9jMBCEGmM
SKENzpOGDTWY+s3Vr9EkJvJ8zCreyycU2UAv9c3HrWCpBQNo1LcQOQiKMLuVcQyA4uWrFrNS/k94
vphyQP1MjRDeEgUkVoP0Rv+hxgy+ImNx7Hu20c/VbdWFvJqRnuPibQ1rFqxu/QHP+CZyCrvtpYwE
iNXPhwiYs85yD85wRJs7X7+thaEfOer+E0Feb6Vk3aUwqeDSmrhwOsQ9F8l+x2zeyaUkOta2Z41O
4PoNWNZTN2IBCBfrulrZnf27OdGkuQBVNBlv/FX2nYGNVA27Jf9j/WGz/u5+4KVUq8hlj7FanGLU
JU3a3MkJpuhgf7hpyGeJQ4rFGOa9GxTKlt6bPvcgNTqZigltNWekzEE1L5v9Ju8ORLreiTtiwqZA
d4UZ2lzJBvpxM3R7vihWz/Cofw96F9o41Egymzj7tDDKx6NbUPcuKXDJ6/SWElCqHUYEXqG/1NZV
NSyEEmGXHoJR0wRVhCrxXc0trNdCJIJjIou33Q0RYdQEIqe52D22TXMQUT3e7PiPujogcwQ/wwOV
uuks9mpQFGjLjeEAqi5YoRfRVlX+UDjWVIyTo+qPGeIE2mXXtys77Oysp4KBqVJw2Y0XI60IH0SH
gpFXJfqRxTTSB4uymB3Lu+7+uUS5p4zWXVSDp/JfY007Dt5jF7m0DfrtAyR2gVfiBeGi/0NEMh3A
xLWsYpDLNJemuBeLJOewNWMmT0lx8fqjacSIOx2k/rDYV8AxTP3vxGdVvsLVNH1nWbWFuYguCgI8
n/Onz/Eb12yG7SOqR55bvyW3fd5DrsqUQZ9rpP/n9qu4ubkAbxN5YbxCVUARnTi60I9QgIckCbgN
S4nn9v/ue9uo5SSNeurKxjzwvCSjD3hmej75Ub1sxgLIRmHAljBYX+LNkm9H8/YokcI/Q4IRWzZT
9XGeg1vODGhLzPuyzacw2a5KoFxGtABYeqBWlujAdhLcZXeW3qG+gb3iFhGoEwo0ztZUUZAycSi2
gT9ucGGKMXJ7xOS2hjRW1JMDAZAlbH6f/6a4IbDuNuo2ChEwMhAQJK5JnSVJz9MOvzzcBZeCRJch
JIhfYccaCx28w+2VQpPMwDPJQCp4+m9ZcD/B2sfBtyh2OmeRWEmaf8Z0J3eUn7PrfdabazWNSn5n
9f/RALKfLDinetSSPxKp3rte3dEQw/cBEkpIw6pmDcgD5TR6/B1sHVrXuiCO5PmZ2oLkmjdC9a4w
DjZrx0O1rIy1QDiRl9/9PPnfve6/jvJEWcNURCJfTr0M02SejSqjj2wEJiBLoxoDtYi7DYqwqBcA
o7hoYVxWwxzpYoi6E2ppcbL6Q28XgS5/gbiARf9QZNgui7FqgaMkRS3W0fXMUL8HsC3OqIdQSYPa
uwIdvC0CPj78hq5ZZ1SyCLPqM7W8G/pYnPEWN23jLomLjSl1lLPkxVjw+EVLLOUHOw3wRnv1yL2r
Is4bfVEHE10BVWJXFAo/wOFz1X4HHeeQjQww7n+rHhfRkuZnrmug/UoMLK2qOozd9dWiJwDA/gt4
lZ2TK33ESry7AVibdEi8QticGB4D1Qhan57d00ZtGtp//DKjWyNvhDpUpV5r7fqsqDlycJOOI3O0
19TfD54/6CM407Q2Bl74Vz3Vf2eLYYbx3utiM5jU/vHjg6WHeiEy31nE0jF1CYlfREvSAg2Heajt
wyuScSOakM40pC/kNqioZd8zIIRgPwkzINGSHrPKCSVvt/crsT1kZjpXq5A7AbboRLTOgFgPlQA7
x1H1MuBtxmVb2CCpesI4OIrZOClUZVNValYqXdckTmlAVj5nCJ2TJ7GUCNjyg6YcDEhUkWitbtAC
FXQ03n6QvztZDv7aS91R7uLvpYjDCBe4vDvO6aM0q1BPVybz1P2YFIJw99albjVVWHYjcVYqiNfw
C3Uudo1xRO75iOPBQvl2rkY+QU5pJjYU6XUxZ0+38Cx+RoOdWDy5FcWhTwt+1x7VTTe85M+wng0P
2rcMlqttX1Anl2x1NzAWQygCywI4fU+yyXTNEdmth3YsFC8eQt9f2rkMD/onX0ozYlva3U9WbLUj
hzezjOhHwNDOew19p7McgYea2mQhghJ5DBgUTutJFRG40byA+b0iXIu1Foqc3hQjWP92AdFJHOX7
A3dkFV/11xKROH5UZ1ELtAcjLrnjoNYk08yIGSOPEUqSUSSnJHtVmvGzGn/TKlo2NMskoyttCyJR
dY4x7dBi2Tbuqw5ejc6D5UziZgy3CBUIxd5MZIzV6SAdGShVV+HTgO23tBYNve4VckQQlNgk/TYa
pUWyYRC3HW1AqGJ+2F7Gt39Div5v75g7TsMAzvVfrHAC1kvseST5Ibhjl17n7JIOW4o5xsmX6wc1
lKHf/GXGf8h9UkpxCqPsTjhSymcJWnLnpUEihSlKXe3YqCViQk6Bjq7czZIDQfSSAVm9oq0166cd
ODZfvpUlTX7YAkObUd9iu6+ap+1DslKOX2VBy5j9g6LhIAX6wwiWU2bM8DVJ/Kem96A3Ud/DtcBE
LtzAdwZCMjdjeHzZ3YfpdjwlNiYx3BBam5AqlmGUt5BKAiL89cX565z5TolRGuZlqRIzhsrKREkH
EdTr+NKozZsxiNoRGPfypuRlLfvC2kqWsBvuLJeq45OatLnlezVd8IQ1ne3g1u0mVR7VWUuM14xJ
LbkidrcmiJkXNZZ3/c+OV+CjWXMgi2Rf5c9WgR10qYcutuIuufkqGQu9AxmJiKIbs5z8gdRKNAzc
HZcvX4ZE/dWDqRAVD/KHULfFwNJkLvyp4IQzeclETzL8lrENvHhr4fMcjeq4fhc48lSehnfLNk2X
k8NzCBxFHsC3lU8LAzdb56OdwoaZcc35aU/q5VdiKU88PZSNEm8w6rk5x6Fy5qymZNmTS/uS44Bl
CxpFzt9VwNLiOfNkuBAdidmkSMc3rdmUf+2eX3WbZkXXfyBHag9AE/Iu+O8zCyNc9yarL9GlYWmN
vyVTXhKp9TS6Ql/B8zCHNAe7WWprWePIE7LkGd2xlu3iGFaY3ht79XAxSPkuJibN2gH1VJgiMjZY
/ntiFMqNxCNOXiUzQpFE8LwUXN3Vzrw1tOhAXfagKBypwjVtCom5TtGRH8if6DMwg2QPOH1OXgKB
qiezkuYy37R1o/beC9sSg97VQeGZ/C0P33RUQEZtQti8yiPIEYtKdHObpbh1n6ycTiNd4lGgAFWx
IhY1ru10ri4PPyJrZe//a6mAbN8ZcGbfrc05qNGMpOCKovuvlB7YJt9k3+2IcRoSDMwlMB1h0CcZ
6FKdBXo+RQPyIEt9YhLVKQnzRiANq4Me1bWAavC9sAPGvC3W4sqvsrmAHmFTKumHi052hdO2JvY9
SW/boH3EFXbEwwS/FOCvtZdRe3zgYSk0zzx5/Wj+FPRyWNWjfBazem54TWCUxIAR8OzoBilA2/DP
8GwPdFUwgai1f8F68hx/YmD6Q1ERtgUtF0nUCrAsn8f/I0yEvwXiFVnWfY0rvVu5KMsSmuqXqOqy
ByvA5dISdwq4lflC+LhtksLVp8r8fmpvr1lLxhy9Dzxm2WtLEqMfSBdFHXIOWZxE5NZHM96QBeMn
NmGONj6FBGum24KkQadXoBvuPZ6YdVMuJuEadaIylH4biPuPXz2+V1Dmsuszc0rogAZ3XqNgrJFF
F3rfJYswfHZeQ8ITvpQhVD1VvzQNTtGPEeEs9UkOzXGU5ee/1buZ0biDh34ePpFaq4oOt5cicXb0
KU8smviPUj3W9oRhXmhSK+HPFClsjhqiMhGxoDP7KwwTN03QS2O8bwHfCaJZ6QTXPKS7FGnpFVwp
O0MkunYk9G7IZwYr6RD2RUPUSn0qTyQ1zd1xne7AWuLNx3znhSbFUfu8usvK1dATllaZhigFKKaX
ldNh59lVcDNaS7fsyWFAehHz3nFyCormyuKIbX1O9J42xs3ntDACJfb9D0yH0pLwLc2WPq1kzAfm
a6twwL26ccRwJHIVqzldlXcIQ456Hxx9oY0BlXJqLyahhPjWx4c4PbE+k4BV71bRD/Nh7694uGK6
mrPqIqjNP7Ls16H3bJhJH360icEhIm21cnv3FnlgKGpe8489hcqg58pS2UREqpbxKbiOBOOb8kKJ
AoKKiIaqjW7MmMNFwGSXDiZV+eJVXg/Qi8ye2mwPh+4E2H3lJrwDC0yJRJWPFxpvW2WKpJtBPYDX
p49gncGRYQVA1/AAVTh6+kQRUhxzBaYWz8njs+x6XmFkqWTu9CBTfBTY+wJowJ2lDMJTqWX5UcD3
3suNa/YXQhxPHcNuhqo2quMuoqpNQgYFIaIgjoKUSWIKz/WeaO/wIBaAd9hqs17tKR5tHbPPt/0A
f2HZg8ZfkiLKAp84XfEfTqdWs6Ool9vkF/k8fAkEk02WPJrPfwl9YIWM91xbv0ELtqZFl7nkrzUH
0Tuk3kIRNO133faahff+otH/OCSbuUcxn6a0IpO0pnW74ZAfaa+FFlaONgRkl7AaOpfOhpxorr3U
XSMawwsMAJvTFNQAOUcGqEu+JibROESWplDDSqQHqc5ax3bCeQwSthNitvQrAlt+R2lK8sekXQJq
65Mj9SAkzh2mU7LRZ6VsmgfF0uBV6SuXsS5SVsanZZyMQv1t+nl0EDUJDQgbuZqzv1JWR6JP5fgh
V5E0jHmEGKM47Y/EPqefg5vh0MuAcgiEMj17gRk+thq2WgjD7I1wiYCn0jjmHJ5+VAKn7d6oVVHG
shXsGE7k/fQd29tR+MFSjxzoMH+tZclfK6OK5HQUMdQXB41/Hnc/fbLcyNFFuVAWRy1LiMpEiuqF
+ceOtTceejLo3f0TS9heByLNQX46uyClcOp8kU/bgpAkZwXEnEuQ1tasGFsNrIqx9s9BlPxXcO3Z
AHcycuVDNuz89+sq6r06FGjyM2OZctxv0vlefeS+oXiCDIckZtU+JEvTVGzNkD884JTZJ7N3BOR8
tWWLQMZdSM+/theAgvw0k7zDdaBPnyOdPXW3cK1IT/doikWhGthg1yMijzsA9Tdlpm0IpjTymdfy
Eey76DS76bq/uLzzbiFCndR6FTwIy+8xlqJNg/DWRAgQGdM54zVRllk2aEawi+W6uxLIjyGEOfUw
DMR6DHHgD8/sht6XcJWJDS8oHnZE0sYS8oWrJZtNN3gvJ6xXedouk/fMkdqLu7qjaRjdj5IU4ntI
hhVVdfBYLbpJKmtlPQyZAKKTM80lq4nh3t6Q5yJ4aREvnxt633rR8bDJfe2oWHULlxC9M3mdtRID
Y09ajPf2+FkvGZ9zHYAR6dwhaFsyRV1BYQ+sOGtOYKXYLRnGzq4Vu8psKIhpeSRwH/JPlf2c4EEl
tDZQKxjz5xP6NTVlp+M9aSJRiWxA1JwjPTtuZlKI1U5sE9pQbLPlvmxvlhUioBgNjGISwmgjmU9C
ONeQeNFGMNc55setyByPDa3WdQujyR/cRMjhK0PGnmcB1bmMCpesai7+AuKfMgwYp+V+NqbGN/Fd
zJ6sOmvhkUsT/+KixxKqh2WqVIcJuW/Rs9EOL5xGx+ClEGLsDwesFQssvH8BLTCRXAH6vldLz3k7
r2X0Y2/gKQLRsUr0EufEapN9hDpEWEJeTwa39171rAHsVbJUQHR456AOOpEvoG9zfbMINZDPXeBy
mlt6vSbOqbetyR2NeI7oaH0bIerFVJOkVRCrc/p7R8d0O9AH0zX6HWeL41EqzTdhk+XsE1ztJuod
Qd3iTdOv+UQhwthYtrJd/+mJRvc3glNb+qayY6kcpvdpiP4mza2pJIACmTXy97hmDZse6/XQJFpQ
vmtr0HRT7opNcC9DuVqMwTx0M44pzhzNciRK/Lu2575yZSSCW2s1AwwmOb7y0Iav2CABmZB4cc0v
V94hAiPQMWzVJ1p+qyG1tOEnSCPOeJ/o4Odm3L6A5lDQZZnjGk7xZNvml5VmaOIIpwL6sRj7zKiT
LYSyyJWeyu88k0MAOoXlFds4zX21MCvU+GnnjFrxT9wffS7sFQ5GUKbTooKRtyMcRm4LWqB9C505
RIvRglllHgtFUYrwcRwjScFcT31Ix9OF0QoumuE2/uwpIu9Wovwto8+QotTUY6QnrwoYyu8HSl17
+dFmLHujtrVRP45zrRRj2hNhp6hrGfGehCPYna2iy+88bXxQvDQCMNf4I0heORo5pgu/qhDdpu9X
U9C5d6TcweJ+MFyn8vOluRFOsEMyq02+UINGpdqxDNO9N3fHZKmJ9RzGMW82IltyM1AmF0IPRcZy
iCmkBWBNUaPRNVDZLn5k53ulpH5jnUekyujuRc+Jcf0ehJFCk69QBkkyN2cNiESmaXVt7KxQTk8S
xagQUyBs5OEIrCqDd+z/ZkUWAcTMsLZxMb3gFGidx64xfzIDF87BrWo5o7Cotcl3TjFt5xFLEpX2
1yzEg1gGcFzXPOSTzc+2rDTmeHPOLhWTg2HCByUOXjwsRewRcZJvqBPqQMAxiklwdxv3vSke2pTG
mAnY1xNKSqAqXxK9vxXIKItsufSli1Sv1RPFsS3l9KPLNLC7BBzl9Z4s+5JL3pUSLR8a70GdWppw
DBl7BufVvyHsZNDommNe4uOQxyqvBeOf5iK2KdwsjF+D8e/2mMxTEScnYjudLj07dEJuESwgiza9
KlcSw+XIvk+Kn82c6LqypdRPGrowGVQDcHP6nodZT02VMQ0ESAagxMLWqmiavu3uOSol/UxpqyKb
wIBEBEcb0KPp3vvqQKr5e7V7ZZrf+F+N6QJd8tzsqS4NpVLJaj8jNa1Ib051kgD4hhq3/F2C/HDr
qvImLsD+bbeFjlOd6HEqs0+xgtiiQ7ovdTiClKhFjbd4lh4JWu5lEt7Uyf6kqpYz4AY3jmzCunJZ
fU02A55EHnv0KYa6MwqMfVyxYnbl3gYvRHTeNtSJ1WCStUE+eUnE1QnBurbi6D310LilksvHJrGG
0R5l+iNW5vfgd5HuoHcapspr81xBFJqeH728IY1/tQk2uXMZVUaxVT5LXxSXXYTJ2ofBFys41d/B
GbkqOKg5CBpyPzpCd9kf0Hr7xSHSIM82EYj3biTxmYearU8ywU3x2VYobkST5W+UZVVnyDasMc6U
r/0mz2aJPAb5f4oGn4IJHB48tpNKZxoZ3CR3ffccNQn3wvPDRWRncwJmcYkP3+C23PgCj02nv4rj
mOf4fbZHUDNxSi4UKJPWmYbZOSqAjl5oHpCn4jmx+mADcJh1Go51kn3+240HmBG7YCfOixAUCX9R
kZLSfNspjkCqb1Cn+1kkaC4cbxumrTMfYPWVDuAkj4dqHXllEU7IH3DMEOhRjb5OjPpowW4LN7NA
sdidYUHoK5pklgUZE9QcyKmQ0d3BagBxjrVIdPUv37hFiWhcaBv25V19josAIWIcIDdqvmgPEC8J
EkUOvUvLWK7L+tEUq8BpFDdGMTUKZxNfEgkbTZyGs7+9MuCADJhOmcrB7Thsxb85qH35Rp9HtvAY
ewLpVGwNTxIX50Qu5tI6hBiA/Z/U3LGB+dWmxVq9yl21plOddEHWsw82cWwNIOkF+prBsRFUBEDU
UUpE7KfyEG+dsr+LvnbA2CiK4+CVq+Q1JZr6eNtqeBeYOngj568q45yanmFqPWnAS4tU1JTV30js
G9a0omFiM31yY0jI+BHyVJa4eG+sfUyK2Qt8eTXWnlRtlomYaL77zod6bfVpJ6mqAIUDg+yS0PPz
nLqHgKc+DvnRH47o3X2oqAZKM6rzqIHfIqW7I+i9DQHlAqYuOJlPhSm8Yd5FBWv4sTKdue/VBWbH
Px4kD3+qtiKH2FXQTXjkDnQAAaSutRWWBE8qUFkiJgBGvZc3TWnKuF41t1OwJlm238kLwlQKpnMt
qOoEaC7J2lNYHKZ/byS8vkhcGs3NsFcOTkCJ/uKIslPeGZIB+mJF9dHssTpFj7YE1O5zWKwIJB5e
PKFr22lpn0xHYRxp7qRmsLfAUfen8L2ah4PSxeZlfl/rl9lZ9MBcmceJegzfKhuM5crYwIuDoi5B
roe3aE7MkuqlDZ5ZPwooo414B0y5GANHZ41Q4vWILgM/DxbUo/XXZBniuSm/rjJ0NigcCHgs3wgM
ZD45rXV9IAGv17KLeTLxazMYn71sTNrwXmJ2uEPcwbK5gVvrtuTWQVVZl309wJeOq8kidTEf9X3g
6TjPUy4q1CrbQNfXqZvECHNx/zAhqA0wSJZZvliCsctEBEWYVXFttyWrrgbVs8xoZuisXWNS3jmS
1XfCGbVF3Pdz8M3AUAhb8glA5Mex+/2K7y/8FaKfEPZm+uH3JGXJFtm/ULLS2iYi8up2EY1d6xKT
3+qK4fhoSRn2ZXkxEPq0YlYhaPNFMx7xzgfjSGYIZLHnZXkwJd054UjeYkw4OajMfRRIzr/ShCb9
i6txKgDLaQmKYjNcLSgAjFOz0ptRG/2eWKajYItoTazam+RF3L8MDw7S2kGE/uHrWqnj0rbDYGMy
08BeJwJKYvgGNVFmoQWQAsOhQQ3588znL382jm3fks7uog9oo+Iqe51Hb+hfDmm1Ikxz1jw65UBu
Rsfq9kAJkbN7dLme1LN/lvn7jj+fFzhpNNzA6hTZcckIYD3gCzxYAS1qXqno9eb0U7PjIxp93LAK
ZMGtGx5VJvzbgUqbeuTKP6O+oIl4TFDU/qrxDYJOvsQnzyrdvwnzRBIcTGdB8zz8yhgd+MPTAsMW
LP0G2/iof8aoYWdIol/IOrk4yPaTSPzAvnOhHbL3g3gfQlHxSDvdUkkizJCSJvjK/lBUSPCANhU3
gwxP81aPCLDybyBl7BS76K+uMFXMkLqcG7ADqfxs5WMr2C3ZEuT3xTu6lvMMHXUUS2bZogrFTB7z
cy5XoQaEkXNPfgBnvXBQH1MnoUz1gbKqu3Jb5d05W+zcTaabGDIzse/trwVExqJPX5IDLjWer4g6
w9ek/bBX72vUu9HHmK73A+xQQF1vqtjowKoyppsy8REoklBqGotdGjLMxTT6BazAOo9Oh84GLhzk
yeK6dVPvpa1K6hsVtPLEI9dcBBbffG5t9e4H1ecL5s8mzd7nx/drUuTNN7oUEV40WNeblVF0T0ok
qZsfPg/VpTy+iYN5VwHotW0VZAQ1LWwc0Gsuk2oZW8xGwdkC/rz873HCZZyO5XwR6fRwwYmmf2lT
WdVuDiehXndmryYtKzlMuUQ1lq6JmdS94nZKnHfL9bwdOtLyLtHv5Yzb5vWDkP5ovMwB4WFv8K7r
+Hjgl32k/PFXUmKEX4Rh3Iw5eOdmuZT3iOP52jdo+C0Z7fUP4b5m0G84YFd+lWHBGqi+OS78ABlJ
cPhHRgWW4CRtqEOx8M2jCr0SIPT9PzvYhBqT/6wMC1xMOEu7Qp7vjY4xGe8Gi/6ir8ZGqfk5tuUP
FW+kf5qi9mZUz/5H83wC3v0Hath16PoW1VCoweCKI0QfRzON6d1YVSSkNmnMgdkhaaZcKfYRsN85
Nic8HGGXmh0GcPFO7XbfS+Gfn+bEP/+V1VnQdzbOb+g80g/Tvy4LUK3/WZ5z5CaPFQOwcJeDvALB
+XMGbX1WuHlT1Nw8sw5FI2zu4ESxudQLOwWigHYx6Ml7T+/ZAT4ce9fYdywLnIzUYgpJ6kEs0kal
erPEXPxl/Ov+QcCbilIM2E1SjTVcjqQUqiho2eES4YWXFpz/kqC6nX/HLmhTpnOs7UGN3p2/Yow4
GH9mwynbH76mZ387Z321BH3OeN2EuaZCpBSfG5q8d+DW7UKe411QznEg289ppkJbgSygPPf5HM/t
duN0rYQ2DyuyB09sR+BeDw5VO+oVUkE1OgTiB00cEBskEUISDLbnQK8842oc5YR1Xu92AiPRaN+6
cBTgHBw8Y59TA48jRn+rSPorbLhsHRYBk5aiK+523JZJndUQe3sa7ewjB1axRg+BHII5lCPBwaah
qEeJJisKa7FLBmrFo4iyUKKLepjf4B6W3CyzpqHpWaBZx/TAQk6aK4+8uJhMuMGCBZWR54Q/4bRc
IuFW0eNCuph/6fMMsyG8rO7iefa6a6Dyqet8GdbedzUP0aAmCeKApRMUWfe1Vvq+7T+YIpCmdmZc
BEfvosy4xwpGVpa1TVsTxznHa8pB0AV5sZUz+KsNzN3CqN9DiEURIPI0mWCj0QFUix1apbpPjm1I
tHkD35uk9+2vQ9BiUw9pjp6eQoZsWP0XUfFac5xHdORbSZCr5iwBFmyGoGuBhRC6+p6hYdfTnh+6
/T7Z11T5m19+7HWamurE1sFpGPh8a2O2PUl5TzjcLYPlGVwyZKBdD7Z+QCDNE+WXN59AC7S641iU
Rx0WLFfibVdMrs574Urc93lCAbibVIrAcJyo27sItrzyq+VVaeaFz7MkuWpMiO0UGdJ4TFMp47lz
YUQ3FW2usxCTq51eMP18Aru9N9iTvTGKnlqMRjQpXUIjTUuHXIKRrXsniwj+GCG7W5JaquCKOabB
jhi6ffuArmn4dY/bgv6q8bakmP/1Pk2LFEuvTmj7CkK89G5VlI/mn992el2EgHj723vt8grkD2wM
HuZ2t/QcujCr33YGM1uOj1RVLydK5AQi1ieArtV79FGKuX/9W+zkchsJsFZj/7rz74H3wKw7lmPm
GO9qAYj8U17TSObR/FFzYNTGOzzOD/zBh7S8UEkSOTSCthaNIH8RLRrIVows6aueRhGdIhOwxdH1
r4MrtOQGPU/gYAuw4umLiIeUqF699ri53SpiNapGh9EeXtq+T8Qmv/W/kFaVFYgOgnB6vd5gW8sz
iomtVThvrmI8qQif4h5ojarLhK9CVB91U2dft9eQ/xrcoP89vQUHJEUUyq3U5Yo9PySn+jZghgnj
N+MqdDIvhp3XFLtvVPHxSCyBGcCeqUxKtQI/8ofhc6Mwv6WVFqoKVDGu+JMhfC7sus6bA90KMtLT
IV4PuJ35sdpu0d0vTjVZN6BjzjubWgKwp0ZWamraLUVUr4F+2UKHw4ePO6lXK7qsBuQ/lAmPewah
0yD5++HREAF5Jsmaa2IEysggEnrWuKbXeaFVfz3OpBgK+GaIRocLPKzWyFkLkWXVF+K8kdCKkeG6
6nw4PU86vOP4QS1aGJsTKnpc56sLhDjmKGThjHa7Jdhx6XBCvQnqbEr6P+W2PYf1iHEzkZdjbOpS
WHeAmxGYBpn2Aye4ip/mIubgJYoB3SNFOw4SGni1cQ0RIyY1iDOY8yP/Z1rcvVffwoQxvoi8T5no
fk1lQ9GIOaFHU7VzidV3wnkhJimh3LNm8DHJIGbskMrJx4Wbq8gsGFF1VYGhBAYPR3iKi7NLhqsx
ONExrv/H1rcHDLCihGU+IshBnGp/sVXrcnR5WrqCBdk0gD9t8qo0rtxFNjZ5Wmn9m9I1PW14nnAj
v7Fv5jwS8U2hB3dfab9U7kwJiO3fwpHlZl1OX1LKQ5N1713sBmINcTbNeHsUQmbsbyft8dUEO9SG
G+/+zlPl+cL/xhxFGRonLmthhKVsLLj96hi2GifImT6Xh+3QO9EEKAUgZGlPYG0bL9V1YutTgbw4
9LGQ1k+EXUSmxrdGAupJA6nynLc5Jasc7nmbH9olbIK+Sk77PoSJYGuV8EH92o9tcX1nk5wNj8nQ
ZRkGFH4f5wB1WvRVV5CFqOgq13nRW/3tZ0H9bE3p5UsRq0wWHH32EP9DVziiLpdXGP1bK3hKCy9V
2FW9GPs+aTCmC1vg3OtgR8OvUTSibRvoDZluTt+ckQ/h8g04MXNKLn+VjWQ3JbOmnEskuM29B+ib
q2BV6kT1Fqc8dSpE0lnqZyyk7YjaK+C0kEmU11k8GqpABv/T/amVuCMKHNqpFAo+MMS2LaGvZjc1
pUzs086KbTf0emFqz21VAPdAhkCNgP+RzTZhJqJqzSd8rFI4hutHl4uZtqjCheEOUX9Zzsy9ax7d
4/vrzPxRdOO9iP2SNy2bHC6+udzS/VT/A2vXoqYDyNG/8/McN5l/78KUqwVQvmv1GbEnhwKzCqM0
+93LDzlzdastPo5XyxnYBnvehiKtgMHF/iVbO0q/jOrxy2vhKpKg7jeQC6/UwtNquIP+4N0HXlnN
9ls1AD2p+6SASsO+rU3+aCwskQ4etysSdzargwEvs206sVXtifyPuPtipDwJBe96QodSUxWRPnqM
9co9kiUO7AKqG+CyaCu83x4PK3h8yVT5aQAbe6OvRlcVW4O3zscrA5bDsfF1f4NrlErvQ1A5qPEL
aZSQl9aE6CCn+5n+jTIAmoYWGawVoo0q3aUzic8dGFwXbayin08O0qhVnQ1zmy7jRZRCBtskEWAb
BZophYoyQzOzG9+tTy+3zB3V5yIPyuhKpoXuVJo2ZfbaJZ/wk76dRX3EVDEqcTjNzml3Xi+0apOH
GSPBZHq2yYhhBosbxvAh2u+e+EZPbVSah6WEA/TKEVPtJgb994eKSAm/L8GA/ZrUYTZ8Z0ueXPzH
jOSm1e01CoNwEsXYfBsWyhNunG8gfJrFrFQcwctgFyjx/6Za5xAgEzsblwVmyeBHhUwZyDTCiyMD
KMVuFW2qlr1ZlulHkNsW2bg0chdmlP7CDFUViLS2bmAqNTDikkaxLeE/tiNbTi6jx0VfmSUIoTBx
J9hLxeVqQcBz9hlGYqXPGxqbg7/szcsFo+QUn8LpbNec8vWeiOtmlIjtrMPN8gILkR/WIXVsHJuS
xJqkZp/uew87ueoPhWWd9AILSvrGOXAkNhW6zvlac/fnawI6K0r1+w7sUJWcWJq/+g9/JSUpuPWJ
BkcQ4pJn9Fx60KSyTTCUYl6V0rfBDzuRvPpjzrx8MESXFhhB7hDpDB7XdsLlVj+8Sx501UvMHUm+
S26Ha0iqaHI0zc+sE2ksnhh5TbgirQGvWfaYb35Zxzk7ocEe9WsIVXSS/Y4AnUECaG6AnHMZh7WL
HdHzR2fi3D/Ujcpo5zz3Gh+Gpk8N9mVukGzz0lKscAANR24wdZnXaPUJ0XxVyplGJMyMSl8p0mPp
JfBAI69l1DLJ3zun/1/f0+cjtbvLB8Z/jPUlBG1yACiPmZNoH15GGjVq8TRo+VDLSPnNjOWdAkBg
QH2sWvKu/c6lA0hXUJNrTvUdHy3O/cigSXHD+SzoOFTfQqVQ8xU+b7nkjz4xPXWChcQqTOYgELzq
3eEdo377qrMKS7zR5FNBNapZyUSTrcwmbeawcraOAWftndhkUz+iA9OtYqfMYxFjRMws1Q7/bd4b
xyGVPXXa3nA5/HmuzpDoxkW7xRhnMTMejTgKe+Q93lkGbErDr1MdBLVoxwNXxel4pljCNZvcFk64
GjNj8egnXsR0jlwB1JWKBKOAa8HBw+SuSIaU+7y/uHW+bAOSejrB8KGE+W3UVadoofqBN3rA+Yiw
fWLwawBlGseFTD0c4JcYEmCMRIdKswXsEgbYeGJzxkBx7QncFpZbx6eDlt8uLtWR7C5FjpiWSZ1n
NO8TegwXOlUETalIeXk5+EY7tdkC5b/Y2Hx7yUqKMKfStLSe71nOIzrYnqMGdH2RnJ9Xq8E9xPGn
P/9LWC4YBbIghnD2oiY88LXk0RCFiaoCjRCOqP/jqI+e379KdZe11xfphSU4hFak72yMNiCalWgT
gGghP8RLGYLLHCBnv7ZDgZPm0kJIdT5hfwR+uH65LI/N+F5YMaZSapAyMul6ZsYGrAZkYRLnjBCb
gnzAk+KpF4CuXBnaI9AJjJjk3TIRSWAk49eQYEKXN3zSwLash6Iaxdff6ku0nHdaK6U5IjOps+77
GB5n4W9rgjsZfXmiPTy5BbgWDlO4OUTWiLYUuGdF+80lNqWjN0h56O39r0L2cjNQ5ftom152mOs8
KG4C410y1pm4d4fWTUHaNXjdgHP8xLINPlkvvRq/QS00jAxrkwljGTmrVXBerUgYOEox93y1pxuQ
u+SznvEchjifPR0AaaWpIn772/3x6WCRPc0rBNKHSIJn9Ko1z+fzUdx/YbMabcj3O18z6ZaHaprJ
E7bktb9ps6vv64oj14ub9PsIL2jtxo6YToAZIr+xBjtvstuYDvG+7BqXViJA2nscUgh8C68XWemT
AA9+mIMKaljK/O1USuE1MJeAYdNe3MWJo7GGZxFJ1djGfcER9V9kAJmCm1OrR8X14Q/WpNnAWBvO
xTJo+dqRVN2m4rkyGJzIFUQA6pGbxuK2BVkX6ZmbDCJwYlrFrc09A7rU/EIyKTybdQq/NIzc+iVS
1mzrqgjy3bxpC7nmTV4mn+t/TeADZfkzgRsdwFnnRMYILLO0dhh4kwI2imDkAdEEg54QHlH+LAGx
CqUhQ85WpBE4LK03OUvY5Oxt668MWgSx490ww1i5wwZ+ANdy5f/e6YMFcXuF9sgrXqJ4rwFU8+Of
qo6eQfskfT84CCVB1XBc5Clok6DR/QEoJpE1GT8zXxEOmHNgyG9PRMmsF0/NvsZ01L2vWXMfkojQ
lqCBh6kPJA7+HnEaZ7LXAVif0at/4cVJFa14yQzITmw98DkfR464Slyo9l+mQJxapwvhPy6EJJ0R
ZVvV5BP/GgA9q83PZzVBekazmRRqMdB9fOFNz5hN6fzpc1shmHGm3FsfPPirWBTTdMD89ePPsaVt
hfQWI9BlcjtdgEfkPhOWxhfiuzOkwDCyl9t5nNv17kFfbzSnJXZCqtIsweWLXxB/zf83/2HzMnmf
gfNX+I99cQs5fHqnttbzpuAI+O9TAI+k+GGPw31zCRQv8LV73tbq3iiinbT79ecaVTHpgmvKKTgF
8ifvTUVb8eiOYuXsfUslnmL+WpjRVtHCDOCtRgDxbFnYOSeZEkv7zAnCawHz1sc4nAd8dRVuuZkp
Vh5CWyvI7exkGO6HIjfYAC/VLh6q7KkXcbxYHkvOsHpVVQKlO5jjadMdxtspZPuHHQyOO5aXAGKq
yVk+Tvqa8Tgq69BikGTO59OKJPJLG8P4pSI4DshtevujuXEoNd9S4XdINPRhpUZD/Yn1bQXp1p+s
0PfhgBuej5Jp+OqYx1o+7RAzBTLdlU3w7tPdfo0a8SwWJsc1dyikEpDgiAiKXsaeK4v2x1P0Nayw
3uI/d7K6jnbA1OXTbiiWQeu0hCCP45uxsbpoGSoEkisP3gZsqm/JgCOvdA0OxdyRrSilCS20CrLo
qNiqKs9nM5vTDXhSkruM0hV7PqUHDXj4UnadqIaod6E5TOue0EzF1/v+iXwnVrWDWKwmQI0d+pEC
OUfu/bGV9DPhMkcG+yP7ILITY4QdMeM4H9r++qOQgTT87I2WnAFEYbKVzdkQXB6/Omr+s6zsqQHk
UQSNRAH/01xWG8rJ270TckU9dEH9XBAUvQmYVp8ya7VJEmMISqpHc/u36J8Fwf2QNVyPIuYqalx6
ps9k9cBGoccb97SlHjY8uZ1u0vbMKIwIguggx9X6cv5QuzEqGG2r02zcGOH629SS+Ey24xfCezxB
LNqTSE+26Z7R+6Rerhib1KMIPZXGIPigURXfYga+NqbepvW3UImRYB+hHR/NXu9F6pOQmcStpksj
xIAk2UGpzPS/ceD9nNhwG+NXMFqtuY6bNIjaKMfzuN7T1uejA1peAHTAA6lcDNXH6r2sLtz3WBGx
9BMSnNjQ3OrtHy+BsCXwsHhd6joxoood/6NAoGmkfW+SlehFVRQStERpza+5/a/hFc9WRqctUxQJ
DIn9FRkcd0jKT5lCKyudVR9RS/6cmHynKEhabIMwpiZHK9F87C0N8ibhZxfRxkzJ/5Z0kTu7Q98D
O7ayAbV0BJG8XSr5OcpuRfrZeuRaNgiFAShvbSxSDQVLZa9SwRILatTKP4fdpyfTH7jhCs2NBcfQ
BGhnNw2KwAoo5NBolQabXiN2W2E9g1Gie4iuQ4eHu/XYDyZFOKlSav97WWhZyvRiGN/n6DczIqKZ
apJqkoB4ASHYIxTY70BdkValx+DIvfU3ArgGtGDXryKfW2ka8XX2khHhjzVO5bM8ciCmDbuNaAlr
p97akpY7ExsZf1CK9XsR9rDa6NUu/V72A/s9OA0Lu1j1/e0hCNCSMKvSJx/2MChmdbDx6O6JMz7i
CjYo3GUe0M2AKTfu2nMaL52z5pTlZrZ5/25VF2Uqo6FVW8G7O8Fu9TAu08bNfPOW1hnsgJKSeyMM
6xymnXUYsRkhyVtkTjdydHbYQuMfMdXWSRjcswNwmJVGIiF0y8LCoQu9TRXDo0tbVjUBNZ7CJl+0
ZjesSwCy/yh8gqqx+LVkVMRBjhXvJtFOpUrurzltSUf1CKzBtytneJWZ/gmZoCtxZPJ9jzIAQjyZ
ZsHdG/gRTnvbrpeuMUD2wFfZ0PZp89jVezPC3k5DdC5mnrPfpa6p46+UpvdA4p1empW514/RRuz+
KZ0fQI93Ny5ZfLE9suSvgM6acBX2grlMhPGmbCsm3cPR8XUUcE0TVRFwwqJ1d8prl/w/ofjG5RKt
2IVh56F6QcbnhCcf3MfV0XFQg2F/VXzGmCiRaorZatsvi0VZSj04i6tb7aqw4VxnQgX2iQJPBrRK
UI/aaG+QYoFI3AHFJ1zhuPsogCoZ+A3wt2drZRgmIYIiN2aA3HJa8962EslJHYe7Po9qfDgPx2fe
j1T4F8yBZ1KgytRa6CEgrqKNf3E7L761hgi2zcr1PRhqV+HrbAJCXX3Dje721ChDtopHTBwagCRN
Ygr9ycmHM11rg1awDa0edTuOMStlFrPT7w9nd1gCI1E17OYbN0e0Ah8UDYRS3XHrVk5SNFATUBYl
60XjObsB4NIx5m0HyKz38y3+Yts2gr3w7ifzItgneRiYuFx9F41MBt+D5CTkFeNa5Zyb8JJxCW7C
sP/QjoHOIkqmykw6pAjQBDF+S8LqMHIxjH+E0wMlpkuuel1Q5Wb8E94J2/25e7UUBCBJBgR85gos
SYqYwcud/xK/OOzN73sb1bSd1TQJ6rS7mKwLdng2WLp8+y4FCZIcQosfIXz8HbD2nGpejfcZjF8H
fIUZZ48UQEJQoI9K8DzCCmzNX+m4JIAQH/9WIgewJrE+P9mRJtFIyWqmqqb70MVw+zH4jA57tF0j
OOUVK/ePWmkcph6cmPJMmw4Vnn4rQ+9/dNdnq/O0jA7Tlk/kQbwu5/557r5rBLIimM5fYMgjRpx6
uzkxNuZ/HHiKCZtaVFCKOrnnlayGNc2JInoMou9EAPog4F+JT2ARed/K3O7vmAI2DkzOaT6gV07S
V/M8Mdom1c5HdUXuWvVnj0LEGAJ+mVa1SefH5PnUL9JhZkZKVBwXPD83IBv1/l+NT6hlRC8u1rcn
qfczKKe1aagyqgu/vtmZsfziZYmgxms+QvZSoM9Xt4WwfGoeKAgdMgbzlGfqhWW/gwh0GZN/q0UU
aD57ZyMjmXn4zCXJzoqSV57YAUjoBCixv974nT1MMuQJ8F92hAP5AxZezjLM6RE54wP6wMvsQpOQ
Siqfqz78xyFhfB/+X6qb6DJY1GMQL8Qxbz6nBmigSfRFJB+0P1XtaEDC+sxle3xNTSSrX3HPT+rp
5bljWA2DuhKxfJNCCMfAWxGNqcdngixmLt6ASVvwuV+jInYHsUuJXG1KFQDGqdMSHIJ9tBZQVaVu
1syzrxosQWv3UlfeQLY+eii/mkDiDEzXbp9n00ly+Yp7ooEyFveAhaRRV2iNY1h1lxC3kTj4FVWH
+Ov2pSi2lBHSYAt7aRQyTSJ0wdNqCUO8Q6R64rDQ0zyF4LQ040Y1Nf9poc7dUfGGC0tjzu/sy60E
9IMqqhZ34AFYUeKsbQtQNYehJK+jkY5moXwR2AcV5BaOrltBfcafWVJtiSCh7PAkBlYa3ncnq2tu
/JekTdz/Rm6dpPmd8jKzhh0+DPR+I2YNTLOGBl7zLlVVHMnosfE4bzmtk9zWxvqKGMVPzpL7OLsQ
dsII8gaFTC1mH5/L4TE9asyq/LaUh49lw7dj7fdcL5LMe9+kRmIt+s4oRiImtsAwO0Z9h2ePYa71
VOlMw0g/heISxhqRqo11AAW4pUo1Yh7Dua+iAhxWfcsYE5IPjhedN5aVR7lGoMt9tbHVzoQ2arM6
MFm4tPs6jMnNfLJ84DxlZesgvBQ5zwzzHk0RNhOCGDgjKsKZeaMdjXMGaJUElwpS6Unm0TjatjI4
7fP7/0ZntBhPK3Yx6GbvqmNJjqlZl886HN3zSWIGQ10zzoHJcw+Pw6M7mDE39nX0dSiEdRYZ3Nd3
jCD6WcvpIypL7OvPhbbVmm1dRBRpytOT0O0ci7+FovXDbFHMIh4dWZKr3zfoZl7Eis7jTIdOdkFO
LKfyd4nKBfRASSLyp8jUNi3gfnLTARAO6GUoKuiL4CekUq+oYaKsUy/w4LM7rsBEzApQXCLuxo5d
+neEm3I+GnYbbGpWeJ4mqFtDCAZg01YhAbE2Ptv4S7nLPyxjHCbXHUtWy3iyZNPVtIT+4+RS8C/d
Pt+KH5al/zYJaaBYQ4T1QCRZqwplUpd01eY5pYBdvoPO8gNf+q37pM4Y2hTGVzsCGM1w6oIu0h7J
Vi93MDAPaUrMQsqgcvOuiI92XuHdJyNUO4LZYnbKd3P1feDoHFtJ40DwDi4I98uVCR/5ZaOZBg1A
Crr+WPewtHjMe5Hf96uAV9OtdZy3hkT9Kl/YHCJDyInYnTx9kaFKpbTSTOFT4J7pT70er/5fF8nI
wVGHg1mv+I0aNtwAcpT54WpUVHJNJctjRA6f1dFffO1V/mpxvUE2x66/mvkDCvkrTYemN/mIGaUm
ux2Z0/szaOq5yJR8gphGr65D7ZD0ymaCuL1X/wT0vepDvKuFxv/zSduUN1MhZ+CI+/trWk7doqW3
BGAOIT7btcuKDxu9rou9jvZrGXiF7Kcp3swgO06e+vKUaav9xyXaKHIErQ+eW4JpPGVngzH6JGZN
8IBBJquPhe3hK7sNEB0l1UFc7g1PPzHb+FzSGrI0tYIPVZ3E4URW1yZtBz2T9tP6dljjWGouXhFP
8W0HDO6cJFTZehtXPzzqKKRKcE+S9+5w6zeGNBo6/ek+wlGvYyB2X/bK/hCg+05kSqBt1Nu9Ngp4
BHKuVmBTDHbbdgiQ/gGFgRH2nuCpVoRPhpaWrA6TUaXQqWCR78frljt3pi+ALqfMTRWlH1WPwsBu
QN7A7ZmRIIUmb/JCXVTV0IIwGgy3460B9CtBMXmk++9q/9TUOsjPS/KbISAXe+R0dEOgP4YWLIiq
tLnObZgBwqlXtaetNGdhhiYy4Z20N5EbixuQ87pfB+j1YwXLeHIRRLEAU3EMcGT1P8BY6eS4nIhR
R1y80kE2F8KY1AcknPF8SD6wHr8BOUvAySOboJ/k19WNoOlX9h0bfaezUxA9j1j7ulAPRYokCfF9
c7/GnjDnIrjjJiTVBX7VQa0OPiLeBRiPQGBlHyDEdvfCJXw4mmE0Td5jl4E8PV6qbcTI7iRKexek
7OgJbJDOK8yVBSRZUgu0P2eYoHdNEpvZQEn2AIgtK09WV/aE2ahSYvtO1jzm5QcsD+KEMSzkdYr/
aviQNrS1YCW5RZbAO4aC/0NFUBoEq5JnjUPxAWCI1T4c86ZfTmxDfwv0iPTMNQXKtMYhWbdzrTe7
KPRXY0xKXQQmJ1/rZKwg/WfTZvC3Z4IKxan8psn6NiuyfDBo+B91wb9lKRI36jOTW5FevxyzyZL4
Ra5tyc9SaKCkae9EPnXvqRGv9aMsFnCyqQAlQQTHp6Tsj2NTmojOmvMdfN4qtzIpotq0ND5o72aG
kRx2jAev+AQa2AGgWQy5c6vDYqQQNHZOsML0SmukDTMGXCZ41zOQu4n9sTGc8C2AehWb7/QH70ZR
jSk/S2K630CarkGtLbX8sWo0VrZ0I4SVckZuBeo/e3TCno9AjL1+l1s6C9qoplbwyoEdUmO4Ka1B
vxz1cM5Rq5/e/qr9GqFqKzS17ptCVxfKhbIhEG+3l1trOx33aC02utWxHbAb7lO1dS8HPP5h5OFG
ay0drZzusF70OYF773aJCzoEgmGVWU4NUVdAsJL/hrhz6FtaEeXKoPeimXsBFqR5qwrgIr24uBQV
CnCuj4VZzGvEwnT9QBRbhpSfZCe4hG/+2TO3BN/d7BlO8Bm2RdtqoJ7/2/6tUqIfnu0DEC9qb40F
ZPpWIWv41bu3Q4InJdCo7jhQJQxrEOGrsdlMcK7smDjUfQyvjs0A+0kmMjr0Y5NrIu2Cmo3fDdCU
vqWK4Cz+qptnEg7NHiMgdT7EcLBeQ1Ex37FDKrTJGNRFPEByqi4nrDa3G7R9twc9ICS10238csnZ
lGUaxESnbP4H9R3Yf5ifshitL7gd5HrfJGE1I5x+yuh6IXjmSQBzAidBfIz6M89qiu9UV2nCZwj1
aWQYxi9b6bhl8gqFgmI1clSasaIZNlvB/7WUEnogr7adUxRXP3Ee5aYQdNvXGQzGHTOVSpd1hsLB
06TZIZRgFNZe7xa/o1oNY4h30mUpdAydPUpQKmJJMNoKYCb4+Mnug+40PGFTJEwuD39XxHvtIMN5
32ZALG8ElTiFn5cWVUA7foK+FwurBLmM4Jf/Acoj96GN+5URtqjcXNUQfkM1JHEhXyuK/ab/DjOf
s1+BLM+1FH5u0XBT7KBoKK2c7AB+Z9O4849/PVLHFb85jnWp55eobvmrMKNnkuukyH/zzYxLMIeP
6ZhAvY4/JaLpVaPSMV5XJQ5IbArGhbJtFa7TkPgexmc5zJd7UrRSjX4r6VzZ4wiypa2UCeLmSZkN
AeYdhqFBx44eOcaBG61Qeo3HIwwOkyWo9WWqzcOrELKxhjvvwqlhznOfS5tlocbnEdIm73pu3M4z
mgXKuNBkszsHyuDsSrb6rQ6nYG5OQLCGs3DT87N0wgln5uGCxZpEKCdiEWV3xOBR85QpesiqM3f+
E1/JxrlMf80fmUHKLw10J+f1thsg3Fl7uxo9p6thpxr3eTZaUwzTX8iEe6ddCDsP+yI4sQMNUonO
mvHFRUSneuJNjncOGzsysf4YZ0s2GPJlaFD/QkM2Dh0BOTHBeczlFflUdAhT5c9AHrqug2WZF/us
jp1Vf67Ci5cudkIWCjIBwFf+MDQUUfLfhyJ87cYo0FzhYc/bd0Bg2nGKNU8AtlDrio/ggP2ieJhF
D7SwLfAJF4yriMbBYd6ejBl7ZhYs5WbD9SUeCCuUGR5WhP+aABsmwjtBb0KEG8Xq931wx1dSls85
9Hc7BkXcR5B33mJVzIknt4YgIanybL+xx3Hg9p2SkTi0su3NWeacHOUe4N2vAenEvcuVHiQlthLL
Azj84jhekYRrXx4HUYFiNW0wHihKv6gSdbWe9srjM+kVLxwbzlnHdhJEXrhwwoXLWUQp348pwnQX
jg0QTrYKzCsIGvgK44gao/AuDq0Y2Ti2gfejYc948wFC9OMDZeS4bYQsGLzmOH/c+/dYUUOP9zqj
+WTuSUEeEG33GSiXl2j/IhZaelqjt0UAxIMor8fYnKTFYlW+YBa3XYjjV51icV0lyZBDIzv5CGBe
sBLKXeB+fVlwU3VPpiEoj/uuCu5fzGP6IInNXffGwiK3Pv/hWk5PEuEbiOUXSWyoi6DMRZzSrLF0
bQWG4NvYCGOPiGEdK99ZGrAuW409SS/2ruxrpRMAT9X6qaof4bRXAKFpwUtbC8SJhrAX0qt3uQ9m
V4/il9ZBI5wnRAuGfyAKMorwOW16ndPya8mBbHlRbFQwneNaKCwUk8qhVZXFoBGEfGcbjfb0fg/X
xD64bKx7KUP853KXBBvh0fLvzZn0Evhd0FDQyF8saYmvBmzaTMRifr4zBH0fQ/AwmqhKi4lT6hAS
vtbfzCpJBpqgAYbuOBCN8VJsJTIazFXgZK0kuKTUm+tWCYWbJJm13N6lccF0Rv3s83rsNnA/YE/F
sX7rzXzA5Kaunge47bt6hDVaxcx9b3PmAnV2cX6JvSRj61tsZ1qEV4qWak+n65kuzqtsmmCTAa8p
EDN10bKu47iVhs4nHfOrKnualKFCDOVdtG65Hk66YIJ9wy61v/3wClyJ2oKQ3fKPyss+t/1sB23o
shRVTHUpSWNRKkgRtGHiXxE1koCq+BjzmaYo3LRTf8+ry/BbXElZouhGdyaIst6Fih1N8Vp73Cdk
WVPb3kJfObFauP+KcEAbBn/EBwZs8JGhfTUm68tCUMLD2MJu+NuxRYU9O41dSOaEiNWVr11s4r9q
yprYK2CQ8la+snlUyKrwWP0Gst+58Fd5CbJja8h5IWwWI1eDdEl4b4kIutlZwQhuWtypz77TPkrP
s6Pb/i+1DGEtYpfbA8070p1dM5DJyYaFpMEU5oFk3N+Taf6SEtUTaZZp10oTIXQH6xu4PeLqHpz9
EE/nQh5hUuKqbG++b4cDa0CmU8uV8JTxDZmOfn6DkOhD3bcXRh9CFeuvyuhj8NkwXYJRd+EQXpk9
nqfwkWryXyDGzkKrEE/q4qB7jlH1xp4bnZOxldozW2rzjkiDJ0HDL5ehfkavXry3gwsItzh0sKY0
DUHW3Sz21d/dOJnJba8Kb02YCnEnJ3zw/8hB2ehXzl8sP68gTMtXF92aouujq2alftngYIyrx3x1
/bd4G3XOTIV9R+VEGbd3bLcAZ05IkNY0oQ1sZuMMOAbsJehOujg7S0SQsjOotIcVvuBO3BC8lGES
JTWn+kQ+51RBljI89ry2pAGUPBSgKo8/BX0xFI4tKyo6rVsB4Y2hGkBtHKl+DZtlVar+KKSJvY6Y
SU08gYpHiBlYwuYUXMCD71TJ1LlOe1ROB4my5Ru4+idzYmwzYDze1420zLs2Oiq24vsPP/EEfeog
kzoDj7IxvDWVjNgHCWaYYW3o3FT9n/wHJ56Ex6/u0HSnfUBcusUsV/7VIZiFpGWIxa6vwGLJk53u
BCHusi7F+NOeTddwHQFRilzK9SdwuSxR2obtgztXnRErUXJKfUJj2h4Fhp5cITlL64FgaeQTRW60
4IJ+u2oR6n0rSaoExsUmRVeiQKfbxyt3bHRzAyD/FQJykmyxOiWoIqAfV7m1AzhHzaiWKOTMv1oE
4vGVey0+UpeRSU3SqBtQ+16IIIctPhBvgsV4mjnxn8X1FyhSD54DW6M0jJ/uEhAJzo7A//81+qzV
a+YJR5IX4awSd0qFNHYlSaKUt40sJM3qDSUGaOf9G1m0rQcgXYb3TLk1kIKJjgF8W2q8n6xK3FX+
HDWrfq2aH5C1Q92skYNODAeQmdjRsWcG5dCa+OFp/i6YsLnb/aNlxm/96kmppJjhTyW89UmcW+AW
SN25X4DMsxXmThwL202qCc+KRVsNDLui0lYDhTLxfhgxCSSjuW9ra6jUTmOx7jjfLVgITialeLh+
nIR9p0RuGGC2FTL8rrtvUyiLKbnYVtLGs85RG1lHP6bbkISc/aD1vthY7FIluA2x3SSXnsbztf5P
YpPnCqvAgAO7+taTrsTdtlUpXx5Z7y8t5CB86HDBkIM489N+J5yB+r4wR75qRLvfLASMBNgzoxff
DRVsKHmBlU2dgRpzo0cP3RJsUajGknlG1Ha/AukU+OEjbuwwGv9O08sdZL0bCUrsMLXK0HJTxDiJ
HOVH+eTnWaEd+xJP9Ghj1B2EWDQmK0H1i2fhvSx0O6MWzrjOvcabe82+Y8B4TCk2+7FHUJQRKuEb
+ynp1koJCJZ563ETHPvZ8xKG37S7eACamjWxnAFWDzSUoZxfKxt59bIa4V+apDPXzahT/htzlXQ2
XtmD2doniAehcT7pHviSi7S1zABOFRJnCetIoGkP0suuBqpcO2wpqF2CUOFAMB0ijkVW/xdl7zMk
oZvV0xqFtVoV4yqPdrGcdd9SemG/Hq8JyW6T7kD3JZ/MtUcm2grQ0tJqA21cjcOv8kNDZiS4TrnP
orWqSJCHh9ePYObsjYRGsaMggK02DLOHVKJxw69EVtZqqCRBIUdBt87YA6j6YJqFgSkkw1Hov/l2
gdQY89Z4uTqh6ftO+lcSS5KqEOdLVqQl+dwVXmMcGNjer/hC+wLQaQse82ePAxF7QcO7G7M1njTh
EIS6kOd27lxnB+nnBLYR/T0rnAL6MRo/R1X/hT/RZeRluHynKpS/tDRIfyAqGImbgQ3Bp6hxuQec
Ncy9AHeM99F3m6xvnhvSxS1b/GTn8OsukDQUB8DqhhjRBfJ4K+pXS1P/l8RRq3aKSPnXK/Ec3Vus
yK1EwwCquchCJTEqoU9C7eZ+wYZFMHwPmStKPJYwT/Qg2rkdocAFjwV4Q0TIZ1/VAoydNLwiMYWZ
GsxP08+mNYk2QYk4CVEM59WgbC1p7oK66jeXdXsxs384mVE78rSqwTrCwdHdJd51B4NwWNeQGhUG
KR/4/q8COS674QYpStnD1CAJdOwcpRUF3yFUl6OeKotG58aWtZ918mGpDtggS5Ft51oPWuwxQdnU
Sfwc09dJxlpiHzr9AhsOU9DGzqtxhlgeAd+spL8wIL7kUluTyzOQ9OzOAsjt/+uzlSY/7t0llCNY
eoKtRwlHyfNp3jbMhOyO9qOC7scLfYqi8pOUbfR+a5nyNp0kWuQiZTRC0iRHogPa5qsIig1XftJl
gMZduIbu+nh9hvIPc148nUt9tdjrxfILTq2FfpMZsXHs5VaQxy3Z5Eu5HjftRo6dUfLjzpsRSPQB
Rui4hHQUuzZaTgUY/eU326Cnr3M617HCmZbKspTAQa55zARNRhvAyOrC+XdMTBrY3S424Uhxn2yB
pkg4JKbT0HBvkfp4TcQ31np2BngeQf33CPxTpnmB2bPJiM3GfFqc3nXHDi55ZGTimU1onqVLnfcY
tJ7XX/cWVsMFDrCL69hYWNK9rKBtHXJnQxw9RzJ6jWGENpJ3EKj61q5xd/madZgR4OWTSXoJtMq4
9KbQ+3tGOHGudDwmnqS7NQ0iYat+OBQeo5WEmMtYnoMqA3lyJNOR3xCuMBS55iCV1VZGE3gZdH8u
9oowxfjwbYPA+Yaxfv1pk0w2+GM7csZVc/1+vIC31zT4DoP8E5GUoGSF9nnHt5c9xv52vBKtcAV3
v+rmuQZ+fiCvycdOT82z8+N+gX1zZyWpoTJ9zw94DD1tFcfu+GuSUhihWngw3GScbDM84EFRzVsc
ju9cF4ZUTAGfOn47hBVcRlgsPiKP/V0baWeqDgwMpzninX6zDkXiWzNl+IEcBSaUt13V9NTuk0O9
KEKAWJoL7079o2f7fiQgIF/C+K1z0qXU5he20XnYJGNsFQhp8MCILqxRYp01Ye1sOU11gd3CRtq8
rSPeb/l3p/64uf0iRsgbPe/Wkk48grZ5T1hTjfZh8xVjtfHHBaPWthcZSrrCCIthIQqjcJEmjU5l
c3cogYuMKOYIo+hEe85+9+O1Yy4EJg7ofmZegShlby9OamXNiwqCYWDjh09w7sU4w2pIpJmB9H4K
LHes7QJbAkPJuakBcWQT/vmdBpIvkO1hHvmg/AMRptdmS/N+5KIZsIjuoZOP1Vslnjwf4R7m7Jhc
De8IyCG4kfzW2xQOj0vW7uSHbTI5qftJAxTtN6Hv2a/9pQ5snNTWVAIPzjud4SrfX4fEROluOIwh
PwH8wKI/jpfp4/9uSRaqslwycSbdnCLoA7dPQkqAVJkcV0for8tm997Jt1IQDjOP5JEHl35uRBjo
3iD0VcILrS5BjL0EPWurGyMGMEBnPevUlduwee1G+EVNjz0PSXP6N+UeRHVBoQorm4ZBEm7xdgSC
WtLCPfRX7yBfyq3M9cFI6zRtAISKxu6fikk/q8fS8OJpLPVW00aXIP/FJ0+DfXu3zT5UBQsbzrew
MljMlAzT5pZh09YftAeZSNDuBCxEMxG+0ePlfAFRvgoHnA+cmWCVBajwlIkfl1gl2X1opaBr23gm
tQMidl7q/XKllAtplMkZOjiqKUF2kxLwRbXfUS4fWxzc5Z0gyTXlooU3sfpLPU7/unL1j6v8MNY8
MWKBuXIumJWz1BcKeAfyZOPHaUJbPjrOpv2S4Z9c3BZO2++Psu4ZJbrhmNQvHVPbC9D1O7UVnqFz
PiKW/mbGZEftE1iyHXrnocdDdR+Jyl6jyoneSl6LOyruRV95n1XaduZEHwJWEVR/Od/0VEf7Ahx7
8eC7oBjcOFH+eK0eNnDkjrU1i016H+BTq3VmLlqTTa5AEM7UCjWlWSl1717/Ksq7GkksFviKPP3x
GJW/iUpDN5yXqirm8eZTGoTZ+rELMWPGUZsXObYlHjswrTA16P2lGgm20C1GvKHFNXeEvRNV6C1Y
xsQjPBLo03fo3Wer0zpenTmbqjR+pGlMFFTzGZEfuDi5RXXanSn1yC9vKEf+2pO5MwZrXCSzu8mU
hIOd94YaVzu4yLVclSMFyntvlq4c9nBXWW67Eldk0x3ltJD+MLCzis/np/n1f00faHaGCZXnqSZc
KM/GG/6Coy4a/KQJZGLG1SyajthQ/DSL4+VVHFuhbeq+oic6eGhCTmn+xwfIVo7nD1/rXbndnn4A
jIKzMR1BDwKwxucHN8L8g//1Wk8nw/KbLucN8CcTFtt0PfuoARJmhEoorpo1vqbaYBh29I3q6DX0
+Um1pvRXG4hTpI4Vb7giwqi/ZcBbHMnDZUJAYH66zNZV2NDo6+HJhDKJJQqYj94QrCp3aii9gObS
DHqvNLt/Rkb+to6vh8LXJg66xXVHUajg85DETGbEbWn8uXCKnM70gucicozrkPhFXsxZD/4qc1rj
p8uEpe0EIqvs4pk8QSzq909OXN5XNi0D4Jjpxk8ijjc+vqUgZkw0d4s1fcutXBphTiapXQFNwsmG
R5jYeM815P9aMErVYOyzkY7vCYBW2Wa2FsJP9bazxlylwRlwswWybAmnkedit7YWR9G0jBXOkgCp
0RXD+3f/p+eF/wlwjCkHP8OJcQDZvHNJKfrzOA1JboW2bjMRFRlohHzD8yvPpLoZ2rVR0bd1iiR5
miHqgnCKbR3PRE6a7kAPmCw/Ll7ofDv0reNhywB+NVPG14oNMjQ10SFcgiJ0fcAIHb2cUKLodIVp
ylOkuVHMcvQSLROfc0b08KXrYmOiyEa8UmUnvcdHqxkNfED+oLcRsd32SnPMbxgqSl3nqWHSs+RY
mMCz/+yCzm7XTbo+n3FhK7S+7+9cJQgXSCjmzSRnSGGAvSpLUAQ6Wo94RqXkgDIlNILYVO768Lns
a/GfGW1notULTyNIO01OIFRUm0xxXhqvsECwV2I93QuRV8dJf+bX/twrip20sV2v1ki1bzlwZm/X
EgEKo9Xi/zf8T4RK6m8YSkW1HvJXfkAx0x0AzDmmsA75nfoR5L7UnbdwhTIxeu7ZRDAzjovQgNB1
jF+4jzt0A6MMoyHIXBTeUJWvYH+YU7YRnXvoLd2Qp+YOD5IOUNsBGBtYJuHnfzq/ohpHRrhHbFhj
A3QpEpEo7HNElqpRzukfdETMJ8rVtVLUrzwtImJA4orHNJiXgaojy+5uo03Hj9jSBHjZzm4y+aVe
j+vg+DV/R1SK/1xWty94JAvva16I5m+G8NmPHoh00mKrv92NqL64YctK8EgUeeFAsSVDhHE1var4
3t4J+ufWtK5lKvIxTrdTdp27q5FdrMIO3iGLC1wNhnC9BgxnZ7yFursW3rR+mYbqaz6plaqahjyY
NCuy2GXgADb8djFhaqaviNt/xwjNnorrN7hR+e/2x/ZSq535Ugh0fj5js6UM54Plbcjn6AZ24Wou
JczG6AvLArh4Ym/Dygv3+pCwNDz1gYzvqD1DwyXxKmYmJaVG2C8RBYtAcnE9+Y7yOx8jAx06Gzbs
tg00y0yu+LEr/WAY+RcsOqYkBpm54orSE7G2pSmm/k8HV/1XBC4wQDeC1dBvGgJIzWZGuGKMQv54
LVCrlQzCegV3NDK+nSklsSajD5/90K5lPblbsSJwCrjvfzpHK5pND47J8WAwI1NhbIF/aIdTAC7L
lIINPvW1Wr/8f+IXMu7e62I9g/vWo6kwgGXFC4AUWHnTtqu2BApOdjoL3NAa0Pe3RkR2elA6Z9yZ
9PUtCSCOZ1S15kN5oc5MscwxpKbf0RXMYC5lwHnNDsNFDeiV4gCl6JqF9Io3ZcqLst5SCAs6jyUu
ny3R6n+fZfHNNXsU96lxH2bpNrBWd6/N9iakMZ/aMtqEAuuCVf0UOTQJtIc2t0UOTPW1uKaBIFTy
x3jlRehHCDeNdDD/5vaI6NgHl6i3VrQsQp8n4rH3o0cMkUp19wwqhuPTFcNlOr0mqZLM9+5S+XO7
JrP2+4D5yy/f2qYjWCpi1aJ8pZTr6piPmTJSmCsevayV/cLCEchKjMf9lu2/Y3Kt7m6xKVIZlgWH
hK+0H7+WDS5XuByIFxsqvuZQ4NUJkSWmgKqZJT65F1RIHvjbrWSFt3IlgPi/zOlAJE3lx8VjSDeN
aZ/DCxLMEuR38NVZceCzRVhn/dDDVMwoGwLQXTTToKgnueXBQVTNKTHcXccQd9MSW0byIFLfwTBG
bJ9mXa75RDpnGuAyGyOy0CkaZcx/knI2OIDE3WYdfsWxDhKj8oNTrGnoa5uTD2iNb3/FQEFVGtQt
426wG3JYZ/oe8+rbF3U27OB664TmeKGTh3il/W/jXMfs36pquQEYbH8Gfh9VduA4SRgrs4HPdMr7
8N4OqEYqEhUG3OF2wpZ2nBu3l3GABx9U+k+khNRvrj+55CEpIKkUZ3m7NtpbjlnQ8Jfad8JAzdZR
eJnZ6ZSSqRb8m73Bec6t77i8ZZ0yd9NbEKrfxwNkvo7613SSs8on6ObpQx9uWCPQV8YTT4mI6rgd
18INDu3DuqLE3802RM1IB5RwQzyu6dm4H0ChD22ozYhrVe4SOzn45e9bejLos79qA/01a10HxSvn
oz0jDR3VUXzLkJbr9e0mTnp/yNleBHHZBm564fEqi7K32TnhYJZGrvegsbmKOrbG5QF5nsTfkEiU
Oj37lscJpZJAw5q3aGe1gg22YhX84t2ie4nt2W01nVEACcxmte9bho853HedPBCfdl9hrlCSD2yJ
V20I47yIPIIPccOSyFSr/27lNJ05AiCmgS/m1l5ekzP/VUvHQLg7t7At3p8CZNZgaOVfsdAp3fiL
9tgZLmNqoxpiEswectUsPZ7ftCUi5h8poi1u01xfGy454jdvIt8vroQ0ljEzPAPCxL7x7+WNz4jR
DYoY0NVd2aWbIoH1YRdWihSlifCVK05aFOFc+EKfMU9N3eSDoWTEry85lVGuKHRn6asAz5hsC91t
mJYkoQ0k0MHAO3gjujQw+KdHsOyxnwR8ZaIadnSzJRcyCdaFAYlQ4E3QXRbeU1Nj7Hxw25Lq30/w
enRMuXODZrIJFXvHWsFrI5Fw28gDcx8C2fdgcRlALZPExs45GI55ZFL/TyLnxWD1T8pjIVAaGG97
hu25W53sE9XSK+qUGzGwYo0goYUuVpi0wcJ+IC16gr82uYiD1bXMxO5mSQUbvnkih1JC/1it4iQP
cb5ZugcBoZxGMZMtAeL7NnTWW4BI3wHLWJkwtdZJNlTEAqaW0G37/hZ0h3HLMbEptFkdAunmDYB9
jVSzmNY7sfWqVyebtN3cPW0nOkFb9RviI1aisGsUTGiQW5EMsFmXa5DuRTrkp/7dTfyJ7gedBhxg
UK0jyrI4vtsv/41lxkbOYwKnwFcyTtdlbET3ivZH4f6B8qSSVnluqZfRO1gg8NiLVJDN4nkf19Ks
FENVm/2Im8BdBPLIZrTK8KppOqz7ZJ4lGVpfuf5wuWGYWPxEaW45zsgf9XIwUMasdHsJxb/erDdS
xhLSCRsgpDaDrK3rhevrVyTRHt/MdTNcaLX1PvGqqgy6jnOsixIsPcIgGrQ6WUWSEY2SKuLqeRH5
mgO+4dryT//Hfn/rpnFx3+rxFWRsuoD5vCybvmsmB/Kw7JmrB6lzuBLDkUOtB7y3WzzGlYg+2ORf
zyX6Bjr6MUVuvNfUlVLV04LWK5Qp1wa0WjxnEcOoUea2fqhQX+kkXjcD97NY31/b1H8d0L/z9wJq
fG9kkbSi/jud8OBSGIGjD/oHPeCpAQvbwlxuQ0pu5EeNdT03UFx4sYI02PGebQKTozrodGyf9q0E
TA0s7Roq41kEe8Y9PaMZQA2KNknZ3mEXWrse7eMTb+39X5ABg0XiwrYI2wL2EHHWOGhBtSQypAQX
gIOVHDAaf5xDGkDONp2VsRQkssc81I/0diT2aSB2+K+EEDNuOGXAIKAV//2T5jJOuJZI0Z0VWlmg
BL/0rfJ+kaHikWXvK0yBEdGqhRvk4coiTDb6aCEmyTBshTzrJTmEXz+zNzc661GDlU5uIqZtbldl
XUmjK3k/mumXHSrceAnfkerfigHKmPqZ4tzFzeRt3WfMZ17fy1v2oPs9cCALCiwrCQkR4oGuRhwu
1k6rPdFA8r6V8Ot5cj2yTeVNHrJBkZ0Dso4o0KWPrWQNA7eEMaWytJz57OVE+QkdB2+ygf2i2DP2
dBSbNCOwN3qf4RtaMDVuSf3OZZoU8/mX9hGmU0JYRxzPCsxzHlD4Y1q2onyse9sbPqw9I87NuRGe
ktqPcSYOjfNz3dJKFv7mz7pv7dyu+J9ZAG6NUF0Bu60xXnqhywsgmWEXGo0oucYWe4YOwGKJKSkN
gDm1G9t1Ngdsp/oUXDAW0LZxnoRxh5LtnVkQsiAFFl0Moq3MWc+uIrjIgSil36XOOnaMjPBBrae3
CQ3h1DBu6K8HGnDxUwWiZj7u+vZu4n5HZ0v3BdLPmTOb5m7KzHq4oP7PNqKkjWBE0K0Gzs37R1AJ
/Af95hyiciyRLTzBmImi4ss+YQLVgUXxg/LtDbvnaYiG9ckZqFsUSuI4I/iX5ELBZ+irUTA2Ba4a
fq7U4h4p2CfYdPG3ZNVx34Ck+yLyHpASGrr7oHp46LQB71pwSjHlOChjemn9K44LyKte1E3tRzJf
Mk0xT2J2o2K5NHHKiCFdyFKTXfuFwGLYXZLxWI8xDGZr9ASL13K7ixWawJVmI+s+iP6supq/rjmz
MmtSjjfFQ96eQkdvbyYrPawMI10LlkW5G8+zxzXuSm8ujmuFiei/LPxWwa61z94a56JQaH4BnEer
svly3KnrAPrZpQQfFj/V55TmggxXeU58RHfIIUVXaVK6h2DX1Cfw9CNlYA3iOnhDeYwCMrFyhlHK
RKTwEZZaSg7QqZfTvagicxcOFwyUWPT6rQONlLvAuIRHZp6XxVuMA7wq/4v70KVXUfQYBEl3F8MS
oGRUUedDVLbeuVWlbSHgQa6lf+e5g/4A0vXLH5fbcI0fOdsdUfTZpd8b2LYTA9/jgYehCR0s1O+n
NM4A9ZVeXgdIaAHe/FacjL+KQeeyjksTTEEIlivkIgI6t7xGypjx8knihITmTZf1BZbCWV5l52rY
6xgKyOcMKFXmKbmC43czjpCm055cZIk3a1FyLIfLExUDXwcq8t4sPXKsBiYucAvQ4fXB38+wM0EG
Xqli2ycZuFU/QqrB9BtDs0OAyCgqTcy0txH8NAA+W81SySRRqLX+2AXng09bTfH0+TZzmGhBG0+S
tzgecYwGPofQfmIOtHTyAXPBDWm98AsFFQ8WTfTF1+M8HyGyUCivGOLIKTV9lr840/aFtNOTkt+y
TP0Nej9so+k+Xq1gmeDgWHbP+tPMXDSbCo9+GwJcr0V0JYlZQdI+kwMz6MIGNOnUjCse0ELIy0MR
eMRdh/MNurpaTapfBVyupSPZ0PRi4GUWf7BXhcy0mF8+iqVcNu4QqdCMTBKXp/+9a3bo1+zDz50Q
PZmUJFo7o+pNUwrNaSqWVMV7AQDnEp7XZju46aIsYw8Q8AvQDB5rBbpPBfQGFegcmHJf2T2vgisV
QkA1ctdhZe9KhXf8bVDtgGqnELlbcygBrSx9HtROyuqh4gUonGy/kj5/BVPZnduIdIf2+lVjp3/1
Q7z2Il0QleWInE3O37Rx2DB36SJ7XQUgk1d6IJEtUlZZx2WJibyP6ygOdIXT0KbaNAXOL62oMpzt
fsUmtj78KAUzqXZ3LG4JWEiiBIlobW2ynOzd0mZFYiwGa6Cn7PNo1D0XxGOjAws/e8SGr0tsJtzP
BDShWnrZqtWXzSacYfRoASVBPJR4CQgf0X0CLHfhQZJ2Ql+XiDeo3bPwKVHYf9gAo23y//3IWAmT
AFM377ibu6dfpjtD+CdQIRytuezEkOpJhi7XvCgl9p+8vVqEaS/phh9DTo9S/f3es3fepvqOaVCi
7s/m4Cf0V9A0rBTAxXY1nfeet5JYe43tNJHBQhLmsA6R4I5G4nx5DIZ0nh8Bf521HYAHoq0KxF0k
ypXM4DqSojykveZQmPAZWNt4v+auhoI9Bm9292Gu51sFDTEavvSYl4btZvEvhJuKPq2BIB8CL5DT
bkLvAQJhzesvYVFd4oxmUaW4UZVqfDnpk27qZ9Bvk9Ecq/93WXO0JdZK61/HD8ENWXWVE0wV16hH
77VtqPU6QeM4IusymNvAgq9a2mmsh2gskeciuwf1RZ1UfMu/ZLsIsSlv7hYekCX9D9SkLZl5bJh0
gHWQE941RsnNuUMv1jLlEkt+m1nKc37oVnYE00TVfxFP5ZJSNebMfF+1G0l2mhsHWGBVtX9y0HT0
c/S2AJYgqW6uAcaLuG4dFiaj8zFMEkMTcUCE1GGon2MPC+IexDYDVxZxJu8+7jeXlbBc/zZfhvh9
Cz1tbJLNzPm7mJ3n9Xq6BRtTuiKhufQ8xqI7iLcCfyzg92YVkM4W3EFpBS/59/qskVdkU9V+GU8Q
xFl8YYKxyPExBeKVEEK8o4XwVtsRNsA2Kpksxz8m9AYqXGYq4pgM4ZrsMgoy984MIKXj5xMvvN0T
nsyuATZ4ZmVGUlfyqpGuWcixdDh6nSkhtY8TA/sRJUhmZvff9TAQdXwPS/B58FDMa39FrNEmYPid
cTBBt/Oz+YS+6cZyIVPDeoqcgI2t9lKRlxu5kijM6yuB2j0WryzORCWUoPSxNIbJRhFf1xDdiK82
HdJz9fEvo/HwC4M9rv76pEZHJpoO/raVlM2k354pjwsZ/EuYQON1WBUJN1xMXwgQq/nQTJkT8Uxn
agQvLwbtxTPMZGwDoK9rey0dKIlpxU0KOVkjElH1TIwyrvPhtnyP5x9PVBQiHdyQIodkx7ecxx/L
fZ3YqQ13sRaB4yMv9rXyyOULM7n6CBB0nFY2lguQEyy5udrQUwqCAMLIq7q7W3ceh2CjFzDSiU5L
OZMaeQdapuCBCalQkrnWwxkz+IibPjTYUm41P6eSoFrNmjV+Ywyji1YGXWi5qVqaZCrNIXu2OUwF
CViKLRAsecTsJKGL5cCiQvN/JtUlsBanZmo2L3hcoRknTsIUmJGuxsNhz5mN7Lo6mEuUdZ06vYt/
iFGDkvBLDDMsZBvdr3tmntwXRej2VVLTY7UOCEKt6ckAGCSEm/3CHXTA6V29sry+5iFsQz/FOTHj
HMRb7ozdknzeRtppOnCpqG+AwENw+nMN/qANOPWEEldadUVxN6XpJIJoqLTxDsDxUv2J1HJFk87d
ePu+usx9yLtTSN2OFl34YLD/7fbRGCc9zRn37vFqCs47AfxX9VrBNGKVkmL1O7dNUS+dMdRyEWXO
upUO14dmBbU6oZLV8sEQDL1aFAut6uy6Ov0CoCJk7+RkmMvjRLAoiyVib8XWecCh7VUwBWFGCB7j
6LgNpB3Lr+obfS1UhSTqCNa9YZgYgDzTx+9PVqYiWNO/VfPYko4KNYuRqq87AZZgQjTjdOIT/6aE
5+WP4T+UCigZ2vPKuHvLRGayNBxHzpXl3aXMaFxLs1ik3LTy8iSkmjf/In4vbnLxbJUVbYAsZLnG
Pmi0/c7SYMcAYyc+tObbWR4edwybfR0wwJ1ldnDx1yQE3yXd9JuzFd2VXOdRo/zyD/p/mlkfbK2h
wamdf7/Odn180Lmor/ylJbLb/fuCiPdDzHVR0w9knLpHQwoSdMsgd7NxNP39jvtqUtJCzjvGkh/u
Kh5gQBK+MdIryZG1rhNq2VvAY9wuLROl7YTjuLgybPWzp3s0ZtsOELJd2TB7dSOQR/0PoM7sDWdC
VIlS2lYCeb1L4glJWMJUyB+8YEMRecVk9j2H6sJYRscqrRzjMf4HL6+I3cM9ImgU0KKz7mC3wcZk
F8swGE5ErlH9T+jNOEbH2earo8uhPCfs/z0oD6K14EZes4bCB6SMlnGumwBdJ/57b1O59SFi4S5R
76YYgSv0GNIIpa7vqsm4VVFnjxnI3jmoaW/Z7UiT3/x2t0FPkjqHMlSL0Db7l7Bu/LJXI4MReiXS
IsKxyBr+KMi0OkB9/wbNdEACFv9V+PnNhrhj04ym08BIPZiSMjJ46Aeh+ghMcq3Phl0JVzBPMTo/
3dwhcoAHsQZwIrVGNZZhzCJoY9hRfiqv0+K+ExSlQGEvpj5rm95PPS8LtnKkuF3X3S01SnB+A4df
WhJUA4j9wjwwXxIY4VLpvS+I065IbwkodQg5jahhL8gn+Zk+a7geAlb+12ql6MP13LTrL0WHSuEB
tfSyXDWZKRFweRPUzMKwP00+nIsuOtYVm5rUZE45htuRAtQBlAsiWRVk1r/e5MgSXD/R7QgCIZQ2
NILZks9BK32B/ZAl6UdUZtJM9nvMr0rKhT1LMG4yD9IL3RLZ71Ou1gQE+GscA4yzveB9A9PmNNNX
QmPvOqKpkEMR5028xp0nAzsXbQh692KUErl4W/W4L215DtaSaLIYcxBae9OG8DBozNZ7UJ5DiZzk
sG8YCCI68ERHKMMSjtON+ze5J+KkU+FJPGQT40eJ7GpyhrfCwK7H58LwT38QrN2FmYDkaGfYtpYt
+tPy+VAF106Ls33FkGsNVDo8bWELlYkDxjHEzRVQtE5z4Ob3cFBn4YvFbAsY/jply983hd7Ix5kL
sXM6IyaaeB0f0t9t5zkq74v598hr4ViQhylCOUvNvyz3vYZ083GL99B0cPV/Zg9rnmmoAu6S3HYr
VPBkR0Tl8yoaQPHMUNrMAUYgnrXiqB37aR6df5jDfQ7A3Q6Q6vhLfdr9CWWHk6KiSjZAvyd7AHsJ
8W2w3GtSJbUqRbxKtRmZoPO22POdZy6QZXz2WKOIbrUwo6jAA0VcZFUefvuaaa38S0CyMeuEMbQJ
3FnL36O3jQSAYe/PZZ7s76dmHq6cHGanehXel2LScvFq/2yxAIRWMf7YAUG1VDhvZ6A1xXcCzv4S
3wCJpuUGi/o8LSk4WYQc+YgN4I+HWg8tPieyv8yjfdKZqAVKMRjgvZnpPhcykf2kkVN6wrErFFyT
yRTURtqEU/ilAlrm7nW19tZuHpLAHXd07SjUDJihDaTz12K7OzkKR8XTpjEpzGJmPJUnKFzvTuD9
dUDiAasDAf2+MYxb/Qw3lyXlMMkN4fw7AeFd0j/vnyp0SyFSnwdhJp79Lt8CgsUN39l2v/yMB7CJ
1NJHVVrJR/HUItdQvWAkGpKiD2VTLBCuZPKgfl5B3IKhcuQh/UjFO5CvOR9Bvi6C7OFu9eg7NXn0
jFo52pi8TZO1ouVYcMapKzeVMjKsCd486FSNZbfgWre49Ms/z5BqshcN4BwXf/SpajJzqBBwTUgQ
0zueAeDnSVatWcoweuF+obUjxaT3gwbINPsG3V3iQAwmzXdtEug59dR9CyEluKoV/U8a3ybhzAOb
a6nkAHOQz8RKIkaH+yKjYU+syb0JqtStfuNqzTaJmiNfq7cZ4+x0tFSGpvr9fawCwJPIr6jd0MSf
74/CbSqiJF0do/sAd1zYGXrD6kNjDd6WWgtb4hSBXjGaUYvHgYKfHIwngORiGcYbv5ipbb8wu69t
pSbgcBJ4g1sxAjOblXNbxL4mIs59LypDkbJZiWVfmocXYAZixNO5Xq20F4UL1hV7qCxEJ5Fsdsv6
VdICS8F6Jk7IU+vCP4A3ylBxvyh+YI/l3S/f9Q4pKvOEdqgRwY4u/6icf6ZYszbG3Gbcb+h3HeLh
B0y9ruiabadR9lb6n4MCUPpx1BWu5WYeQqI9Ew0q3X4Sh0b0mCjXjvSbJ0oyAhm+oMAcigYkmDbW
I9VUYJsR3Zb16K4LLogfzVMXbRcNcvKFddWt6por0db7EMu2Ej42Fp1olkZMtz2iIGqe5hphhOW7
ACeYMJptl/OjpAsdILIOZy2/edZtMnO7MHkG+PG6uyae3v7AlB6IbZHqRnx02tFtVJ6ZyR0b3VNE
NUrn97Vozr9A3yq3tnH4bGI0WIbHo4Nvq7/ixJjQKczQZgdEH5phiiMplRJsh/mgSCS5j+di2e6G
ZGWJNUIGnhNozzHmt7+9X1Tv21EyT5RIAorqsARyyVmSOriPWuTPqteqIz7F3TeoWrjNFDRtA56X
ggWtdoMq32A2IDAnGwUC8wmuHb7Zir23XizC9wmwJPIgL3xsDyLpUFceLkwNNgq2jF+21py/gVvi
RnPIYADlOTTe7UjQZnBHxIJYWmbbpAeekHFE6RwPmjLH2gQqyoaemetLhzfhc+tkIMNk1+f41R0Z
F29IByt5gi1GNtoDOvBjT3IHfmrQcHmVjgh0FxcqaNuWxpJAcZY73ZOCvI22e9ywjix1QCXNKz8v
ci2H9DFP104kNuyWj+RdHFmZrmUwuIjIn4HNsJBEnAo4+HQmE7ug0PCax4eYEFCsod89I490NLkN
hH01RYX9FdYYr/mu1kMAKCEckTupBQ3ckk5BIyEv3t0cQRSwaAyjK4jSDLiNYRYbDdHScNYMskzc
Av050tE+0XLBjriX5OPQmyWSrlTQYsObh7w6iYzJry2vq8aC9uXDnC28jjwmtLa+U+GopFgSStRN
yyw3foowS7YrVgwYQbA7ZAOC50szFVo7deNt2i10PzYO4SjDHlZTB0rvJ85JBA8NICrsp6jc4cgF
YCEzeVwrF59Kfev6L2X+YcqspGwibWlfdjAHriHOFwWOW69b0Hnq+psgDt4lQ9o+D+wdL2sjsGBK
AhtZZqayOgmTxkShUMOTg/4BUD7cSF8bEL5aEVJD9Q/jOndhHKy37UbJFRN1uK0wgEY0WeMLjOj2
e/GSiwho9uznJNt4SL5m09GC0bp/KmzMumAGRIC0BiJ2whMcXd8O3udFjJmGTfgJR9WbDHX7E9wE
QSo/PnrCUeTClSYwMX1Iek+LBcbct87WtiY+7JLfzNAWNC9sIQRdjJxagvg7k6x5L2SoNczJibuI
NUuLzSvYLHb50Qos0ZaVJvs+ZMTyoMroV6eezlX5oezbzOTpkxBmiNodn5iQe0d8TV3FxIZ8DKWP
vniiOfIAY1AueYW7uc9XsYt3OOUnbL6NdM+tYzw2zfFjilyz616XbBFbNPBh4KkcPquqCHishWLJ
D7UXA3lUaSbx02Usd+NvUKYbBvZpjxBWwVvo0ORduUd2dxnIdawAsgRYMckSWtB572ijpplG4ei7
wAVLJyFj+403LGwmKkyngUr1bp/XcREXwCk89PMnOkr3X72yRXksDrQIVHfxWQIfZe5AUWdaQEUM
7CI3Qb5MMM6UUoTifRDqBQO8NjAxgiQLbyaiJrgJHWHhkCLMMvhqRD3exk0zhWNiuU6/Nc7528IP
yAqsJmOZaE9T9iUk9VEaNR5vb/KgOeRr2rz8NGn+3oWs5E4BUCUK0yRf2tZfvbCELTk7QHIQBqed
A9+SCgcLeACAT1/SrvY2WnceqMR/dcy7Chx4N1GVZuSL8MpRc8/suOf4+n5vqY6pnl5fmqPpXOfY
2Uo6Cn+9vjKZHEoYavLlgi/umihmy2BG5Avbu1q0a2v2HOBMDHQhV0xCdsfDXcYojdcNxqBhqAbY
qDWjO89+/ggFi2fZ5pRwOUbgjjTj4EYYx3lbGjO30XrTRPCDQ0gwqCXLu5HmKcuX4BoGsipav77U
Jr+4LHjEb/dtt2yWs4nTsgD53mGJcPa2vbymNHgNIdb7Np9eTvBFOcu3MTHRMx5Uxxo1Tps3XGAD
gqKiwdlkS71ctQg6lKLmJfS14kIBfkki3PIPuYh/9aDf3KIbhpQcGs9ZBfCUeWBIDc0FTFJsCJ26
6m2FrkQVx0vc4M4TbUuAcCDhtKjBUMYUygqo6I0KmGxwxmpiNQIh2pUZnCX59XkaWIO1EcyrNlrg
sZNV5B7cgN7ElTNrnnOsE26fMjUjULlKf4XXDBBOnPZoS42w1dZ6P2rBoFoCHMJTAs/7pcFRby+8
SvOFTMLcd84qyjKeRiNIomyX2jp8Sy+ePxmXbUSWtJsG2ERWenQUSrsDlpO0cAncEkGz843xIAzL
2YlM5ds3fULMsJXAsXZ9R4BY4r+UGftTJ4qu+c8RiFoBUVEf7KHlogi6PigqtEvtn1LsX+sZjtnH
oIf0HOxsy4bP16TV/Nut7qsdGsZi9uFG8Dvoikr4teOOYMfBW8bn9vOJia/IIEt+KpPXM+MOk1Yw
jqDyJwKq/nVhBbuJGQFYENqVFfJLFAMwpGcavChSorpReT2DVD8RpQRYc0JEXqiwGtBKmuzfP/DO
odwdLI9zuZkfYtHT/A0ZHR+KVuvaFzi0IJanK52iPMQU5xJ6vhR3Q/P3YG27LyI8N8FhCEUqlT07
8+nr4tm4734hnWvBz9q0UtuCoFtAoa9JoGw4s4nldnK4YOiwn75iMiAFyEjjN4hz+n6b4isD57M5
s5+k8ZIMHv+EFwSOHcM17n/WaT1FScvM8dYkZv7fJjJi7G5QnCdZjwVn0D34wiGWQGigi4CM02/W
k8kxxXtF4fWwmEcgns+TJMRQ9A6CCIV4GEIw6OrOX/lkEFw5kdWwkhwO0XeGTl3yG9TuAzRdIJJZ
dAMn0QZ+bQv92OkqMMPwZajJbtX+YzWUuoyqKz92+FEpsjmoi3bVaKpmROZuGw8KQ8inGxijmdKe
EuC+3H88BVv8HQNbbOTEe1+FNqOd3pDg00vOKBGaMz9HrmHuo8Ih3CXhL94RpbKuV7CLFEOnSHZ7
pz4v46sgbTPRptbTcYZNao5d82IDYEXzP5HbnmsIFJto0dPogBYsYLXTG7nevXPP1bxUfcbCqfsc
mxwKOks+G2N7fukufz7xR2Z28be69n6yrezQqGv3rBrRFxZtF79KeriSBrdJC4qSy7JRcAtD6HS+
SCLckVDu4xFYGatVJYttVot0tw9n1AffRWxerHzvQr9xLaRMl3OKKFFwEOjwd2SDxXId7PZjQaVK
kVMhRK/knhHCxAOldkJ5zzhmZB/oa2bIjoeP1J00VQUoMBLT5xSEKZI0olbgglqoFDuhZUwOd03P
HGLnuUq2i9RRO7RWaTLEL8mYIm/iTAVThneqB8AUdzAavGFxZfANugqtshUSBEkCJDgTaYSxcpFe
BihNyyzip/cPpfrP2WeJDVdHa91PA1EyyhINYC5RMzBHKFUMOuXmKnZiW4Q9TqXr4PbvObdfNpvT
dnDYZIAceaggIbVXzYJz1F0FWza7BrmXlvSkHm11aj/LUJYh/6pb7QMhQprEGwcuDFIGUADCWOi1
Cd7mDT9r1ZYoZ1rQOUKLdlOrN6QtEYeGlsn9gfWxcSUh0q3pUsk41ClLt/Pw6q47yOf885S4DS5r
/dk/8+x76QqFH6jiT//kogCkGNm28TF9g1S+Mk+UrItXJe3yKlZfrH29trbdTojl2dArzMRFT8cb
72Wa2lsP4D7Bvg4CO0IuNqFS1TD84O0/fLf5kBIA+539VIeM+iD4RHinUqV9SSwdrFawvFlY4bw+
5arF+dRn3XvivyjnXQSq5bcEZboa/DkRH6JWGyazVoZblKa4ToHq1MyUNloIroF2BcXTIcx0+PVs
hQnNCmDmq5wGF0ufZIB1/Lif9TT36SNk81tXUOW2fGm9cw73Fq3yvPG9oV1wGkgGSpQsgCv5mDd4
vthr77xEqSro5SSZ4HK+n8YHnOb+7LeesNagSM12AGj3nIzW3znUEaoS4hqshmPCHkpOMSmvPxLb
oP5PuJabKh+NDo5zToROC//PLEMXEWylOrrrTdgfPC7vnMND8WvaDN42u7ZgWh212v6tmvaL7Fef
9sbEQmEJshwa7DR7NXbOC60Pdc/o7UpKxUR0ndzEXNbsb5yUnntC/ZeGgzu1KcEDjwfeI/OBszY6
8zjbgAWu0uaUCcD82Y5KbmQ9RDm8VDRqudw3St3ttru6iZTGdSi6WTY5FD6wxcVT9loK1+OC77E+
JOVRSkNI8EnA/7T1AC6is6OQkiAB38AXDkPc5B5lmTr2TADLp0zrXMWoaeR01Vn7LBB5yPBThfoc
1PulvKxts0/AdIcGasXBasy7IlUAeQ0J4kAX1z0pMbrrGN5bFrgCbWel0S0n2TCPK0dNETSsiBVJ
g5U/aAIg2yfW2uewhz52bN96hz5CBCbkZ4vFfBz8ro1LUVuh0XSfKso9wwsSQA7Jrvg01a2RYwwP
MJHMMoNOB4LKQngE6l3gYxJ3RUYFcl+yHKNUWO5jqrIGx7vSGwuJkpzfIRlh1LkFKncN7uTDiW9f
DrUThCN8zMzYVm7ObO6L4pFIYGpHf8mueZnzEXFIXzdpXI1GAhu87ZY+8o9TJbO+Mk9ux8yMkrca
S96wzROqofkAamxYkGEk9dS8WXDjrMrBMNzFxBKNtGA+VH0hqZUlE4Bs4WgUmnEx2EdP8zd2xOpM
ABuE/NJaa4kUZU50ZPiZ6q2I7bExV2/+kpO2OLXnOzd87jxRaiovyWu1+WiOB6rDJOYm8BLR13iB
kmbbCuFPPTTQgz5DducDPmERa5QJT7FSVxOBnxjAuuTy/vczFBm4ljlKw2GcIs1k11czCC4FPuHK
lvCgPiQm3eLgbSlNT5GvLJGjU65KI8eFgCqTXNBWZZLLqJhmHLu/CIawW//axyAQZYPuC2/72QX2
rja1wOQFV61jGoF2h4Ujtdabt9qPwu0VVmLaJ5022epN0nN1sBme3/d17Khb2vsLf02b002dx463
0aMk6l+hJQsN+De4IkH/CowJNhmxuclEyh1J2OQNgbpvNEL8SAcRnVPhG5jsn7yFbY55+Ris6W/T
nendJMcyDP+YM/UJeJlBtjOtnsLaaSb95EaWJT1FvzipgIYbXPXOvFCQjhJ4xCutpga7iuV7klq2
j9r6bH4YWNVD0dOOy4IWKMQCxkKQl4HLr/18WE+BNedDsQa9fu6As47Qh827pHHcNrdkXpg6sGbf
BLaWm7pWO2dqgDYy4vZ2K3h7M+m+0FS8xwF8eEr9YZ1yZ0JAPSD4KDgI9j4ybEoPP8SJ9awr5L8P
AqNXxa+xjOPvEs7uwCeloNJ0lyC6oEKFstZ/Yi9OriiwYaQBRVlj3tt8Q8cLH9GK8qf9F4TQCjVH
/uKsxvNxAopQLxMDN4iaAdgdmu9Cbthfj34eMG+Q7iNFVCqdSWiwvYWdEF8W3aI4uHMpEHnV8vHU
l9iOLdRcEzSaSFYGRN+WQ+ioTEezr8H3JdxEOe1LEwn0fZhBQaSMXRB6DzRPGCEQGj1EzDo2/yoU
VKFuJcbJmTaQit+KxJrPrvcE0EuaCUAyZmReY/Vqa9Y3lzw7wrSLo/9hcXZxmrj56IDhP07e6mSp
TFrAvuDT9129D1RNdayibdAnfF9B2fJq2H17KLpIm1Qxdwwy5kbY/KB8IL63iAsPhfW6nKg9tcjK
cAVofLrolB52R4Nbv/dwfpb3BqH5nyAuTbXEanARZ1KpcWAzK0aYeVoL5CKvRJ2zPg3uL8sfaAxe
AgdUsvKcriXAb6c5k1mktA/B2Q4CsFPbCd6mOzxTQDxGwle5lA+gGMXQrerebv4gKzV1sQO2xneC
FZRlRDdfbs7vUPPfmWTQR52JiV5NI6+NsNBr9o/t1wffUbvLXYj/rJ/hh79+lHSE7iUMt/ieeQOo
/c5S4+AizWqHD7KEonGFTs0QADQiGOy2MF72fzN7hccJYLfCvP/3N9uXXHWAoMf/TPJXVBD4M3+B
2YaRLld5Q66D2qSCztk4SIPxmtEdFF7jbHXQfFEPvxxGun4xqPbA72oEXjTs8MtJwmP9TU2gcO97
/5b4CSihpmCYQCxVgkHuVxRPiUnwZ9Ja2r3eI5978vAPzlOOD+sv5LuMZqHot18F7Ob9l8yr3HdF
Nf19yAfAD8p/XQxlD/p4yq0HfLyupJVgpTlne6G7YaOZtsuWgXfOD1V6HLAYmiaU97+6Sicppzwv
/J9LDQhdUnkiMbJNVV5qb9zUuKc6CrxnuYii7D9EWsi16qwWVV7CQoj4ClZkI4mdSQXUKTXFak97
ndrlNvUTr8hcvpEEHYekPAKllHp5EJJI2VYnS5gB6KEK9UwxTLdHVERpMllHh0yvhA9H3XRgPkKl
UNviajSyKjtR7GG6vCtROdg9hpTOHflSdOBjwecFeGKRTaCSWAXKtD2umpv0wDfWRIZro1otCXDN
DUIkLgOD0VAb2/F+F09AG/AF02tqQt2OBZ+zv4q1b+G5PYlW9yCx9tu/Ho7Mc4T96sNZIksYpKx7
lurAr9z6bOsLSs6ewdFVWgzsISfmAp8fgk3d5/ODj846wKOOEq8Yi7UlzaNbBui2GCYBx4aDcjNp
VgguZl6RIgItpN6ez+jjEkbL8xL8fDyuZLDGIcYyCURylh9VfXeKNO+wNglbCmOdqFcMIvTRAvF4
HRMivhY6OC5TrIiNciTzl/CWhB1I0fVIanqGvi6strRDvz5xmHjlFOQtWeRp7/nrJvKv44Wh7uCH
EMNU5ZVkT2AHnUCnBws+6whenTRwbDyU75JPJ1JxhEh9kfI9Tm45mFQmpF0A+T6mPa+fVm0HV2vA
GUd+aQZnqJ7X/pjH7Jt94eXRyzNkRiR54dwHyFC8qQfF9ugW5LVZzk/fXp4+3INFjy41UegrHefZ
4zJ/SZ22vIGu6MjoifVogZ1gdcOTQyZLDtY16B4SW8p/DQZ+mcUSq+B03pYO2SMfJUo+S6si/EUR
+bb3ep2eOtf2cq8ZRT2g6rFdWo1t5LeaXWldR7gVscws0byxIulJKf5LRbY5nDzT9Cn2cQU8NmUb
9RBE1V+dEEHzy35JpSPEbeLHSdCPAs7zwaawj+dxyGZW2whKgTCKa9QrGuVZVi63Kn2a8UwtgHn+
SKCbQu7vu++ZEjAe73StvXVGRwG/YunYPA5/82kLEk1PxJHHZ4sm+TlFdn92qfpsiTJpTBTuGUHe
aZI3rWb3qAbnJAlZCeNlk8tgtf4+plFl5bqWJGt8MW/uYj8PUXxU1Gp26GG7mOLJe6qzz6Kfe6FY
kPvGBHPd6EXGosldRw/ymmEkutrZdlwwBuD9fGmk0qy6B0Wk5Et65FurKNl5pGC1cXiKSqW4hpF4
Wu6Vhb067n1Zj+PGv3poIEaZprOzXZBsmi8bOgHP8PRGuoBPQ5myiveV+DH5x0A73HuCHjgM2iaw
XP59kAcV8BDTSPTtKT3AHfdD00afKjQ8xir7dwmhpc4byA+Zfe86BokZgKqRgbA001e2EOj83pA4
/PPcU7RkIpvO+s0mKBslk9kN37+F916KT7wRshGDgZ0RVroD0iKKVSgk6OHbWChUMEL8FaGNdGTQ
w0qXmQ7Ip10x0BTiSQBIMVKayK6B/Sy97ZmbHGowKvm2AIyAvKY9/zh9MKp0tY8CSDw3MMuFcbY+
yqJA5kYV/zBFLdPf7rJgZO88leh9RR9JXbHvMRMywGL2JSXb/MmiCuZzcYKBmvFrvPN1/XXWvd9i
W9kAWAJqFE6F3TGyLC4uYOPpc6SlWaph42c0jF3l1BXXyUc+A4sPM3NCoFAlXhP40wuEC5GwMa+s
2WyaAU6lPeSC7NP3Ym4IiPgEy3iyHrCFweW4DbrLuF5Angksimr3iC3rbdmhrpHFtXqFrS9F+mz6
OpaVocNEo+Hbeo42/jbWXItE2YtjXrnBhOkY/3EtEZiw1jcbBG0DwQK2KK/L+oUIo5dw208jbSuI
f0rgTrmBrHox+5ctL5WTqh/dBOMQzemKgA13XDM+wZnkG/YWEyZgKO/EOGbqPEpY/X7YknbMOkt6
xdXNRa7+n8T2uU4T0x41uiTjk+nqdvU0ZctQqgR/AQjqawbqTOPDFvPokMz6CR4F+OIOXG9limYs
OOgovoy7hMNEDGD8ahcoc+2FuZq6zlDqKMc8cs7zbxyiz58a19hpq2ob6JwNz3bD7MaB942kaeqV
xxrde+zpGmlfDOIYssKAMkUE8mnwW6bdjzZbt152D2Mj4udvOsn8MIjj9O48/y6Uz+aSaS3NYk6Y
KRQkWopL2l4TSY6sPizx1xljtEBXpbdQPRTrdBCyhbKn7sLRyvobG90HIt15BUgQSBXgz2NpBoln
j5+sZBZKfmbNNc2WMIU3hCtFBU99OVxPsT9q5uJGtOp2hSi2kMGBYdEjPzOwj/ELiUP1kuOWtL7a
4rl75igHraUJvhuejGShF5coXVKSOOJpNdxyPDr6UdPnEwRHh1+of+ePBSREFR8OlpbzfMR96ECT
MiLNZoxiX32Ne5AXGaA2VtGw+ssU59eRYW5kYrX9/rZ7lxYc4qHbsrv0j+X9qID2c4lwc9mO7DQK
EnEPHITafX2NJem2MUMZtknf6OneVvWzUMAwG84XR7UN3faUQ4fmscDR45hW6vBRMDntekB7iPxH
AaA0f2t3OTa8gE+ofEKcdcoaJXIhgG3UYC6B0u1UBDHXjy7H4I2kFvezaFMFVXDTaDFYuKml/KUq
GQUVzNqcXTzoQ8FHzKB0dYpwRWd5CUr7ccIyumpb+B8xzZKOGGA4GNCH/6EFfTq7nGBArloX3VDJ
DlMzIgJyXSXJWjfjnF5+OwRdmQZ+I9rGpjCzD8CXrrimiWnz9/C+HrW2IiiuNKa8sY6sFV1JdcYC
NGo+Am01CT2GnE1IbFiLetyY1YIoRR+q0JAt6TwxFpktRK6dwZj8Lcy+XMnCfG+G7A59YIoABXDb
nl1NrLTCSNF/YllbHoMnx4uDOfIz5eWeeBD9LbNVkB+uMqBANsnLoGu0ay26fzCVsjkO8Mn+nLKC
+8zO1c/HiCQrd/cjVawkIQ+qSUT144FmLNZxan9bIpvOts8du/DLQXyVPyFRRo+q+cSVzRu6hCO3
gtYX6Ebj7aRwyXXmw4/O7WAESWlzsSAgUcuhDTrwJiMTpbcWkiGrBBGq742Ui85mGzfuEITAkpqk
xlmC7wLbQHi+4xtpOKvM+Q/NfVrFXNTEGjlrbIQ+ApIZNzPmI++yRc34RI2KIDW3sfp8il0KeBbx
5Bg2eXxqCommAywNiFiBimrQDUnJXxKIcIB1l19ZPCiTQjwMHAgWdVH5nncMx9QOgRlcTWYjfehh
I2v7Pcg2dbrm7fShexvjbk99HkOgV0qGlT4aqYE3iJZB3kDVDEKLBhJ47wl3RtmhxzyU4uWquYHR
JgP1j9L4q35E9OrvwpnhjT6+orOt2Gg7s/7B9/TPe7uRNJuJ3Uins1hxJDvt84h0p+l0FW5FX8bD
U2C6vpno30vsHhOIuJBP15k3UuMcE05A+D8t28yfKhXDmdbzxdioG5TPBlfrsUPCPqPhmSkSL6IB
WCsBdrUxU2XLD68eKdfPxEpuiUG0WI5z3uiHs8RdwxPVi1MUG2CvHxDG5jF0oAy6AKL5Wx192DgW
xBQM42qUZ4BW/bkCV2PIdQcvCVAbKge6ANpTGsqNGRWzy9oD8uGLpiUAv7nPqOIDITTQ50nCJ8LZ
5v31J7rF+mPDnPe0oHztw0P8mFHz4o92FOtYMSlevtSQdPPE725Wh9wttTvT2E31TgGBP83hduJ2
kmUFga4UcClqHbm18vZVUjhbdTAkDHyiBRSuWDSFsv9qzYiPztdavO1Oqi41TNuC9QiLdq2F/66E
J65SkZ6G8aI8AKTGECJeM55l9oCNwNWvXLcMQ8NtsD2ZIvbScskGGgXNvG7la3ykL6YT1tLHLQGz
E5lFfIYjoNg+tNypC1R+NTgLyzhvfAKB4j+argqZFmsj6zW9cn5pgRiSHK/lPQbLAtwrDkBqhhcm
g1uSJi5nhstcSV2JnmhmcIUU35K5EFY5vnLFcJBKo34HxlWw1tfh1vGUniFqijpNeD7NHYh+F9z1
qojg3Ya/1OtK6rCz+hEQzVdgt7s8VIeOnMK/lNlb60nFhN+f5D60J0/gQDCScPNDPZOk0t56pCYk
bUlSZkqFVqE7rMi01qYtW9e8sF6gS/SWqp+si/s/oeLEDZPGGYBD/ZAKa3mAN0y6P1ZjiaNiResZ
FTcmwEkhtsb5+usrW1Z2wtR+10jlf1K9N/qH7iHfMiRI2dPcqdhjBlSt0+0Eg3CtEoZER6+Sa0+1
DxKEHaQcBEE2m4tCVFF+EALvmSh2HoqYlpjQ8RDE3AcS19dzfWK68gbav1sKSskZiOd85K+PsxEN
Iad9DQ2W4YUuvAqU42M7s02FFrU51fcHlKDfOQUl4mlhay80FkNygrY0fSSJEE0UCLA9abpg7ioQ
Cf2ZDhHLdKBAVbPwbE+wKBWlipMYy5XFj/QSGc1/5hA3r4tHHObR3UGVZRjHMPEUw+ND0YH34ODQ
i3VWgtHTNZDtG4NoqVxzO2iUITUoXnpZbE5O9YViv0b9K4kwdYpKNdhSbxEIajFsWdjFx2RejQH0
FdKic0coy8WvT4sogacgGYjxJGiuKRs4nalHqPGpdCDqvuJYTfrfqzyd1Com5ApYQZBXK16igLm6
O4ouO0gTm+fSoPV7bW0ysxO7eHB8wpklFENfyW7a1enwsrj4Rp9MX70PHLKH6pObHnBnB+oyuiTE
5c5yWHq9EPJk9/+MCxujnI7hDKTSwopqfiy9hy2+sAq+x/ED1nqcz7EWvF94FSzF7/9+C2ji2kUY
SBedC8Znor3/sGBrz05TWPT3iJ9R8IML7oMMHAMtHk3jSv2KC/bckcC1ueGNW6QJZ8ays/z47M3o
6+f1FR5t2Ip03auiRT6L7LlMlnJLVwc5I0htWfJMbuoWD7NoUG3zI5g1zHObfxG3zlBEUF47/7q1
76LA6QeRVVBcQuSoFQJcGL6dtKbob2khYpswFDTWPtQ9vz0q5WKsLYevWme21hSJoMTZ66qoFDye
/AYKbeIJFdY0HubE5N2pdu5zvWAhaXpNCjjQATG5Y17YxUsTP0hI3RHKdCKP1Z/MzNaJO2bYpplG
1+xkrqkVIds7EwN6pZo+wG6VNLqS5XKtmL4jQtpa8emmUdRJyk9WyR8vxB8nFFLz803M783UkrC1
Uj6CvZCVEj6jRCx5yFhnG7gPcGnvi4SrVWh1zUd8iPCNhTid0sOl+6SHolQtfZS8nMR8XeMu0P5z
NWz1UjK4SyEC3CjJ5RWTNe8gIc8rJtAsXdTwhVJNZdS24DZrg/Q2IMBu2mveJTcUtcfYjNkviTZg
5WtEDrs6G/74ayuqEApJRnMfz/TucmC3fgtD10eHkxjiDF9rSqVOTiTk9AKuOYH5SZpfJp1Dhnq/
bm86R6vT4ixl8EWtpfVj+D5+DAc7Hf41ydeKpTBZhsb4BpH2i/fXm5nVQ3H0squZS+ZgEC6pHFd1
WSkY6lflSvJeW69m+lxWcGmI+0eI8GfWGLdbwNa7HEt5AGt6jotQJ6VAZ1X4CrDHfHD988Jx28gf
iNDSG4Ull9edSjDMs/zf2QGz43HC0xdBHd06IcOouqoeynv+5uZUZvMjrANEo0YtwUAT1FLSD6yY
p7QnEvWO7AOx8TRNdahyay1lY7LsZzgJS46csCZ3sG20BokKbRCaKkNOdLBdzRY4C5cUqO/cQzFm
ClRutq6K8N9YHSrvxu4l/13jrPKHFq3jyryNQFyDfLK85RwUy88zVYzGARiXGcvUMWYNsLOQDnWi
huQhuQj1JwoEHgZfGKMsrO59O4pwRE73XkXe7Cz82RmxOC2FDmXwsxSt+Bz5mr7qmuF6bkCKJPoN
tC4+nL8pewyd3qs44dXNSX2hTFIvLOBcBSTslSYXTiKSOntZAoPQUQLrZodB+y6LcYEwcTvKCahU
omuLZZIEHlBYkmL+3vw62jivPIaTGO7v/PkkpJ3P/1w94KUAzqbxvZFmqWpkPXc5jmVfB0r8dKVb
WmEC9qlx+u6mFgPqgLHLwsPZxK4e4r+Czhwbtow4nnKGyQZgSAkAZdwKZd7TRP+Xqctkjzohhl0q
2fXWRq5AaWU00fKdcT/1rpO0MFh49EXACxnQxCCBljLdUc+WazeRKxSlBC9ReprC3Lhvz1V2e14k
hJYN5NUSMHHuZblfYxniERbHQPdqGxN+WDJb974jtj0/K4+jifo4ohEKktZiTQOiJZvJ56LOQZL0
QrajX6JP+aeYsvg+1naL5B0+xX77liVXWb6rfJ5G3uzwnWOVLG9L23AoYz7nVjI5FryebKBKOwe2
u9woq4nFSnENke8D6nxfrz1b9cprcA282sc7ymiXY+vMZJBfysPwrzOcnzO9FMFdocVJ/eSCDqop
4cUZ5IlcfffAPVEMH05aoesnPrxoLzy/aCFa9p1WNkjArUW32EAIW3CID/CgOYKsW2wUqPcnjCX+
l+fBhh1qEGj/7HroDc81gecxfPEsHGH4eWrdZobrclBpwPEdJEW9LxQMu8UVNVcOjCqg4CSKjiUl
rf0vFQ4stF0MCLbNe8XLxmNmJWgSnpKX/c8ruKZ4vLpwVhH26+e91ppgrKPIfyeqz7xiFrBzTbji
+/lf9Eotpnx0sxEyUC6tnKiQ1kduJscy4DwHbXEJjg7CEIhQAZdrm2C8LESKsePdsb2k8GKyHwXj
m0Z7DFZVeM3MlNQU4eMGJcOlKU6iw2AWfZZsrtLY5xf7zCkTL4OSYxH5PmSIKGugKQjQ/fjVCs4I
mBEhuAvpNcaQhqC70GeG9B7wVu3Qej9ZrAIKy6aIy0tKlwRnrlVeCb15FG3WbCAAhpVM41S4bU4O
laGTF6gqAxjzdM+PIEfBVI4Hkwh22dIMOPeZ9Kbt0DjNNzqWsBbzff1yCtWOaih/eDf2m2m1uCJ3
AURqMVVR+xlE4IPxDe2jaUahkiU1RWWYK3wn1QUTZ10egWOJQr15Q9Fm0lR8fF8btyP7Xk2o+rO1
nPvVnfYFfGgVxRshPOgW99ReHivcn/Cg4g050esh2r5gC00iMYrym1sKfhyzgj/HeiAfHkRNKZ4y
ckm6+/ukrhX8uJanh8w7wKRIX7qiOsydRwv8G5/ZI12AAl7MKDsHRjU5Da3nBo2OJBP30ybtArUJ
9Bk9kQwvNuYzKOlwk8uIOAmOsu1MKKAmD2vBaHMMsokpGBfHODPBOIusE9/29all9OEWaeDFcRG0
vmvg8oR5bUNlHqLn+hN5h5rcel6cmxeKznrds2r5tZpQmdqw6TiLt8LqOs1jRPHs0UhbvryMEzZs
Pxz9aFd6Ig5M5QQD8c9zBRTQ59a8ET4t4U86MlcHyWBs8mIHEa/MQiDPgsm1j9I+fXVscPdZUf/k
oRwHEwUh5npatmutXEcy7oTCx8oKdhPWO/o7/E+FV1YlRzKCgkVn6R72rgK4mES3UkLZyZVYteLI
bgXB9ZtvLmmU8NGLwGYHcCXYuBxB+AdpprQJVxaqx8LsgnqxaCodpLaUIapz63LqS8ZSILhF3k3h
g8YfAn26II/0w233pIaNj+lt8Na43FycJUA4K/k5Nr7cd+uWw7UDa+WbQttrUpnJYEB39Zm1FzzG
yWGY7HzWg5bzjCY6hkEWaDO301fhj1DfMgbSglPvNZPLckvu/GyXku077ARm7VHNtbZ3WXg8xRxx
2uK4AYy4o8fD5JqqIsNAqw3lMD7xnp1iwq455cM0e5p7jV3qTQXb8XdRViYdAmlzaf2UvxDiZtTg
RFd5APizDiPFi8izl7Nb3c1TIO43lyLLxpqxxBaNcm/FhBH54hw4JOdi/EXbMMIA05VtS6I5avKg
aIEEg4iVNqtQI4G3NL2c3ARiCQuAWYFIx5fSUT/9PoY6N5sgI30Lz/oX/LS5N0kVo9hpXFkm3rEz
cyKj3wT/VCll55QIEpXhoYac1dPPGFzIfEMxwBM6idVQPrGYmbVq2k3Wj+htykrfwcU0tOGF868z
Lwa9bMc5D1veTE3Q2LBM/VNwhnSyIrrJzUiQyB+3jIpfa4imLgL1vZYMWG92MicFxwf7MiFzAPT1
qpRRDQwBOLudTZLmlcCXox/DzC9r10LpRnJ0SArtguxTER6tL/xPZSNhQ4YFRmAnZbawn7Br0EnR
dH0N4XmJSCcks3FqRTZyBiSriDqH3dM6hLYltRplQOq9FHdvugYFKKhga94rAUmzMjygFwLKGG+K
LQZtnHBVAAGX+0XHKFLtjxLctJt53Q6os//bz5kscXU76p2nJD7XKEu2EMjDEff79U/e5405Ow0+
TiOEXXipKK4FEro2L4ron6Tr1u9fl/PgNv4q5JfrNDZOWPKwrPD3XQtYWLm27lGEe7GhVhGsRHSJ
rprEnwyppAogF7Nzefu7lWWvtfOL1u92kpfCZWy+s64sEK+vCHmURzxC9Pco8VwCGSGLIa2DaJJO
uOADWR5iREFCG/GDbew5m6xAhpFLaf8QrN8m6ReVsNjuR46RMUccOYT/QQtibe1rmJOqOSelOSQt
iggt5/lchtnRE9lcjjLpRUHddEqsqfUA/DFVeUVI4gqGQz6IWl/yo+oKyvVAUer9dOCVA/mtdS5x
nlgR5Gvjh3fdWz+IwICx1uYP11taKo7wD7OVwYZBrEPrv77Hm1iEWv/DIVfc0ka3wKL5kYD8meIX
TePgVW4TnKsfEGgEImJs6uamu2XCYZ8skt/279w7n8/IvWXx4egc5+eAu+EyDIFuze9UI9J0S6jV
JVtzZvgeY9Y/7y+GeSxTX6K5lr49hxb4XdL+6MlKhpWZLb7ZvaN1OPOsg9Mu3TdwOt2MITJ5a3F/
IyFvyYOwx8gg+YjUsVkoGDjpTnx3IJ2wFmL0D7DJdTY7ljo83H9zm0m+YEqSP+AFxCQLlxHkh3G0
JmaezLup6Z4arqlJRNqtBjZ0RW0V5/n0lte8cn59tyHjb6m5x7/Jrkm3no9AUvoNoeUncROQoxyM
SEBjJgvhb3+qGgfwMrvizLEw9qUfGib43qfXyPEYQBPNmwVdpqBvdrp1bvcAG0ribIbXQcBgpugj
g8H61NEuvjCwu+CcGgmDNsXDbVdw4Nvkw4YBE/Elrxz/9YHy4LrWo6HNGeAhKdizuxFx7xFnTmHC
rFvttrDzGK+w0RyJlU3zB96F72z6BgQ6BSLhCAlnqkItRrm7+yjSl1ML7DgyRRRr1GayN/wHhmKO
2TlRtwV5m9KuvaJyBCuww/eKpemtYBFqv5BEox0Px9MUdPX7DXmsCcf9kekZEAtgQC9nQwd3SJ4D
zJFU64SCzgdjnFuB2bHZ78erh5Qe5oOJWQNtnvluYfHVAbq9XuhA26LDs5Cgy2dg2U0fFuG0vx6q
2fNRR+COOhopiE3i/+LVsrPXTyo0IFXvASj+fzWruPr5zxzP3qnBr6eiMLl1XWP4iqtL3I3icfLT
bvVGH/t+Ut032Laaae+whSoSBiCCIzI/PJRJ7Tyb6gcAsd7kBjKZApF40Bm5gho07oyh03pXvpu2
AGJH0sSr3psjhFhzVP55OscgWYKDNHwoaqoQevCCKW6Sfg28qWBzsoZkVM7AleDqJzltktIDdCFq
cvzNN614bJtfGUsnadXjLAqmGXfXBfBlecyRl4F2a5Fy8fPmVk7tL05RTv/F4vflkxHJqqFrL+ka
3zeI1MEkPnHeNb/1Ywm88STlGi2wGRInJr8PGWtHEokaKjCrybdYEgoQ1jTJB12GrcSOrr7XmnGe
wrvyuLZYd69ke66Cyg9Kno/j55DJXuWccZGDgaxc6FbikkP5n6GGchOyYIf5Tk1zqorHt6ghzDOE
m1FsU/48uuV9TOrOznqpPQC4fMzaJZN36PNKaJgImspMPOV0kN7NsEz2FqAYcNNFJogzEF4fte1p
vzCICbkRi1MUKZWP3fgOHaJf2Z/Ab6HxAV+E+x4oQ684kLhaQ22GkdMnTgaMTFve3cavYHtLQtXu
fH8RWMAPGH+Ps2wjVyBNshNY3pvEAIqoiHRyNSw5mF5ZYTVY8WgsC/Qrf/xqpFVuKRof2VEwSXVL
us/llIWgYDeEEJ+eaTbng6idlkAlmXsthPpZIPQ4xXItpLeGnWpqLnlAECzA8NlV15CEATaACKnX
ExJH69if4a27naxKo9srl6kHW5JiS5VYqLxdESs1KJhM8XIW74CXA5ajqn1ANckFcj4cJlTJAW+s
aGlyOAreTC2iLeCpw0B7Bwx3uq72JAefZDEoNsS+x1L1ymyGDy7/Z5ceHNFw9+E2kgE6MBl14o1c
Qa16UdXOCsSlzdTwa6cHuYj39gKqSGDzBC4AtnWufOloUJwOJNbEfm8WyuLj4cVKrVgspJi6SD66
d9LfpbgH42Qb08Ko7f7pNyPugIelmgMXh7kcd0UcS6ZrfVU0SICGbkg2sBaXxDRhS18Kz0Ub5vBG
iMdWKkmun+kxPbIULZIT1FhT1xdvMKdMgYg5Goh4ApUh65EEhtFrMYBgZWQhN1cW5eXRabHLo/LN
tD3yo7wvq5h5B454CEvCqRQipuPrtHdz5cbWHbbQhe6bsvEVpQaHB2xw+hv1/UbmMCSRaa8G6bFd
mi/anb65EHyK6CsrRDoMp+wI3jNB0GkwJZkqtmdDtCv4JCupkOAvApbNDL8yBwY7nicjhlpRQDlB
5acg55hxfIFujbd3ny2TgtdWhEkop97zxOe7lXhsVKZLI+5d0tIqjn5PiQn0B/EXc+KYigOgrRgT
i2F7PYrk0te9q6XDQRHJoQ7qNPL8lxO5QIiQa5LArwN533cA+VXicVE70LVLIxGjAhkywSEOvOAE
ZBF8fOGaSNrrbNWjFuv4IQ152ClVkr2CbC0igoiQknSP6lepKK+YKNkUVYiFdhXH+k/uoOV8FyPf
3V1OshtnD+dHWmqx3JZddKgdWm6ATpbbkap/RcqBfdCvAyn8xYOTM68TVX5AbK0qfMgGWZHPyeVf
tp1hEyRN/mzcljw8eGcoGQq9CX+5SzHXgptYWVwY3Evr9iI3iD0YEVAfFT9cTsKJOF0kIRlFU+mD
bRlMjw05E+TTkgdHS5PyOXK3386mlX/sWxaTjIVhbKIJBUJw+HGvHF3GkBV5mOd1jfpcn+UZLriC
GpptknpRawE/YPaWDPIbZORIVrqfRZMWFhLTphP+wZylW08IcsUz7DZcqXMTHcjPa31uUy6rhoBT
N2kQ78E71qm2N4eFh+qPr3+yx0EPj7QooX6Lvn4FGaI2yNZ33dx/qBObRNguZNwlGqfPC52h3ANJ
hI/eODTViOa7bDMFVhmbFhEAJa+/qYKhaYQdM0nCfgGFAT1yeV6QvMLN5xBz0lUNoNxcwchY1Z2A
OWbN9ME7f5gmjolHIJmycKvsdy1amoZ5GqZjqVEwQ8OiLUn8tMWOmW/4cISAz/tTlYfAEOp9f9vR
bRMwdiMcKh76Yo88iJKIqByOPx4rD8WQAaqwmB4rGc4pNjrAZFuewn777vgqER5ijJ+53ljzG/PT
O3Nl2pli70T59gorFf1eQBY0/5h4uN6v2pPUoLnSJ7sznaRPX2D5NiohClQ9LOQpx6ksOd9s1zX8
zC9+b/cCHby5iIT6BNI6mmoCO32M68wyVJLVanaz8RcV3vy6VeZ4b+5pGWmMxcqjRWLzUalqj+S3
KH0g5RQueVrf3kDKaNvLRdYyEtvCUMbsfWsrw2Vwp/NKGm7xfDisRy/MbGGg8wU1YYgkYnG5T70t
hdvuZVQmc8LQDxCKc3mLAFovpG4E3mJxELgmxLmqbk3nQJ9gqIeyzVBkXEGZIgZXdebuMTWvWfKV
kXVEjLL8ZU1KstgYOFvlI0raGgXK1uT0gK2eJ86i7oqmVg/5whRpMmlXhHQrCo2B9BXq7fmScB2/
VWfHfubqb7KwedsrS8+hjxfpJHLU64PVCefK3zETXvpDnxl9MRkdHDO/2Rfi6gqjnr6KU0nfcHrW
VZEBoiu7kMDn+KkwZrQDqGqzCTigotJlsX9Tp1ALV//6cE3BiyIOXOC0U1mkAtgM7UJeOjHFZBKl
ve0w3AGaFH9W5O4ECCFQNQYSO3FsBal2JdFhV+sDDAPWjpn2Qk9kXRFTUEIWcVDuz83vNiLTmEoj
BzAiMdKiAvUkGlkQPZaE4fnGUZcnP1B+mO7VTp7Xiy69yNIy7Ep2mhtUpjnI154neQPd5V7nL84H
riDLPTMAZ84wVMnvzfYHf9g0OURQ75zusRK8ylNLY5cTu3F/LTs2GrGY4/qQLN/s+rKs5tGq7ZQe
UpnaIFJ7AgQ48P9Bb0QFUr1Nc4XPyFT336+Z99G7PwKRQuHeL900qKnV0VHZIQv/QimfBN+gOBsV
LUxcmctqlzuAx8I+CGfGjFj5YjgwxRdSiBCSeMM2/k4o+j8l1uWOMasS4LR5sxatkJ8Bq55Q8iuS
0PWDghXUrJJDzWGuqalSvLrT9/sdFrsUKWzyI4804DahaX+9DmRrpYc011Do6YQ91bB78TC2DPzL
yNdHoZW6ud+MHCC31LzWpceA5mNOF4UNFpC387xtUaSVpuBDz5D6ZICCPpJOgP2rrCXCVqFxnV37
y3ZTByGgcy/8TrzvSuAX08J5uKl7ShT6PpGS4uE3WDIPkpRe9zJY6cKh55vsLhsAP+nWchLDVYFg
IgNT3omkjGD4hrfXNlwAyOokBd2nN+mJv6X7JxTLo7vZ4wrjKkoYSi7z0Dvg4PM2gc/epL86CSbn
ZG3H/lSRtzSeg5foZY4Wqyf7WWR+wTreoDBPyDc0k1lT6z3saV/NYSxSuEV7OMO+sxoSWqG3v08G
pyj44m9PIClRWZIfc06q91itK39b1uVBHOH+eTVOFQRVj1v9yCjVaiapBqBJ/7GVUxbH6tfov8Z2
QWpTBsFP9tMUn8nv4btygP/5gcfoKY7pSsPUPlpnGvbax9CA91p02DlSaFvUC6eEb7CV8Ob8UEok
9qJYTZk6OO0HWNIdFMqIbp9cTyXTURaZqw/Vld9rS6r+4SnbwI3pN7NMJxqa3/LJdP0tJrcf6YD7
Sne1tJBNLaD0hDD73IaKHwecaQ3YN1rDnCXxFv+KFt5N9ibT2TAkWnSF91GkRXkDC6n7l4V7dFit
WvO4R/yRduucvuKf/mnpyxuC8JXSKCHD1WHGuymvlnZ3XOBfhXmN1ILI5r9tkTngm5RtzgQ9cH+0
VuUyS5iZ1DSM643jiwvG9iL2ac5NWCb7ca7l6yx/YRuJmrceqNDTSRzPUGrg9kyq9lWMVC/k76Jn
HSFftfCfnpmkCdVH7vmxMJE0VIcG5Ja96ovHliMISvo7KuGnc8LfXLoRk2tREOWyJpDAfDLib/Cy
LPS1HD30QLu+wQ1aBYUVzX8SnClgetgGA98kovtVffKU1dCwN+8ymiDANqRERP7a5M+/xyp8Nlji
zdDdAbKaSaDPzyg7ToLfNssn0dkDs+XkGDvBfhbudsPswif/+X6n1YFanFNWCIpdKew0PUk5IBf7
8qW+khlZq6TeiNgel7KxJLBhXRikeSn7ta1UUUOGbjV6B1PqakQdXdYQ6RA04hnO4bFfBXvNWHGp
8dCsjBIqn4sxFwp3gQ7tUMWLHXKl/mhua1mDtndPH9y5HF9yWznhimLPp8TuTW5h6mzzoYwRpONf
wqoFA8jOml868xWgKxT1rN4xLl6YfUY8vDkCk+Hu8AA8R8uzS7vVVWS3xRyR9U7x+oHQGZOgUOgo
Z14wEUwCnsAmtm0alghRdnGbVUms+tRVKDHdSzpmLa2S9g5R67nfPnG6hpAZqi0GjaHeD0y5dqoq
19hegR5FhJHXbUTFAHb7TvQxV5zr/4DJdti89zaym8aSBMqIRPVXbjCoAPb/dw0Bo5UYADZxyr2z
ejQmmC5Rugrww9nOceYkzSxR+oDVUZUgRK/Oeb7JF4UzpWGUgF3I5laCWmnUTvjbWO9+ecKcXLhZ
dR6Q6PTKRda9mfg+AB4Lij69MzaQKqw9qzr/5saJFjKM2Wl2z/9LTi7UwwNhM+/XsRKdkIkbHHzU
GzFXioKGPl243ZdskPe1x7mXL0EbP1Y2w3b3yVbJ+PaebRAn7IG8I7fwROQLf4RdRPTU7lh7SoEa
O6hBJcwUKIIwwnocM7MgyFDwba114bPW8wgQwmDb280Pj+MQ6L5PvOLHDZGrGVl35gF4ticNUGNc
t9c6NXB7RBLBneMlHWKo+RNiyhhc4DRAB/foSN0I32Z78VHY2YtqMmc+djm9rTA7a60NvZJWEyYV
//Ho/1DkUkqqXQ5Y4089AEXGQqTdwjUv1lJmcvsrGf/mfVAW1nnpDGvzJFqj6bRsxiB5ciw/TCNT
3WJcsOyxiZbrK/JyyTHOo+sLRBXkxAV35QN+OluIxF83bjeETY7WyNCm4iw7ifANLhKI2F7MO/lw
F9QeM9UDuZ3AnwXecogvk8iRWnHhnlzvEMs5CF+2+qLrFHu0v04V80R49euzn7k/pOmZGaxCx0zj
yWuJSWuy4d67R6uroLvafXD3ZbNG0ervtrZpGRtNdNt6+vkokWl5PMf6sM6jtE8lN+lmwGYXvaMC
akhDSU0BuzjJ+8xPmg8CI0chBEip0Qko+gnlf7uUEiz5nk1OCXXsVrZNy1YEcc7lUTcHXBdGtPM6
AquQYBmyapOas5K7uWcd4hBDlck6flVd4CA5nlLy2w9WkhcPwXhaYa5BKC02T8IrAgiiWSdDSksq
2LC0EoC7vHxEILl+zYN0oataiAyJbxA6UAK6o5G/efpRN62WTzfq5GIzVEIOSETOMHvoy5Ym/w9G
i0ff86dkgTOkFuEJ6kCh0xEZkzcfiqsbuSvdFGUPBMLYMkRQDUNl458BtEObENyiMCW2icLyV9ld
rHD8/13lyRfGMTV9dZ32su2BxH4O4ua1tCywQI9hMJQ0zILK2lScdn6ok68BuTQHRenkahfVh4zA
CDUwTM+ZnIwwhwk+IMTouZ0qedNDc4+bzldw5eK1fT5LTlS8ubSqBLvF96JVeZLEILVC+UbbKXw7
qQBxzIi2CeuRIq4g+KVN3Q7FnMhKoYxy48Li45P2P/aQFZY+Jd1+XO4E8bwyvr1KUlrNU56QH20O
gwsQZs0rWr0EsYBo7JRUOS/xX5BcVavDMbPKn9U52fWoMfWSh1BWl4zcPEQmdcUqakKw/JRJOZQI
ml5v9fcBVZT47ZidRgRmMmoYoRiTw4dsEttOH92eAzEFJBfh3iGvPzZZDh0qQUbi06DDTvV4U4Lf
9ZxlC03GUWAnhgnfJ6NiWNJgQ5IU7hZfMnRB3bSZv3fo44q1vicIlF1bOHbCFvMSjZJaLYTVR5QD
JSVwyQYmW+0/mR/Gs8+p5qDvwynuFmCLHJMa4+4ZoKr+DHSz2chakz2n+S39U3sAxm6Bl6AGDHBz
MAd5jekUjhxb23WpEO42XnlK1g+65yFHWrX54w6cCGq9ZtGL0FlalluwhmJG3S7V767jbVaONxBw
6cXJNykaJLQDAkZfuhX/0BqPLQGPx7F5vBRxkKgDqSG15l5UCmDdUP3zNeG+mpV1NASfAHqzxjfY
/AcMlHnuHJNCLY5BMtLUSgHZCdVqnekj9T2WGbAJJVXoc+8s9VzTn6eosuCxbUhSxEhoxVPzuf9W
QwFZxHPwObe28cMT72FF8sAz7+AMsK/Zdet/mWcugGLkIoZAF32hC6IayFQ/P0dikTBSPjoG9EHQ
gy80v2bLOdn2gdGSW7pr03Pqj1ruJLyCVzI0jNW/hvC0jyrVPZPL2WMXOOG865P8EuhjZF3qd0rZ
mVIbJVGSw4xMz4m1Alytj416sroyUyIGa6F+OIPED/4JQHDCTmoER6qxw43OT2ovl/UPnvC9GqEa
/62M1TpECZDZwLtDepoG2+pUuwleNOA6BXmqM2Cf7OM5JzlUYUzWNpc3th9yMW8HV0QuzVtggpHS
nvK2syZaVnM+V9ouzN4yQAQDZTT7XeVBSG2+9FTvKEPk6PEgA2lf42quZ9umlGZ3Z3zjkeGR1F/c
PEOSlHKTia59ghJGfgIYizz+oQ1EVgsyWiYO3upkAGamK0I0nZVbOYvvbS9He/saw4Iajdct934a
MDkaKj+u2wR+hWEcAg2Gno2cvKo4thToJ8N21u+Z5nIlGvtVKWoULMQ9GLWigDOyS0C/ddxLohJX
XYQg6tl2eeQD7sI7RxJgNnwhS8iJQ5rm0Oph3f3pHLtNP7dkPUBwZWdoaQe150W4gASG1/dnB3jH
/U4oM14rDeT7/xMz/QvCNYS0+9zkEcyATmslDg+pDlyFXjrvByow7rl8V/3cFVr971xp/kxnxR1g
+7n4OeRu8bO/7ymWvHxyewosbLGVITAq/iwm5R4QenOX3FgdO9KU7AmpF7gmlcl+YYnuNdhTDP7A
1v2K/UK5FEd9C/uxSTsXI2UC3FUYI+IuSb/SMtZ+t6SuaDQXS3NN/w1uXS49eRdsi8g660pQjiev
K+hhVMsB6aVqz4+lm2on0YQ27BoBU3b6QpnT6cE2aPIV/tm7D2J3274w205RSgNhI71q/LXx5D7K
x7XVpsWVLXLpnG5hSdGZp1Q9RO3rzNoeuGVkZ6wW9RSO6vg4ymNqFZiC0+AvvI5y/Oj7UHLS5KX2
ogNlIYCzzDXTbG3YvKinXDmviVUp4vuiT3CHSvnfPxwo+mMOHsvuREpt3TZpvgy9ysFaeJIMO84V
WX/KU+Kc5EjTw1T2a3s8JWrXdRpdko1rbfcb3sd1KUEizJ/Y0Oi7855QzyyU75u22rWMDTogEBLz
fp9MC1SJta3wagdJ2/EY1Kpt/kWRqhmg6L5wcfWNh3OIrkp6En7uUJGNscBbKAYJ+0oI8ZECoBjx
9JSlTgMnfNa33pFQofh1dJlOyRxMNFNqo63M+hErWKfE7POHixDfYy9WHaHrpYrNI3Crx0NloxfQ
Eicy403GVQvcgkXRxhmSPXtE3LWnh+WKADhATAGJ2tScmHmdKjve9cbonbN79K27ykmBa0MbRfQM
bN59n0FUJX1jH+A8jdNUk1oDr8HjpnMVkSp5is/WgrhoUFUiycI03TJbhKTD1JexWYObJQpLTpW7
/iw0JcQjFV+2lgrk35aoz3kjQhrpV9Rlpu+/MMWxGLG6kRwHayvbA3fN/z4HzKepHWMIl1+oGwxt
8lhXzFCHUFpTjl7T/SLsSHeBVAVk/BLcsUb8S+PLYh4F2g7dRsWUAasy9WiPSYA44/htx3wIAOiA
gIAQOG0IzCK6KsTP35W3XjpoigqYHccodKRqc1KsFwS6dri+nvOShsIZGpMsxLrmyxkNwUBqIIL6
6emzySXUJLIc/Vz/W2MFQavo3zd8+NC7fT0Nn5lis7HgpyreiuspWr2WEoPMkDcFUknXa0QxllY2
eMEdoZJ7b3MH7ayRX79wTfJNpQlRFmwoNVMvuIIV76fI2B6vuZWr+lzCw5QezNuZUF9ZXu2D+0Ep
aU5di2ainwRCW5RJOV0xGDcW0Waudf1lrBbS2b5VFnnZh3KzhMgeIxK0x7u0sjptogKQVFmWHhWC
4ysVafb/HEJAihu8/T+5pg2+dszfaAasvpezo60kF2e+yvToWdHG4CNdryyclvtbxs5Xlq2ZGm+K
SzUqhMMETcpfdN38LvrWPIUroTYeO5wnn5ksE/htiPNqW2uDGo8NsxuW3bVFocvy5TbykepfAKLS
p0F1cc17BzHZMa7qkbUOaIVcd3tkUW+9qH1FVFcAW+Y98uCCj49Ulin+qIlRjKJFjQv52O2PI9Os
oNdmvEZ9f8ILjBrKwjJql4xuYznW9PNOJr/AnO2B+QrJ/JVSjKjpAQBFg9PJbJZmESBMhM+XKrHl
Yz2b1kr7ujPgCAb9PSu1og3/19EsMpJw5HxxcTWrAWlD9jR27fn+RVeB1ZWfglq9rk6A4fGUh9H7
UHW3hEtj3emDuT1VBptATTgx2J8eQR3k45J0i1tDefTv2zfOvQAyHr8sM4jGLos/UmcSTvKVN8uZ
BCe6wtUWlwf1XiVsSDQqc34/NpH/RbNQiEgLCJywiAy/bU5Tv1TbfIJ90SIYNIotSnJiuGaVKdtH
LhmwXr9WktffqJ7dvMaZb5/FjerOHnkoPRXWpdSeerekUKefan4tWjJwrdYamrZXwgw4+8vMfzQg
Vk2XNGr+D0In3lq+aCaGj4uwzUhJ3Pj61A3gZTaK8dkiDb8b1Oy2D3fDDwICbzKgnFGMWT1PE9ms
Dx6UJ18CCTKtaetsqj8CNAh1mfXWNoENuacAZuFvCBWE5l3O+5/e4OlwHVmGXVZP3z7c83GV+Bwk
aTkMDbvZKBPJKoWEkG6bCxsHPEeRheOhSDEHaFdKBTTOLU1KMcZSw6TGW9JcEwJ7v7SX6mvkGuGY
cb25xzaQ+cPkcIle9TCuSH09CvH9QRRJUwMBLxZT/8pnW7/LkXDYefp+O9RieX42Jl3B1JCKcnex
PTaqcpiNGZMm3qKR0tIm44HjquPYYwyb4h7qH1emRYdDL7KRHnxi2ygqoNSlgNAJ5QGBrcfegVzU
MBYHJbhrufZyNdsCqOuMgI2350fQ6Zp4ZmsJzR5UmCoc5FD5n+eXgTbeuYJQvc7+gZxBj21gqPyL
WQM3vbSmEdJXNsmqjDV8Bn6ye5ICivonFK3PKkVUCKiRdU4Bh5dDIdHRhXaJ3nQbc2b610PF9dvg
rzK8rVhPDDpR1BqrqvtnDsrdbk1jaonUmmX2O4apnvX76dWCiQHRYVOMrRnWuoxoIZEhf0V66cdP
tQkasP+FGYqUNYcPB8QvVIciPJmVAkUZh9KC2PPgyqi+Dt6EvZbCZ3ppQq+f+7veGPIOGXzdS60/
HemHFBmFUZ25j0eUE77IOn9sqVMIvUOZQAPAd0ZHpY6lfY+hv+LTbhG7UysWh4IIHUKCVvoYTGvO
Dag8VTTAiXFdtzel68ItTkUccOgS7Ry21TbYGMizj3fSshJdObjH+r03DUa6/dA8EvWs4mN/WYe2
7s9GDlvBN7hxIT8qCAb+l5riYWYIli9ThLOHvNz8ctV9ceTtAfUtcaTmD6/3m6IMcwIItKISYamR
witZ4sDesejJeWWyroz+DvavY9dTOTPYKbirqWUifTR8zCZSiUlLfjNw7B/8AQ1+npEYYg4RoTre
/SvmsCG5iitlRkJm9l/Et7ad2V/fGzl5HmLD45DO54S/uWKdwMoSve1XVMQCY6q8448/78m/IUbz
tkx4lTNo7Z5QTYyiwXWu0y/Q13PM1rtLglN3tiXwD7KBg/Vh4KbdQezuqTWANN+8czV6Bj3SkE86
CFM9hPJH+fDgsSYtA1AJqU1Kn7ppowQE8SzYNA+zFA5FX6cBoQlJxkh0NfLr44ZzIUCsXoZ3x21J
XGprrNk4HAWkreyyL/dvctki0pdgxCGp8p6QPOx9QXVbwKG2C26TPZDrVCUC0zpDyvxaVg3caLNa
zkF6KZ1Qbh1eJGeQSU1Wk5lOg6sPTDvgWBYjjGg5cq8NBqRcyAmqh0ObXrAQe5l4GZRWxixG8EZY
YjbyMzDYDQ9rA6Bu40hroFQAOdqLLdgWUTNSwXN5ftgb+pJfNAiqUrUullRZLerDsy6ksuDMZZS5
Xa63pCUJBGTmgDZFgEK8wCdIW5Ls97N4iMSKqZy///Y9yH898T0TrAKW6uCeJfmiTMhEwRiBvh9k
CYKMF6D9VsmsJ6O8P4zcNE2Jp3mQ8qr9keIksbB0w4tajjvRfN3Hx7kwOYVZkutQ7pC4JqY6EhyH
zG5Ha2dTNsRs30BPVwKfnm5pscDFAWna10UcocJnfrdT9P6zZUX8/LGX1suVIyDvzUm121PupxGf
PvKwBmrxn1WbWihiisJuRtrK9gMkbLz2JXE7JQVgHBRslu9Pwy1nXCwNhcBbcaS/NVYOVJPkUcb3
ybs65bknJxlVqXcEbrL56AE873kSBKJfcQYx3Z4yQDE+FocfMWqL0MEa2k5iKfWAmmZQb1q80QTJ
diriY00w9XFny0jLu/N/qR4cUKZmwGOA1J3r1Ev9bQkyphpK7DXko0GYe9MfAlmZ4OBrICPMGFqH
RDoVpZOgVzTnFm04G70BPUIx2yAIKCk2cXSljUV5BdHNxFV/5rhRnP+/8mDQ0r6fAD9FD9WCOV52
Qxwnsq4FV77CfKnBB0dvZOFcCGlRglxWM4FTkiEsV6fs83zWiAOh9n0HYRKipRYUNkbHZkXXXqNj
Dm8IV1ZOA+RpBQzmYHVddbEZnG0AyM7jPekhzkWDXzgYSOu2fwxIpVo1D2ZAtdIS54d28SwqltN3
DcyIityN5k34g2Y1HxwXblAr5aA61Ysd6S7uYMkSJ0vQd4bzBVt4m6d5/i6padBRoJPOBtvGoEMI
krPxIsIP0dl3fBfZOJY0NKGYdRz9ixvFPAlokWF3USOZ8pYcjjw2MTdF8H70sX0KpaskYt+XPYTM
szeD/dloG05ec+m3S9yr38PQ/J6buJ7D8K+hzHPuLqVWNeQV+LMwqWjapkuaya3oRlpgXM/UU6dW
RZenUf2CiYqJ2sveWeZWJF+ct9TQNEb0WzkXwwJ+9124qrlLCDogTYAtcQ2YfmDibVEtKfqvjV8r
SVSmd8iYwe0W/8E21K9ymtUet+cpOjkuwWRXEIoCnLNYEGNmlBVYyNPATk5iFC5x92H0PVvrme6Z
NikryR6nvs9bLZYZP5WYxix65Ce64I3X9qGBnt06+RiRC9BU4x/pR+mj7rIqt2cMWJFO2Pg+CB1u
REuoL/Ml1nivZ6GgB88Ip1AV64gErFJLcEUnB5E2kCI6EnLL1kWoUPytw9GDgfTAh1Y8LVZtw7t/
xVTUfhnioNxl+ryJO5DUZNwrDp0jEnpOeTKQgXUddsOOsmF82XeUiUZWZPWd9u8QwmhRa98tVPSo
4HfA6ptDfx1gg342EanDudPKdXuLYr5n/hp2TmebxWaN41e9RzWYemsdsBCqGnmeWETM5kEmK6xl
TdUFb5sjTAEn+sk1fGMKj7q5nLBPzFF8qQxYcKpXksq19kz0ymy9K25jHnROR68Ejq7X/URq8Y4I
Dtt6TL+yY5MF5dNHr2zRh5tzU1KPUZRSwBQ1wx1P2yi3wD5gFKL91Ea2Rh3GtopjV00Zzn6JpM9q
L8eX/8IkG/3eFgRSl79rjcHrFXuFcrrVLxWnDOkIIpFv3lyXHYNsk40yp1ifJTaNic46Nvpbaml5
tlfIPW7VLUxDaOjfpjgBB9LWCR3GcSwSh3e/eWSLiJ5MSHQrYdIm3VCyg6soKZZYeicGXC+Wu11u
Ot128YFxOD+CTuE7kifTq1CGFtIKrmtgUjlVcgeZfck2++WK2hG852zr71qnd5xq9Aj3klkGmaVv
AWqE3CcZ62r97OpbhmQuHbFMRHU9TbwWIiuYZ+Lj4WdPoYleAMFG0i3oAWScqZM40srwMGsBpChM
PSgcSF9JfVFbaftgZEdQcacYP40m6umpUsgPTRU0i5mAtbPxmcIoyUYSLZyCBF1Y/lI09WWy8Tol
apET9ONlaz2qy7y4lXlR1s+rft5nxKPlt15IQiZipQQ7nsQTiEmWOcXPde2CECPlVtyv4QyBHXn/
NkQ7ZqS44cikGbk5t6vgKyI4wIjbfzvAMNAas5++Y5/081/q+yDqKHLFyfuGsNJQKsfhSxd85p1z
bOiHaFC4VSUwOgrzgaORpiQU/dOYUauvn9dEVY2cGNpNiJ5BHcc6cyPg3OOWpRR7YcaupFtlQ6Ip
XCEbn4Z9qozNG1zisE3ZeCbodFqjRblOQw04ZaIRAXNe2mOfLbyNWflPzAR/SVJDHjdmF+s0xjqF
qS90BH2AG+1DTiParUoSZpW0sdAdo8vApuO6AxutmvYzpDHh1gn4Ap6UXdT34MKKwUwfV2L1jvH4
6OSNVxHEzTUnB4cUDyY3TrOoWUd56UGk+C5G80PE+1ZCLl7lXhBjI4zKMW0j2qUxgGnrWihw46zy
+CeA4DaM+SLRoPRn+6hhEfxKLYKIuZaFxggCk8gze8QHDyX50ZZgnEvZoW27Q0gzLWCetrYY3dfz
19dh8ssM2lTFixrK2tIIr+rAGfs6dyRryxf/v9fW8uPmJ/rX4b2O+GJ8JX3fzs5BUnDm60RfHeCI
3EYdXJuyTg3p4UO3xhK0iFIqsIFawv1R32jQTQrxj7OhLbVHQLEP233TBbNPYvKgpC1WCl5UhS7W
qapxxDxTamHgYNyE0jVCisormSVqOZmpStzlu3OqRnjoxU7vEQVPCnRK9i9TghTRnn0NFpUKpS8N
EbZ0tVGl4ZyRh4mTQwHlIxPpsTGflkHZKiuyOXam7wUhXSsZTE/YZqTyE3y0DNOW45EFSEgMz1BU
+e7YlthhSnZ99q+13MUytxD+QDSy5idF+Vy6jJJFYTk6BYLBA9KE385+HEfFrNKjAqJC/gzZ88Kf
wZKYTS6SGBwYDrtP04pEk7QaffhLeYe376L8HFHcvw1KMH2/Cwa1hgdea1zKFu+A98mQ7H5k5zai
15CL+xv0MQCaqAyjRC/ErCvDoeTHNOr2urFyYyLfzozha2tCRsX2uuGK1lsf6kAXpiGEWIaFwriP
jBaeePgg1XqrZzYpY1O9oZiFIFZ3VKEZR8N8JjW6FzG+evvJPNa4q5Kvl/Aho0dRfF/M6WReCvBC
S+vV0YWS0xHc4Fq6f9/xcQvmynp3xmUJv0+zYts1G/WV0RL5WKIG0kc9m9k3/pCXHo+GeZ7Ge7/X
wDWnhSFTJ+PUX0TUxvtc8vTGqRKb+6WP6iQOYsFaQQsayJUdTD6UWb71j+abCsd2pCm3ijWcFdZP
171zq+iufFcEdwC1WieGCCnBy5HKDnzUp6S2Hp3LA/GgJY5DrH70pxhvSm6LQKeFT80DKJTlXG5E
sdK1lbuPHyY6SmvGvXEgH4MGV4O8HuAwAvKYfoGlwiAEI6Ce7oJpcc6GWwWVDYzs//lf77RO3Y7s
T/6SOh7TGAf1DGYyEecxMJumj48c5PBH8UxsmQpK4iHZr0Jx1aXItgAAeVcVLqJEU3K1+IVtOcVR
9y2CvUlQGZbK+gmXk5zhULd7WJQhhth7vZvYTXqZxRi0IdVok+eRTvGiGGTr0d9e+tM8e8sKC5M0
y81fGGLSBqvUxIM4W99lXAK3Vkw1yhiHAl01Zzbu3B3556X/S7dPnJDZLI9UKNhDJru5EI0tDkWx
uxez2fgwN2xhThbzG7U52ju2X+SopImfkBY/zQiR1xJq582Mi2BWVLcIY5Jq570lQnWfd4OYdDoG
MepqnR0GN4nK/hr9JKgwUCRlaJK8rs7OzZWtQSPBY2qF4G4CdkXQWFGIRml5otK2tgUBp9Pth4md
g7ZTuXLkcjIe8JfZX/nVpZ2rw8Kfnw6U6NVlGxQsc/sUmu4+7tHQmiJ1idzHEYwhNAZA7qi23Vie
A63TDXHfofSSt+kx1C+vamX1g5n9l9eN63jCLVj1aZ2CvRE+2Wmex5Me2tFj1B1TR+rg95gG4PA7
7mSSxQoEF5IiZ1ZLmx3zbKMZWmSYDgWm/i7KyHlOv+pZkUUQdAGJWeaJqsZisHpxRSzn74PzZURz
sPV6sTETY1oWs3BibUfLAJ/IrXDju64gcCurATBpDMBCNHDnlSPoh5IM3qnZ09Ira8VreR4sqJuE
K3B63jzuXCb6l5thnF6meWv3HX7L0gTSWKGueLSCthRplI41OLKngJSYxeYqFae5akDSasUfgyq/
kbjL/HFQq/s4H9ol0vLYjIvs7cJukGbgl/KlUB/FXpGcR9pNbBJcZnse/Wsu1D/z3SgKUFkJcp+w
ieWZaGM2+Wpt8kNzoHDfmPZxVxJ8bM1pX32zLgo8yTPD14OI1BdYEnMOypme7LCSkMnLGJfhGgxx
TyuTVpYBjP32BFMu1hV7gQ2U3MuyYj/EDAwcjOoAHZPpSF2K0RKM14e8cpPJtHk4NYvbYcA0xBE0
8yIAPUgHYfH9dcXMQ2pgk25BwXygsM/LZ+I+2U+Msxu1wA72dz89I7o1aLXUGX3UQyMaGvTx7kFl
Fu1xc3nfeyfmAYKHlBvnuZLSP31FJp8KS0D10xIKNghrAcSW9+B5PkXqRfRX9MIlymzwLgQKVkAh
orSCLF69dGgk8BDxLnD7mf37NmKV+D5qayeiUOkzjYYjgxu6A6xLHCSnQcYYZlufX6c4uIZQ0kS0
deFuomwDVw23XC0Bwp2JMEINRzkxieNejd7wjH+dN9iQEgjpiPrDjGY0aYD3ca1HnpqkEd2p051T
z418EMpJ7qOXC4p8ajU0/D+f99geQPyW+Ne9OOhljvfWeF7FblzyVsDgxzD9OwBBCMTKE0nuIXS9
FE8ver8Soaj7FtiSu+yS23zWleCZ0Ti17TIay3EbUD1oKkTuW3EgwC8WEV7omwqLmep98Homq1zX
jGYvpDgheQE5IJ8M6GOOmzSGA8VK9yednchlDD3KcGfoOUTaPFOqQZUpVv2ezcfRgLXI5a3fnD5f
bbSujtViS+quqi/2sqFQ+NTZwuHovHmJ56Ptv4fNk8X+Cfit7Qyi5U8F7p/f+rCyVu+y3r8oOKMU
OCXtQqPIRSvzgKHhBXZZxNwuWZ87wiZuc2m7XoSKxJ8E6S/PGpjRqC0Y0tCiQcqMp6LACVPWtGuS
tjo+TSD9UerqyAuUxjEEE8zOOV94b3y5Cd69qvrTslCkgjP16IzSm5MDfAMB34QWpUkS9nfEWJe3
d/TKyDj+uljhPDF0L9f7dFAid/cV7eumTOGxi4NduM/Hbos8PMoK/3aY7K2PHevkz8SaDH51WNr8
8djxoE4uSsVCcigm9bOedC7kbx8enmoaIVDERi7EIPKOwpWGgjViGGJpwKaYz4enKuts7MZl381x
mqjoRwz/DtexLnAnFfA7GkkQ5k6p34G03vIRH6GprWx2YF/rh2I7h9XvqGqaI8obVR8Wu8gbO60X
NAOn/y7hHbcMk/0wXRfTQnkJs+ReYPqK/9MEU8z42tJEJ72HDL9mttoYThHdrIiFBjLUR9IqyrVC
APXpQQJPL4Jf6kb48agkMpnXmpu3mhLqtwtEZ/3jJaOpWONqZYFnE0eLQgKA6yFTBA590hOd/09y
zt7n9fKKHiC+ZBQbEjoEZaudVQzZi4Kj5af+Fp/nTX94PWlqHZTIWJQ51Q+NdzeNuzKxNHwMJOEF
efjqfi5BUF/LM+TGaP1moy7Ujzp3bya7CTKqHy0+A9GG9Vh5/GH8KSsDEEx1sLafAuVyI7jfssb7
J7LseURnt/Xe0AeaGH6ZsbtjmPtb8ff34dXMkWJjEj7MIbOykHFpoO08SYRBzH4TfRYDkkN0ya3E
DBNDCJyKmACRzi5k25sqtMAO4NqpG0onGZwt8qFMRCa2ugENgQAU/Nyk+Bue+XhUR7DsUKPnvv/g
oUd/2OLk303ejXehWitvss3xxAAcvbz8VdNAqaUXTmt9UxzmovIUbN/2USrwQXhMdj2nn1Hlq4ef
zNEze/4kdHgN5rAjDViZ4J2NyOGgEw37rHrRyjxC+POAw3d2aubw1PT8q4NAoogvkBD1En+V5Eq2
f4YCcbo3OCvxzTTYcFmeFUFFMiFonONn0PVHwOHBXpcDcRKfwbxQKpz+zakMEDs/hajl7BtiuR8n
99w71CB6VoTCtFCczVc5qqPL4ZxHi+6VwUVgNSm43EwutJTJxBQ/A3HF+F8+89MRoWZyCXXmeGfG
3KSLZ2vIGb+R49j258R9s5nYE1Vt8/OFTMlk1YNr/lUjekIroZxaIFmSP6NiSjTqMLeEJS6hoY84
IWOg8Ig+ntQar4+abkQvwTPWv8K23n7gPcER9xaCwiXyXyN7t3YyXpqQbJaHY/mefdTQPUyUENZh
BXjVv028hAa7cpBcLVMnbWWhVAOnVeQTuzU17WujWM6RqW3EktvGeEwSicRryTcDKfs/p+o7Ctx7
/CI4jQzsSlvCI8k/m8T/TtV6TcdNSjy/614JzbkpZCDSlU8+fHUKqitrdf4Jm2O2Mko5wDGFLFAN
XvSNBksxbTIcexSasA+sUa1GwnNgcdCmEPg+AiFnDmV4qLQSYgsRJVL0Q0k2gaHi5210nP0OpIh1
/9hSXlc8ftk7wzeVpHHH3rIhoWgiRzn3Mh1NE7HFK1FiG82pdmWZj7VyGi3qraob6PNn9QEu0vLX
/c/6lvwVlLWGgCC+yOlumf5jVCxAkQcIrN1ODAxLwWAvMfEr54N/h0YV2njVRFK5dAIzaQHwwtQP
O1JGa3rr7AbkrNfXUHuZ1sCTc9PmxxMHPzg86SOvcSmda8PdgQzwQdHzqtfJgA3OtqvBkWJqQYfY
YYPMl42XmaFM6UEogIkMf/ZFNgFCfLAlHFNR3dAcSeoV4W4v1xQGsERJ6rvx02ilIy86T9UBIZB0
VQQuYfaPgg3pYBn6NpBvwg21Y5tHrw1FY6NQ34Ov1WRdEDqraiusnPJwNTSTw0cEj0FhoNQC7tY7
BCzagkLANpN7w9didKR2sHBPttIYEeovyphuanLSLxWCBz/+uM0kDPHu5O8Obq/YIgUlIzkeNvlr
UESkN2a4EJZv+yiXTyIxwxcW7UvZkQb8bPxRjMCWrV4JzNWlbb8NmwxZZaFpyIbCN8FARte6lTxd
6P042f8z2KKUcvdnK7zFZHHAI8Q+q5k3bFOgaobzyPsfYsPb3mUSgwDVYrBJMr6n+M//Ypn7Pjf7
ghfVHcbRA1hV6z0vFoEDIMlIrOLAywKzPQcwgYSUqlTx4B30WURBjPszi4n4C2035T8zmp9VLUfl
UZhvxhNnQFD6c0TUR6o27HsxsGsxYdBpy8WcE5Vc9kDlbXduljm1DfWLZj2V6pLp4Binl7FdhMDQ
QvQ5jRZPmmIDj+LT4q075oKM/G4dl03GaoaFuZmPuYyt+HqCEHoTFMfH3WXeT3CfU5ATS+lwKKHk
nMmsThC+Mp2HKm6PChlBTZQc79DiO2eIqM44SNtev35WqvmxGG8xm3WiBeWj1PuvOQzYGOSGXiqb
c6WnBTDdvCKrcKhBvi9ArC4aaqeItNA9omQUzyidNmhnZ9oYsUNtcUjGHGowT/Hd3vm46GmpTI1G
7+oiOpbsk8IM9ct99Df8eHuUJU1l6x0wA3In8oTWfjalpn5z/Eac0+ThE8DdWKOAyF6g1JSTD8kq
SCCwPsH4YD3ph+KuN+fxICvgeRED8D3HtzR8vaFy15MbY1JeK+VIWiRcINE2xpjNAkhTBqyMO/BX
/QEol5VFHI6UeAkm0pnQNATK/FZcc6gZyS46hZ1NJybfvIhpepYMk6Gh7+qpFCoQl+uGvGde3uth
aonH7PAeNxJNvCKQpHmAjaYKsTGKDCpcdYimFl0sDeeePXdOXXQVyDIYocCfWaWmSR5AStMXSpo9
wmIVxy3BLu34O0teZgS6UhXkpPbSjyL9pKYKgJTo3+8ORhbbMT/jvhCUbVD9JKb1/R87ItEogAiw
LSE/7z3XRIIOsijbrdBS9jaI4BtVzrzt/qZWgW6Bhsh2zLn/omfCLE+LHxwP6Fmr9+e5Ukq7BkRY
bew9F/A7pkYMmK9tQH+VEdR7zZ6OBP5TQ4pk/17xYcgANNeQ7ickeiboTbbyWofHixLpoNWUKG+4
nAqy+Nedz96gbEbhxWt109MGwVv3L1L2Z9peRXh6s3Ba7gP3hQ3cT7Usn2f3uX65+KIkLUjYtZIf
6OxiRzV+ISGYdbhX+2XjfZ9AyAMRXY5pfXUuwNrhbhDf15Ub6hN4k4amNKKVn3+Q7U2UOot3xRYd
cBRLIKtJzWNiDqivVHnPbH5egYZn1zvRHfp2/kwC3UukN3i2NcawI6MqRac1YWSt49M/c0xsj6K2
2/x1vGq8Z6MfMyVgIVwGc4CbdSGtUgaI471La88qY3UnlqeFnacM5dpoml9iUEGcXXLz5BK9fpaH
wu5JiiENbuHCgMMqhR/jMa+TOGKBOjxxAg5hiRi2oe6LNfHYZwpS1fVrLjMABqr0VS59BwpPtw/5
D2g8IJ3k6YbkwYUJMWxGJmPwWmyBWI54dP/25r/sFSDpyN6CmeScIUW37zRkXnJ88V27asEI6CI7
O8XYgg0/pinaRxGLvN/us7YGA3izLrZMQGsBREQNCqhQLjhv7JXnPcMM9zP34hwR5pTwdin6NkoP
zGxlntx4WdvCi6/BBiT+lX5DmyXBs+fLmiVMoLnnyA5CJvhaay6OYCq+gIcYb9AT3o4mXa4gGfKI
U+hynV96+/yPmApDMjcYGaNc+lP9rO3Dt/61hP5polAasnbeW5udU0A6ww1CUvX5lDSKIN2kEBXc
TBhdEyLWdabjVheQhyATL1yqIZBGiLs+AFgVlTOebxBt8oY/UoJ5Ph9R96nFZ5yoc09wo62A2A2u
XzT9BydT+WbhOiBjV0SLk522uSxTLkjNM0juBOqYeZod5zCvaD6zQ4hBR6b55KJyy/RXbpZVFhs4
1e3CGnBQ4e5VGOnRCrKsdY9+hAL5FtVUhpCJ8OjvQGzrgXDXFRld3Bzz60FM8Z9VVwpEyMvAq0bh
txkn2l8MRRNiP1f8nlJoTGOVuOi3kVYcFJ451w/IUOkR9yKnojlankq8pvuN32aRtH4WSMJz/MVh
S/iLnF8BbqmTFpkJhuUQym9s8mcavmZ/p1MJWwJ04K1aOKOlaB8/D8sT6LrRuINTocYyW44hnoAi
u4C8Ps7z7OCunKJdfZtYTU3JvCOKGzof7BUOWrbYYytXJgrTtjA0Dfp/Yp67e1pJt8zG8P9hPi6T
PZPBe/owjuIyTWfMtr2ZGqWHICamICnODvn1Rf7Gs5/QjpFxWOIEPDEGVz3+VDclFjZreENQorX1
K2JrVak2yDV23C4Uf1M+7DVZjs4kYU9O/ei4jlh2uy9tmb9wtElLMV9IP5+D8pPEo+mgyddyx0N3
38PcXpFfXXR5IvinUJLV9KWnXpI9bdHG1XQJJWndG9vpRi/PY9BEl18CArN4WSgF4sYPy+KAEipx
6LvCo3xeFV2qt4LzRONtxk37h4csNHtioZ0vfaDl+ll1/BfQ3JP0Uv/8diDSH0noLCL4ykmFu+vq
FlAotrOaZRm5pc4NpuJiS7Uu+edj4yKqeSUXyBXAxABodRCMl0OlKnMFIvYoRKjOUPx64bn8BLyZ
dsJsr3/N8K+GABqI9doRtG/Zm5FVL+nG7F4u3ZbB+X3rVxu490EOKwZxqR39x9XRkQrbPL8iR/e1
rBPcBcYisEDlYbuI/Ha0jbAB4p3f0vtBL1DJw6EJ80Jj9eA/Kz2NVDwuVMiKQheQdNhK3N+coiGq
ZUBs4FzU3tdsmOQ06mOrme5rqDOAS2I5n/EPN7IzHenfaK/PSZfAaXM2p0Vttk/sgsUTirLGLgIK
b28/bcOJmtZ8EovxT/L3xmhW+WItnAA34tH1frno7ul6KVLPgmJOtcrlYsitECTe7QOY4stxSyIW
ksQdyP6Qhw0cFSUCrr2VECSOcR5R8QA4fUdnPR0p6zl4cK7wNcdMgTIk5zoc1yZkG7CeevaguP7B
fFd2WDwHQp11UZdYI9CdFVIwWptuav776PI5Bqd6WzyQlTmZ9FHdcw2bOCjtfehxWaYzKZ2nPqI/
RHAb87IyKPeOQx1slJ8+IwfqzCyGokPiImo15ynFSjIsshl6zlLBSMPJ3Db+5FMPT+XAxIxqQBn/
ty2wKS4rutpD0ypcMBLNSUPXeeCOfYs/aILS4naI9Jh4mP68NKuxp6hrS89Zy0gHWjDGF7QnTrOr
uZVsQmd4888eQDKVASuRks2bpYp0+gdWv+8C/vDJPCCNXyBkQ0N/Y5rUXDxocuhs7JiP9Qu2MyIF
o8i4hbW3KlHNvN0hEgEuksDD137gfRt+rcvXAIbY/uDI28tY8+wjtw3q1o1DsCkmCA23CAil1hso
U+F5X4pA1g3RxA4EalHVcOLG0QzuhKIWsqEGpilpA5ABqG/r5VL+NMYldTxdRNiPl4TjstgnKPv3
D49yaEd3YZ+n5KWFHnxJz4IcyA6tnPU96JhT1BZA5MXAGXFlRCx7gnuvxVibEJKCEV6XZZWQ/O0C
7r3OF48G+xru4Vn/nYIGlAhiwxjsFZrjwV46dMES6buf+GRhWv1uro6iGTTp3vkPdPCQkgUFLJ1k
JN/txBbXaEW4z2Olzrujf9lAJgE8LmZHOxlhrzs6HTb0EgrnDAlY6ozhC+j3IzS1IP6+yXh+1+Oa
6JlCldFv9CpCPbLxSK5MBFAw06DIXHfkfBSC521CgbDAxZW9em61NGek/R6PmX8sJqA9DsKeMohB
BppEQGbwbdwp4fCIIdKC7Rv7VXXq6aukAcwi75ubBfNEXlo2wjWIYx/lgje4Tw1W49dIkSk4/A8Y
tH+p6AXwGOg3I8YpxFcEzUVqhw6Q+cwAv7h76560C6lBHIJOywseTl5sfnNCSEJTETtL18hPupAj
BpX8LhX6alUFuX6FkRQuWQ4yedNF/DQiY27pjzp18mh9hRdbUfrP3AaVDYVSOt8fTu9mTci7MxaK
o3Uf7iCEl8itil8oc142yEddLKUxmdDJMEtyIGTefsFpQ+BK5qRTaakNv1NopaXUCN8iTAfPYkjx
1wwHmjNr6+CM6sUbku+9nrnYE+ZTWKYpmk6hv7n1T+GN80l1gdRASEqhaZzvUpWc+w2ESpXyuitp
jjJM5WjODeVvKmHGuPCCm4HfSHvlOgjgXH+ML6+oLUQ/nlJEQTyHCBkGBb3hOAw1sZm/JepdutB5
XmVL96R4vpkK1fEyTrX6GfHyVdV0g38AIl6lSjMuLiKI94K5RojJWQ79C7r9fCq/g/Nti1aV3vxP
VjmUBnWF16NezshF0SQgHzT0MbKEMdKxNdFt6I5FaOvbAYU0jQWfMLSEQxQhQVJ0Y7GIQ3JwiLyq
2ofeKHP5RVeRjdkU7enfbMbBui2t4fhylSYyw2Eonje9ns5yW82fnP+mG7C8yr/hzdIZ3tb1bRCj
nEdTwuBJS8FIDj/wMnoObIlHW8XPp+j5VBAfAt2khoCcIh8OEMaaXayTJyjckK/73bmhQZh++mTB
AbxPufZGg77/vlmcS5z0kRxk6KX7ZNuJUF+W2ybov6OuBoE+NOWiEDWDkbu6fNVOh6WugVletTtD
rMsl6Iy+fJJHvoyJxLNBYuIDQPLK4oN8mjIQflhDGYvp6hut4qIMm3JGt8GbDA3bKCingTY+F37U
sxyVL+EKGonrmf1RSKUrd7PshPn/x1iqtdb/AuwaXY9faAd9JfeDzaj3aoYGi0lLPHOUojBbrGhH
7hBBHi7LrpdAsGr04J1tjTCwIbTBCTM1YpPrmFW37Q9Whs4MDgUwRKUsTmkP4B3qQZJC847V+CFR
LYjFRtabBQVr89cf8FbzWurdjQbv2GMNrRhR9D5Z+GL77CYCrN1o11zlrUKKBL9DH2ZlBw3XZf3G
AILen0Ha70ITN1CJC/hreJUs2OM81RDT9bfwo1EanPswimP9jR113jnyISf9XNT6CtR3nrnwcRmQ
P+shoPi4oXjnaBdJcoBnKJ68zUfGFd6D4U8uLH3UasSAzuZOpyca7j07HiefLf0d1um5olM58k5x
khDjAoPBsemznOlm2X43v4V56qPHWzVC2wGKsggfSITXd5e1z663JnWgNHW8/DnmmSdy9maXrHVV
aDqqgVsWdYI1H0GK3LFTMqfQZ6aGm+K54XK5T6tI2Py0Mn2FJjTKw/VAWDY3LgSKf+cZpgvIrydu
n5Hzo/WYQqhElcbYStCys5CiuStQau4hrUOQmWuKAEd1mbRcro+s/H1/WB62IuP63ycQ84mLtWwW
8CVOcKyJgHSaI1BWJNyRrX3MZ6FhCKDUW1kD2Ojm73mPmYWXHaac5cTzplH0Qib+W8zFjSC49+ws
GxFV1jjjY1NMGJzV4YVa7/6b2j0mILZ/nM1p2yFPmiMSN1+M942pNP3B4JkLzfNCowd0kHnwVp2H
6FqpS2XHBF0pmsyXZWD18qInCw80REx/w9oRl/m4Vjhy37ul7Xl9oZ46eT1IdeKyIAaycE0cpiyX
6ChJhvs+mkLkdU69HfxDV6KJQNb+oZXaB5Z5DvPASJDS9fsypFrZCLkLeIqgHBafK7b5DHDIMy8b
LzQ7DJwt1MmjSQ+YlKg+krkNfsQDaIp14+hahbvN/fENzQsiX43wqqW0Tg1IO70GdHGVe9JkBXAC
HKex+NQ5vv45jGTc2l8zhknOZ/y/JzbetDYzTbRANtTO4wPZELRhAlnMlCZS8LgNXvqh8lKhh/eU
185871h1MyM/UtLXC6GSg1SdF04woE5xW06P+09XDvOAnE8rRgOHQNb88YmGbsPjIdVNZEWQIit3
oD3cqTBEl9wtiaJk+bYVuw0Ra40bZ80K6Mp1D3B6bAaZ9kfuN0w+I+hMlyuIBrMHx1blsUp+Pd3v
Je9CUvfVebwaTKhbYbejYtw5e9yH+vUaqLIja/X0C18YIXu9Il87JHUMSAjFP6TonkkSUsrE/n6n
zbs57tW2U/W5rXc/rNMA4XVzrP5p9xMm2l6/GW0FBkPCLRqv86s7geeVciyyG+xJjecelrZavsWE
P2tbzN575LiQuLmA757cZLJkwozXVGeVmBicvHWx3AxsQawwCjrqBOvBJwk6IOBD2Atod5Al0R/o
F2U1pxouyZwoxHYBvYkKO+FmozAlhyA/mccPFDaEe44oMe5BFX2mDJT0F160x6OsbOFU6rIkbV/7
BNsB3NH2EBZQSN2nLnwlCx7RYw4efM8cQa0vb6JtIHZh1NlllI4QFXZ2440QOjfrBsyF1AcRu+ag
wbPvfVMsed+JMV/KDiYoJZawEuHoysRhkPjdDgynUQSJuTWSyrio3zRPzcm89oKViI3V54WjRsdL
97jm3RG+puWuPP6kBFSr61WlQ5SfXhXWNS12HwTTh8Iz8q6TKOdXhl99v6FySiuzSYmCCznm4q3u
aXLew4ekacrxGoxKWuRu5EHQsv/lJKutlHEdjh0l+InMnkfouWkPGDiou2BaMB8d75rWbVvGBxcS
S+M0sgyitKUlr6o61ntEZsvnVKLqnjPxb6gTXFgbezCZMKqtrdhICMJnVty1sPUHT2svyQgorZ0g
CjkHUfnl7g8xLEni4zpbWSd0YlohlLbwAuoWYb1KJE8rmAZFy+25fsBdPSr+naNWbGGbWhYABACF
tUym/MgFsi9yjXOlwyDXPmpnRrvqtLi608xHiAnn0tfXoXv8pLiLl0VagB8BozusNTT2X1Jdwj52
Z5SaqmwjKw/oSBJ3YH9Wiks87hZew4wM0BopbUSHgo31W/L3Grp+zzr73Jd5lbhYil3MQURSGQGc
/+n4Flq7CkleQNNwx7OKpkLKmVClkpBqs7nAWhqtEzCeNTHIkxiGA1pb5+Wk26G+skYykD30vEZT
JVpb6uBvbeoxnWqsM4rSe22u5QoHmhPrqek68VAwU/rucw7WfizGSGLr3UORjW5eR/euvYWg7xCg
5HcZHfzPaRNPbvFBhIQf9G9xwrrQS5XR/OUcCXhV8e35UW0fEWrT8hC0hHMl4AC86EIn5FN50H8X
caKw8ZPL2rFGx2tdJg5i1nHbg2+4cyMU99t9YJ7ob/6Ls7h2V5M0BHHAW6iBaAVGYREXxs5MPfl+
zqIl6ujhuTn5rSrixZOOoXXmM9kt2HvNzM+oUk9wt8PPfLNepkB8YjZ/OsqsFerQ+thQXtJAJsY6
YYUZUrN+sj9AKRDbPXhWOQbTHj6lXUbtxtNeH0m46EKzRlCbPc+ocXPsuHQk5172b7Hd4NVkHQc3
L6jsmtcCjVUGce8OvTXCYpz9clyV2mQBibfM/d1ipiXxO6HAWlbWvhZKVDeGXi4GvspkLY5fiucy
gTtVNf+5OnRTznBmiyrb72HivLgeW46PUMjxu2wzCRwvJgR2WewwSK9lfjTUJvZ0Ayz3ZsGBgMt4
zNd9DUs1AoctsOKRpK4vNOhZjcp6hopQRV+2ClidZNgpCYbtD3kLADUXY18r6Vdv43ZCMsAvqYAx
jKHbOlSKFGHBnYGjbZrlKLk6ZtHDaipL1KpaE8vBWQuTtvk98CirJBYItdh/xWgEGReD9efN8hSY
9gDkY61EaQrkC7jJxdNTvMjXsyqxdl+zt/4eo6JamvU218A3QMIbO7NtAOP1A6mGUkm7EYYOzxSg
7I1HtSCNVwhThME7QBE/jFQhQFSJxboXJedZlDgb1ngiBTlCUqi4+Bow4QTkphkRqJvupFmciTd4
AblWw0B7HZIyQ1t4tgTRE39gXuWSK8eja2ix12TkffXKJLNeW1p6f40l9q53ZM/lOCG//IEqVIfo
cMBWQsX6eByqXenuxnzkVE05qSQKntoVdIjMvRVc3bYBO7PKaWQzMZ5YIA0nJXedC3G/jICh1pBn
CxYPbKshO5kBEYMPNo/r5r0KrlGGd8TuqWw61dhzlON9gIUD+OKcQ8EhJoofZsXyra6VKHUMMUNv
NfQGgRUZK7AnsCck40Fn+Y2d3QZU2/OxSvZ2w5CHwLJd1jRphCzQiFwuklyiGxjsT5tjmBZPVump
E2UmTlQBdu20r/jNvZtbTg8udMLS4c2t8YYDnPhmwzemXj7gEfSnQGFHPif0GRdxtxgGmLTWOYPP
R/QrTdwsQZ0MQ0mYPMPSHPYEDfoW6zyvHNj7qO0Ipo0n3vY/f6uiPriI2awp1Osmo/OHyXJ3zvIF
4YvxcfczKIefpgZty49uidkMLLLNVY6pQYCcNmDFGx/WFh3mKaJay+bpysKbCKB/Q8TRfNqXbQd/
y9sYxEl18tfiTnv033VRJcK/6XzACWiP1Sz49QSVCBNPvhKZlIW7c4MDpYj14zUvYSqPy0NT9r0q
OhZ6gj0hAIwRxcMVQlznkDMA9gT8ZIJzB6XpHoZh8XkFwhzgL9Agvu9ruKI3BHYxEaqieabLkMJ6
TeMiv4NLsOpH6Us0r+0HtvHf+ztNGzYUWhTeZ3pto+1K6YPDAHsZyzXASezdei4q73CoKcJz56p0
diIqIA8hKEIx6/MorEzAP9VkXRzyDtrD1q5E6RqVdT+Tm9iZBGd4BegVcN7mGMRUbJT/b/z3rUe/
t8/VIR5tWmDNfoP8uKe11FL3lA6XDzM6bd5uaOpbAgv7y3I2vA2oqvcSVDpWPPvEgTVpOBvAEHor
UpfRa48Xf3hn8pUryBG1Wia+Y8hEy+TCyBNJw1KmHISt9cNXocTQ2PYEyBb1D1+YcpFMJDiiFIP8
JfGNMFuCFv6HpOPfa2WcoBaHgkBVKd1OF8s2FcglIkNpU7ww3El+V26OzCf4dO6t15g0dlU5oaoG
2pHruiJ3UNszHhDT6w8o1lTlzpNATexRjOO+inJTicOno+F1SJP+yDiQZ2HeWQ3wvGKOO/GFii9F
mskpLs1XTQ1ZjPnqvJ5t0aTAPZSfBvDGHmWsSw8wFFzCdHC13CSN3Q/lwasWvn8lmdYwyDzyz/Zh
71VKhppX01nIB9D4d58taFSvcghNH/Dp/xZtG79P3vWMNXYqScDe4ds45lT1vtu2Cyt75/bqamXj
/etRbQ6rX7nfCNL/IMDCS4xoTATBdD80BOmqL8J5edftaE/yC3PbzeNMCV6eCDlAZ1h+qXaGwqQc
sjYVcNKn8GJ46lmkM00YzOrIAYKlgoxlwV5ASFyiikLDF6uS5C9A/PLQi00+TYUqgtlvNTut/hyf
262Ipf1gtZBlAEQRHiwm31Ac1nrkXg+H7PmCsI9beH6hlz139a8EaB63sFDHJWj+waTBPy0BWnhK
fRDA1qpPsVXxg4rzmJq3PU6p+7vaMpSY8JojwTlUhy5pDAywCDW2YkFbUIQ+KEtN1RAmjTySwe1o
jqZhk+KK8m5lzAfUsdeenNj9czv6XEh38sGrmo0kXwtJ176FUv13mjU7DhtC/R+FJX0zfhWzjjVD
jf6qJnu53wMQvkCsViEZtdwDDrQmNX7nsikKJi4PfZhUYpTk3WYfYAIEFwoF8XTEfH9LHipVV6c/
jsVEGMxfXPpxeZO/V1UqxMknSoQXNkOrldb8ZvALWJlZxY2qRQ/TeG4VPZYsgpiDF2sG5C84EWlG
Nz6N+j9QwId3b1TAfiFuDVmR5TnLCWgtPxBZn5dLAErYZ0sG7PVVZ0EnmUBI1AiY3H9S4nc0P8gq
wAjrF1fk+fTYCJHOiadm7obHf6iEV2NEg1GlZpQ1kBMdAZN0/f1RsChiuIAZMgqwGqicdGaQtyk0
xIRQkrZeTmsUuOcQoiuNV9J4/f1Fzw1+IhbFdOjqvzFOc2GFIwNGcrPl2hs7qIrb6jjMQwqSQpxH
Xn1BUdt+R83OnnrDoZ282sM5w0LBG7J6IPN++gS6dKIoBp0ehQRnQlVuheoyJ9RpyofHwWv6oDCF
exGdEEEHmmIO5Xy6cJufuheR07yR8i/Ve2vPp3oyvXTq+B/3csTOJznT29VbU7yF6Y/vC1saOF21
GInqZqHyJlhDqsMdCPXCVaqJabiYG7qPs6gliI16bYnul54Ib5qfPRbr3iVB3rH/GGMzOCA+uT2y
yFV/rZJbqqhQE3mg6e7PYgrVI69Ml7/YfrpS94wYcibgmVJqR/aepTcMaksDMyqxF1+OZ02etu3F
XufZVmGYRliQDWL9cGCq0ABViiE1GRReF39p2K/m+p7viULGOWrqPfSUMcmK5Pq5g389FyLfWO8P
6A26CfWFnMzNmsov8y+GvnY3XorrT+/2uIq9VH7QwqLDUJkK/kWDDyUWbAzZzzG2iEeLDPCs+yTT
1uYMCMmjQBlv5cw55+LIQpRFd92zQ/nqU0Emi+7mds36s+r857TDbWJcHj8iO2UAkmPQ/ZjScm/X
Mr8ApQntLoxbmXDNZ2J2PuO/ifA21qYSrIWvoie460ip/xivD9AJJcFrwI5TksvXgEFstNIKV/Br
5O4tlbTDACJnRQVcrwyRBwdNuXhUbv1XMdOzxAr17loeS4j7bwyRK55u0IuCHKji0JLPhYD3CA1I
yjTWoUvmO+TxOSTR8jWhJqXFruX+T9f7XWC3WhDg9qrJRY+6CkqeCX+oAa2vjq4ELKTB3HVn9UZN
J3OFc4fa2dDDc1L23qrUHmWn9k/fvFID+CB4en3CWEAmYp+115PnlHqUPTmx/xFGxZEjBiZk3zFm
LbhvKEX3q9LgfhAbdg45MXyUUV7YzdnGk36bNGGR/TUMrDmNh3kLWBuiTVUW6j9nb13+RuKYv8l9
u3UZi9RWdu7qxRvY9ymhxF1oHLHfJUPBjnyoX94wq2T7J+kw19PL4QofEOtsqAGmB6mUhhYBO+ek
0tX/nfmUqFIufgC7JIyAO1fjQ60o9ozKcBapkpZG8vN1JAqj1zdCSOfXqRAMxyaTftXfD+hgb2e5
lCz5QOs9UOnU1tIAJKFGjfa4PgfdVq1iFZ/rXTfmiCINTysejg4Sr7KmntMkeSbcKWzt8ZM5e1+z
CFh2T42njchVM+92wjSAGHoqhqGt7P5rpK1YVRGnmYter0fTHpV7hKYpA9ZGtw1FL4vybSor+vX4
DWkBB3yPobPZirzy2nxiDlzo/drqG2XIKCoRtM2hbzcog32cE7pdJv4kjPJ+chDMBfkj0Fb1pa2O
P7+SlnrL+YtmtWqOWUul7XuySfbkZ/NPZ+9xQs7BXp8QaDERSfXp1uwNxGgfufjx7DNVMonLWWE2
kQpzTJK1rbwjJP5yvqFa5Q6zswXKjm79WaQSGYCVzcKEFohjrlyDs8LRY77METEegp7w9u38dNBh
orLg7wFupuskyZH7aqr+Lr6MA6E7CrVnqTJBYXXspiTsfeC2EPbL100mglBujK+r9+5Z9gokhH8q
jm6/sCmxaKNrcj0nBloq+SkD2IAnGtchDLtDfrdHMcl2VO7Nxeme+LsIVwbzRbyQem9pfI35+vjW
0bq4TNA0zObsyhGDCS8bH4JCIMUuirkav76ILDvoEeP0zwMVQo5Su3a7vutw5q9iNeWiqpFBSbu3
v8kwx7CFMM6bwVfmoFLfAzjf0BA9BDBHfge2IZil6QAvFMT1Cw5A5CSRaQgE61BWZ8aB+eCFqFoD
JpuR1bUbQyxeTuN1DblMlvkSziSyjqZmldlnfhg6KXGXrL9bRv7ARBjW4vzok7kE+656n2ozRa1q
aygRBpBqMpqlkxH68TJgQVRci3bnm3juFFUt3zOINpgD+mfBdO+Delp1fsj9wOPonhlhsKNt1wl4
efUfp6oJ3rG0lMpU3vKS+rrD39H5h6B5pIWliAGngctkjVdlD8umSmfqSn3yEa/24mzmO90+Opbs
aIC2vZo/p8ITBBBECd4pxXMPo8lE2+aylYEaDZgQyMgnD5iJvEcH0xWep1pPzfn8yJ0KBEGK3HpB
6hM/MDta/KhxaVJNIwYvBQ+eAPn39NiGuAQCz+F6y3xahurFJFuReYrK4FE35h/HM4ZostpCWFeY
X/8LIaVQxFwIznRGPJHEoeIrkou0bbq+p+jIbb/Cc2vOoxyjiHM91Jo9xqiQPbrZ6JWG076PIJ6/
4U8tgJbDOBKpaHj5/eCMyQ7lc6K2Eob0q5d3yXG9wYM8s44K/zRiCdNLEhHmtf+CFRTy+CKmpfKr
AljYaA8YQOYlNNGv7P7ddYG4SGDh0p3TPognGxG9rStQl3pSKTHdCWU5xUxl40IlQ1M+svc/bufh
bEgEkalX2wyKbVHwp5e8SC0RFUtC6hVjEqFGzlovxxcNK9UNXnqQg4E+BWKgZmIayg/2p9fZG6eM
v0rEQDF8iOY73LgW4HlpImAVJ5ivPA6OUtLHGnTe96bvCg/V3vdZPhlioXm/FSUyBtf/lzGLhIeU
y7oWQFzoSoqiDEbnEWE5/CjZ84L/8mRWp9fEWgNYE3l33WiRWIy1ZT2q2fNk73dNPa9v2tiB7eJd
0I8ELeEsRGqwsUUEHWB+fke9nK2nMGZkZi+mI75RjoC4gbw/H1oTdOiVuaQnHnusdtrNmuCnok/G
FAbgevqLvsGFft2OlZ/ug9ZAggvP7JSewH2wUC5mw7f5FPCdz+VYungqZveM+sOJYKmB7X/B1tDr
zO2MWHB5j8qtBwWRfLumFWaNLuHmfEzKxbulZdIJwfJ87+RcflJH/1alDJCKGJZpUYeRBTQyw68a
5XebIj+YQx1q2n3FJFTiuTQzEnLjP2Wq+SSIizq8ZNQGs6KHtN8is+MN3Zy93CrlSPEC6fWZJ5my
z6NyMOo0dDlJm4UShGED9hB64oCtQ5sKcEESHmzbftPyxbQBNTy7ByiziFX/iwk9AK9muCSiMi8N
taokMqSQ8NauOppb94g2dx+VNoZ2oCSwdZknS0nRrK7rJxjBIPNUjNf8zsd64NBitzeTzlJOfFtO
JSHfu2g9JtA7nvChIZL4PEkFHeJLy0//ipCcc3v8CYmn+S+MIXTQ7//M/VzY7ybyLAaIxkYLVeDh
BMms6YCizxZS9bqc4JDm2TEnhJ8WC2dmZXSRBhO/8tKowZtsj5ZXMQ62+XWqwJooycjqdsqJb0Rv
C/wCeq610Kr1KMSToiiOaqdkJq1xPPxwPagOPrLicA70F4Fumk4vgNrNXnPBm1xp+eaxi6ZhkSNM
tbDCpEDbqwUlIr9zS4dlxz2fZVIFTU/u7ZZn43m003N82rDL6KTb8s/4/k9F/+j73aFeAUl/5pVC
ESHq5q53zD2tqb53DmO3QFfUkK5PJxd85ldIcGzlgHsKkJICQcpE1Xi7AmUUHudfRlEfPAXk5+kT
UIBI0pzOQejwbP3NKR1vR/1y8IkDDQvxy38jNnIGNHH2pLyLusI9Z629Hxt4OQk4/d9TRXWFlcOa
nkBeRmXky/YON+93+GP71TMDNX9woTXbBfsZ99+hhKHJCDdiTD4EU+LbyKkNAlNQGpa2YfBIxWBh
0oxr8u/WvTCq8yC2z5nRWcwdtGj/VzpdAdyI0HWv1F8M4attn41/AArgCeucDqGzbm+xFxKmpOil
4y4RZ+MZ/MMlBlsPuQOxegpz9CJnAmeYRpzCDeb3GaOW0PvEl0B4vpPgsSxlBNnoAcpzVwhzNkA+
lfwQ7w/tQp/mCTD4dU+vtJacfGjIA6X8bYq+ZaQwvRNRM3xO1eDhCB5VfeIjdy+QvdzE40qpCx41
91GuV0PPXIcYaq6VKzS+P/bQeWDjA2Cjd70Z4gLws69KNgsm4xBypsTZKlR5hGfd8NjtG9fmga/Q
td3m2R9Jlt+nd8kFYHOJ3gYQ4yDIc2wQgRBkjg9UY3tGefUWQ/4G+2HoKEvuPB22peq1iTr/eBz6
722XyZWktTzEasOkc8YkWuiuby3l+qpVpNHf3ASUE3KZtyzQnNZsy0UKMDh9aqa6HqJztGDtFjZ/
6YPj2qTFI67mzxgRTjB1qoSLNrKd630e/dcmKWyC8Rep0+a+sz3xsW3DKMnkNoR3a1lxWPjtOCaf
N57K67hHw+/5Z9lb78LNoqwQt+UnbkEfHxLxkTrXtI6iltsZPSaqaBjp1gJbndf/eQxpQx/rpnOg
XyDmOeH35EReA357aD1vhLKu6j5IPSLKHvp1+hQkf//s9Qi/5FJmAJRu/PoEhpBTjubmN7k+AN1Z
KKV4Puwt/UWwh49kNoIMh1RzBAj7UofZ0vcf46pxMELHvJNUXTYmwagca63GTSRz6K+ndB1mGxKv
qmYtQLyTO7Cdjbw1uv83ruLM7+hyQPh2m9DlpCP1jBqhFd8k8IJxZnh6hqkO9Ca48TpewgIKn+5c
nNQsfkHXbp7y1tyonEWojLtRd39O0rf/c84HlB48FEybiLQUaGBzAlu4pec8jBwJ8D8bfCY6YJhJ
2R50x6tfDh4IN/R5YZG2UzW2xIwXbmCu1X85ThRr50c6gr1hsMoCv+j4PpWtWAszYV9FrAY0Ml+2
TioQy7VZZVdrKn24TGcZjEs3nl7iCS08AiISjL+5xfP65W30CGe7lkwE0k6lSju3S913Ah/5VHoc
scfaJa0v9lR4O5MKg8lxrg+J+PchZWbvd1cMdQo1Aw1cq8IFQrNcQEKPUBSdKd1ceuryl8cIWnAm
Zli+tfcT1NviBtfpdJ7bkFsDALyIt8u2QfDCSqVDfb860Qhd1R0bo+ngRmrM1xI2tfh5yS29oOxN
zaHVmvBFKfdchNzHGebT0fjUPc06FThDo4PaXRPJiXxOdVb+L947sE8HEALvf57UdhEOpSXe3rUa
57jdzqq/AgSvSLRIafx9W4RVhj2G91EZLdaVh1mkbmVk0Ah1RTOg5We56lpRo4Q1xZZLwbHAhWWp
yNl15IBBldsXwz8CTONK3hNR5B1OimQfphB6ZR7Tm7f5nX+a2/xaslsgmGmfbKR3HsEcO0Cyrbfo
LJg3nEKqLc86HaNCpw2P4cufNlFPQc/ILoYNR6orw7rgrJqlOgnCE4WVCh9qvbOGPPsltFHmUmY2
Ip823GRuYBxOLEum6ohTg76mWsGiSK2l1mNhurJBU2TGdwDuTrFcZxZCT0sjXpT1zVg7Nz5ocYtH
NO3aBU4KReH9DxU+3EYQrVfYAssu3w1VGZiLtTeAGw+CMU6jnQVYV0KtRMz3y1q16OOFfIp38UU/
GxPuLPpDXY5mJuqQ3n8+uSYbFcR4j5neJYIOs8bfnpp4QeQ0HO4gt3ToN0m9QoxXCq6+CV4IdPQy
bpbn89M/d2lxxk0XN+dFj9fujXxjQzH1s/TNxX54xqOWRbFApf+q8rbvIE9Em0ow8r7IF7HuHIYS
2/w4p/YB9iSxq8aazPchHPGgWziejWZ362ISstxXdot1puSFZNAHELLrKKyqvRy18uCmjbgpSQ3Y
ASt8hbWdNMgJDe/5cVsxn7basa4M1cdysB6Ytn2rs83GcweK+lZm4T2J2Ia7QjthRQGlFDOK/adh
IFxpwertDrp7J0S0yqHqL2XFBAQgRiu9iGnRqfTEiu9k+gR9k1oWs+wU0jK3d4VU4DHjpICoX5w7
2XqEDs5Rfmirqa2fMQDgSNOVUVVUk6uKD7fSEiPAAYYaIdJYfavJ2SRx6LZhlSLIrb9Ri5o4tZGG
dkAEn3eF9yQsIbql6oVKoyQywKRfDjdzadE2IeDepQ1i6ehXmJxZpaGlQzNuGbaBzHHgRkfLB8zW
Sco+q45wgNRMlQc/woelc4FClOLuFEx5dCm69AXH0edby38OWNTxinod0uwJb7jMIhPob7B6hrZl
Clse5n/wlLPaeBtuZm08v5ESRAhKaJ+XBAA02ePPMRM4TFqjWSIjhspajnMTDx10CUyXYuR64qfv
KO+3C2EUjMn8vftMLRegB4qlc0WrRvw0LiQ+xfQqN8pdtXfItuKGw8ErmFfk5jTGFqjndep9mx2g
7rzl5qW1x6u2mSYd3cvt7D5GuEZdXVfYOK9AIu8xmMM9vmzJxtNjtgoAux4LXGfWSD820gkH/HhF
PoiDhOuIv6OI/fn3TMaYZCDEhKZndUJHVJF2AY8FwUyaea6qp/sKiFzsC4WdMqefkT6BsA3svw7/
06JxHfrpOiusvLd7fGWV1fM8giZLTwMCxhlPlV5/C+PhtzN5HZ5qKf/flOqwQxaLl5TnjjKzHuX4
2hOZjBX9k6ZDDcoQ6ig9v3f7jdooIt5Aa8CclDdqs1QF/wzE7BtqAvKUvunNXei0EEkRo7WNGz9r
QEnR/UUZI8bZQr+dyCbyuEB60mN5iAism38JHYKmNG9G3B2PmLKZQIJHmdLsa+G9e4iADSLEG2NH
zb1QcU9QGdGW74g29ozmhK41ZkBqxPRdRYTUA7UA88OxZ1jnaBxl3gu3NgISiNlvTN9ZKBMZVfkI
9QREfec1JKlnxUixBhpdBVA6/kK5mqXkyjBIydRqYjJUqHczqvcmh/HWEWLIo5N0m5tRP/cnVqA5
a3zfzWYo2/9SGsFMNKbLPTOv4vGwgQxWGtpPdFSf33wl+L4MxCLE3xj04x3Tk5PD1amjpP/qwy+s
9t1tf/q+Gf3hX59h8eTXmQPxMyY0z+EYuVRtgKW2Jum+XfU4ZeZQrt2tCm0nDfbbciN8VBD5XtVw
Fqw9D7EX7rYK/jNIugzEC/LRr7ffIx2RfLfD+xywvB2HaXxU8Jboa62ea+P8ZqzYEVlWp8saypfE
IniNoWRXqmY5jbX6b4/GexGCD93CWjPWHEzn171JtxSXyz16WXoJKjs+mBt2GT8jx8njY+ELnEy5
uMNyrsBE6JVWXJI0Y5TWXzG3ZwtNsGc5LEkN/NjH2fJRxqrMDAdhtm9w4hTpPju2CBf6OiSoelK8
5QQIH1k8WgSOaWmRt5wdoWk50VfMcapggwxuR8XLAGIo9+nbhS0QyeLvhUt2JaEY+mZxYE0afXP7
1D7MOytrxLB4FsbFUSbPGzicunLJjbJu+8NL5t4VAuONEikE5vPmPuHYzHRDY1G2m33neUSugUXx
wARQxKRE1tR6AOlB+8GDMOuA8srlpeIxG6UuovkWCO5/GzQX9Ze0FTkOsp0DgjZ8DAYoS+MkILW6
xhlgWduP4qOHFYAYSAMunD5zySuy/hcYDPkbC52Dd5spNAEOwtyGVwfBmTWmou4qhSl3p0nvVwZY
wGy9DZd2uyMWamt6Uc5B0pjkjGV8AO1eAD+4wwuQx11Qa4Nthyr95Q2K7uJF11dvdIGDQUZmwSK6
N20Dm9diNKM8euDmrUGKx8OglVQsJO6agPLGKPCbOVOeyCeiKFUy+1DvatVDTnhOu5txJ+eLs9uD
IN4kuEo2QlbCzlca6rieIPSD2Gy6hl2w/103D69/AHf6iGaIkW36Qldd5ODb2xdiG22LPBwXV5NJ
Mti6C/6S89QXmEd4WK7RR5ZXgH2JFdRRHIarRatN4PTuIhgIISNQfjnoIwi9VUHxMAdKcekl1e9s
a0YU2WHt/G29oOtD+4yW45L1rTcTZXaUBZTc1S6uBiuga7CBT6itcAiEhykkpUHg/qlo0mzLPg7N
e5oIPN/xAgNL/bgspUJqru1F+/ZL2gFzLRE6nOMRsdBBGAp93tP+m8ID8AOp1AE/G9sshjB0p1/U
0VcXY8RhSf1DzDz2MsNgkgopa2802/dahl2+B9hexNpKgt4A07dUfebG1142yFDKlhZE+TJRGJ8j
b0tmgn+oaXCsGCI1chcCg6MNaKqRfq4cBiofmv0wKYq+iyUYd+IFgBBaKHC2/EBrq5YWQwO3AZHN
rNnlE7QYbLTb5gVisEQ+mnBtpeV6pqGUrpYew7Hpcg4fUEfZkKhJnGcoGu3wfEssgk/KZ/3TCFl3
4docv7dzo5lX19XAHdle3b3CKev0jinWyQhWgH3OQFyTfGiiXPMVg07dW5qX9d6FSV4kdVRWKW1p
dpMLsS1F17xUFBWEt9xKXLl3dB/IvyaDKaQ1J6b5Lvc5QbHPK7kIK/wuN2wDE4E7WV2uC1YSHYq4
HeZN0hajK8fw8UEMQRKgvBsKanwI2+oK/6+5zQKCijGkmmF4WmbkYneXUyuGDF//r2RzPisGU4wT
XaDuXmkMnMyRIKtP6EayyeEW3Qml4KocXa0BdwAE6k/rk9Ntf8SzkUxGeUb27QHDIMezYcyqryLQ
UCWofomP+paA9StquX2VtnphNdxBLlvQs+Njfxg8wqC9TucvRLXeXpSCuz87VALOtlHUH7fmoKCA
TSM4XCFC6b2nuZXUKezJcDreGMtlIWLo9utK8Er2o7TtqG3JA4o96HvOBCy/rzvFBi8XIfSbPZ2L
EszsB4CSiYOYCNbdPL6GZV3jz/7vc5ehoVQJZuUf1qEVzMOTaR2+9rZX/gQRUDFYb2xzpqIetBOo
V/lf7epsOq61MB/Hgh7UYJo5Yf5T1S1YKiXoBk7q5Ly5FC8RcfLF4YJM0hLa0ER2lQZZ6OMpbQdy
8V1cjJGom+JgSkHmLs7kgybApLP+IMX8uU8v9ZWjIHurmp+WKJLtslKF46GyAxNlu0JRA0wJR3p4
+3GMPLjGEqzeg3p8cWNonCjNTGhb9ApRuKb0X667qmY2IrGPZ8ZXjt7ATV8tDn/LlP2VoYYx5jy9
pRWxLRENFc0B5OUZ/WFMXJATMmSUrOEWRrT6bxK2nUe81EUTNNm8Ul/sB4B6MVFsHdI14QAsjS4i
sw68bsFsuJ3qmk77M0hviCWTO3CK4SVTYQulvf/5q6mRXi0c5T8WgQPp9r0wnUmy35cXqzMo3ZyR
orMttySKoD7qQdCJCPqMuFJzLZlRN2aA3HAa9vaQ0HP/lloXnSSypJRmeGK8goGQRQ3Adhwo2Pph
VTwfrs5n2iZvPaVha9xRHkROnmxpmW4S7qjRHYFYfj2mZVHX9Ou7H0Oi9p+xdpl5J8eIyJnLbrsI
PitE3vPA+gCnQhKf27921hycgd2i4FLwybYv7TgsXt9n/63JbTn6vq0IEZXVRn5agiq9BsgzvVwD
Sjhh474sqNU3vI0/icK3wchi+vPoQzSj2rs2tU/kZFbZEwiYxJz/N/hFwA6zHO3sX3REY8nw0TrV
yMaP2h22AqefGGlwfKAg9ZhC9nN6w6WEtkmcrKVFfqumfRu3FVWutOlakD15VqsPBBR/5DQKaZTm
6WoNcuOC8HhssOsLb95qLDGbbLd+iOetGeQ7ijoE4QWbWKwOFNg4DMAz+5OI33tZtiRpesMfoRKA
ch9CZHzTqXm5kaFXPrUyNNOxqAtuAd5JCmVSjYuwHBiEdRY4csoZAslkRlpGZ+kJYxb2W9klh4TK
HKS7CKRQJK6LVtv8cHlyAl9abupmXk2yvnJkJ3uIcRa5dhRdu1nwbOTs2Fh+BdlLjbKZvTlrPHuo
uYNqO3WMFFXSMpFU0nbzEZ1+GJvNtKHrJRTKA+kQtguZ9TvT2SAdWbLcmQWx70FDHbwt59MydVQ8
v16qzKKFuNCsVjGSqLC0HE6qbFLh7k+8G1eUmfnM/DkwDPqOH9b7z4SWB8/uhI3+U4tbP6pEXKz9
GlX4Gwmx29QZDke6hE3SNh7SYGuQdT/KAP+fCE7PRWCwZoRV5Hl0rJIIEhO2g9nB5jaQ/CB5z08H
qfpdLAMYZ6iE2tP7fDSBryppI+o1xMbEo5RvGEsSlnSfzN+lBJ+JlNxDHTmlt3bGD1Oyh/LdZHn7
y7R8+soJWx128tun5gD/ZlsG3VmHRSgXmCiuRi2U46Cz18T1eNcI68XH6r+bx9EX0BI0gcV21yYr
LW+zh9BlsnVHl5bIkYVd0pbnskxU4Cq9b1bSHRmibTh58VOXIyhUdyD+NJ2ETX/y6uBVMxJTXBbX
YE/wy2J9F/Qi8r6MUgcxFA1BARHfJNkAEKlZ7CgXZYRNWYrUsVNtd09KskR9dcuqbnp0yk2CiwW5
uDq5ObDArLM6+U0YDtXUoqiScIL7z/2DXyK4pO7akexvbfim7vh6csvdvfKhGbU32+4lKc5yY09s
Oj8s4qRewOkPmsHG44A26CQ2nHY7J+BAT/AA31tCHYQQZWljsR6hEtRaThiIDa3PgsPGf8QzTN4Z
Kfz1i0PXvwbrz0u2VNWlP88N7SuIDzKjCKt+f7iGsWA//I8Its9mEYJjkQ98sTHP0KK5I24px4pA
UePMDvonit1ZKAiTFaQT4TCYk/Lo0aUNb7gb6ioqQbXQFgHZxB0rCbi6W2hD8EbZmtiN2MTwDb+G
Pttq1UDLsqilZltnzUbJKNM0vLlEoT5qZkDUn2xqJY9ScZ+GBBW71rSIkOEvIhlYQ3xHRryTRGjM
3r+03rCsixDBLh7Q5mIaoCKvCsh7MvQmOsuzXbdsHsCsdSNJHnPk0nYoVvLuaj4J/tqYuC8T9NN+
shnjh4DRgv5ZrNTbP1uuaH6xf43ZAEn1l+6ET+RNqs9B++P6qmNdfjq9SPSqOsBiHfeNUBEgRoL7
JkXDX6/ha7p1iMV9C2rGtShHhfipephPaZWkxkC/VkFIUSk/ohbNcNfyJlK4mRrBd44p7Ta0Bav+
ZmgR1d8lqqWcg3coIxaHOVMQvffvIqzhaxT312wTlg4YqyrOB/3X4dTCGVuF3S7reP7+wzewreWj
IqwjXpm5JaoronUWBjWnwgHZYIoyvgN7ZiqpG72ozt17bqzeuOwH6DHFpf81kjkqY6vCrOFjW9PO
7ITtiTRCjUhC03hCcE+aBuQzsyFnXH6CVA1qUTkfwC+Zmxa6QdPng7tJLfduppD++qhwNkeepmYe
Xt/Dws5XEhN7G5NrzaMQgErwTzak9aVkYmXr6u9TDt+sK8UyawZ4sLxO6jPY54CAfJLvjtw2aeD/
HCojuqsF2S15M2ghMHOL84jIzGJQ1cbm6XZiqTY+qvHSBubVR96KoKIFRIXoJS1tcA/1t3QoamiZ
HLdtAExGn0lH/VBgq4GdM3rhRMPyNixaeNvrY2JUM/gvnj7Ss6CVHK73C9J8dDYQYPeN8B7r8R4g
TXlA2lFIQmXhDZcWPeqgkxN1PHj6mf1QQ33RcDe8x72zIYtx/Z98paUVKwnaKlRkKC3U1GQL3V+q
zEV0RBED3SbsHofJBWLooofhsXVd8w6SZ0SbcCiItbWCjAISYZRqSw1i9+HTzjA83cuInrTzZ1k8
nYY9Zu+gGfFTJWXJtsgdlcHVX3arhFUqvYc3tTzfKiidErpfE/DwtQLqzoNtLsztnyT2r8kVVOEX
qty5RG6zg7I2VBRcLLFMvk7bm10zs2eD46EjzKKGKZ2KrHa+4XgDqSdRbqU4hTDOqyn6iQq9SsgU
o65QC4RwK3HgjZCn+N6PqGuznArl9t60OO+Op/VS5wtSo/yZbM1q9XJ/P+WGIHjco0c8nnxGYqat
AhWSKVLpTbBuYXt8wWsq/kMi0D9bBjEfBu2vXQgPHCbYcT1lPiwwbEgUlG3mUUazixFpLOJPPsHJ
JNkESy8puedFsoeTkPDSFyJniMjWtpGlrYVLhMnkBbXenC37aL2C46uOGnqbzPd9cMbw76Hp71o6
huKESFvNEiGrAtRHF1t5ID45FfAReD2EX+hp13h76d3vH0axLy9r9Yimx81Zt6ICu+4EK9DQPsxL
ORB3kLjCA3/XSyntR9SqCyZBe9AUzVB7DIMhgt8Bq5BPWMBbjiXVYFwMtSMkiv3ArV5sPiCZnya3
sdwq8SK+l2pHKY8JfgtelltXy8qt35n24H804IUb+QX3PJsaVN+tDHHDuARLv0wsMVCX82g4lkfa
acRIT7NrPhr1B+6n7guMfmLS1ZuYTuEa7ClTQop751SrOws6968pKshK4cbDtX114d5RYJPXsMWd
wD4VrYC8beLypPknumxepXorl7a/9CnMIJNELNL/GTLaEdPlY8bgzPcH9NOfJ7UUc3W91upQUjV3
aPu1ls+cuF7SKCTjCL29rx4vlfRTMreyCZqYvwt1QL3VBqnowILZMTIBRIVtUh0eLf0ykzqfH/qQ
71qbzg6P+VegYcU6W8lbPuRMULx2EBeBzuiUo6qalPDpBOMMQq9Bq11aWmmLWe4l17skd4LqELyQ
DWOTAQ8t0NkNgVXDeg8FRMafvucySvDPvLEFl02Tt4H+fsWRsdT/KMZaNjseZlMB7PGLan8fwgKt
6+yNlSKjeetaJHv8EbrLpaWRs8Oz13jAiduZhgB0UX13WKlJvICpyKZ9CQY6A9ex3v9dLI8BgxLO
+fyMI9rMU8BrKDx7XxPCGc475PjxRRh3QPWs+gKUSqDHySz3zbqLRdU6r5aYH+zbMsj/RLti7foP
z1J5PRcJyYefwc4BYPxOq9WJO6kXqLtuIs7NaGUt600D1/gJiIm6pDoHUBpqNR4iwpcrYZ4itYlf
zan7c14TFmp+nwgiSWtpwYgPhsq61QtK4IPoi1em5RlVLS1Bzd+hVab/xurnERyBKnnnn/LGdfFC
y6lDoeiMTa2hba36ZzHfNo6WDUJhtzOfGjMJr52hbLPug46GlBE2IImjykuIguQJgK/22DucxOSs
IkNETXGiuvvSFsppwGdnVIQ2RwGuj7q6c7nhA+VQ/xzDH4gzjgjtjT9PSzhCLStqAq+gGVn7fv87
Eg5rrIelpI6CFLbUY7E2leSCtUqojif8SVCBPxIdbfdTZ+prxjGBTEK0oPNbIwSaR9QtysJwq+cI
4h81C35bttcs4KGM+FGcCJEjDelRfermAILmUhCBg/HLF6CPfYdwU/rx6fXr0Ii0qb5bmVabFxPo
Qz/p2dcKD7I85Al8ntUTUFPsuUb10kqjTjkzr53KE1cbl/z4GABOaaDyXLNenR0NLrNcO1CmsF8/
vegf3QSHnFup5VdSUF+dzvGs4pxajAgv04sGdV6VtM2GKpx1Lr/60Uq4pN3UdrCLnjlS5D4hjEFC
mTkRhy8i6qml6G2bq36W6KX3wthI3XSBj2pRXYtdeJDRkrRD8XobX7tbiSNej+pnpBwDqlzSh7tF
tNcUx/aPebsfFEos3KyMhxiYAFK5INo/0GZyPqLsiBOY6fv+AAL+2qY6OzFDxb6qc6BjdRenHmmo
Gn7VhO3YMnAat8Kb7ucl/6NGaLs4LgTJ5Io0lRBEKHwvgm/yIGD9xL/64YfHUQGHSNAq7da8GWwO
/CkuQd7Oqp1d19ZJpdKEtEjaCqG2GiECXxvYHyRay2Hx2a0nYZwA8T4eOB5zLJYiG0I8loSFXKcV
llVyvjOGfPfScsyCcNDnVGHAKmi0OYVbEEnAZokJnJH42hoKQ6rmv+2RX8VyTBaqz2J36RLKcl6Q
AbVz28oobC8Cmef98NI9HAkZvF1QLl3hKI0RHaXNHCJtvqNf0B6a7XvxrZFgWoNu0QJcJppmyLUL
/i1imW4AxocNuZxsmiloyuWJzlvJRQQiO2ORrVep0+1rLuYpfDLS9Ami8vcBdT4JS1a3L/wnOy0K
OEoYmz7d9hlI0FJI2PGk2UKiR9k4Hf/yDyeTtk0FG7OdnfvuAlMXYZMpiEhKKUudPgQ5bMhIK6ax
c3S0W7FAh5zvHnL7pej0vnRaHO6hMebvZkCXTLaVtJRRiy5KVJFT8egSKpHHWkM2T7etiFrITMon
EWn/DbsQeUyNYiGsAaQOrWBpFNWQ7mqPmHdblzZ+hmqAJIy6s6mQaIGKX3t0GPiWYTaO9ITiAA3I
UmqZc7xqLUqIvVc4Ik5fbWz/oAOn+9EHokcf/2USqVY5e/PeGKsZFbpih3eS7JZkS0qgJhGsKy07
FVX+qCxKSgeqPvwm4D6t3hnVm5cjVJ99G7tWMCBYcMRpM3T6ke1Kh+qDa9288BUFZCzXruBVyU7k
0khMzEgvKpunQR+i5lI2ywZWi0oeeiN7MmTr4JklVhj7O8EsKaIV6UM3IStgAR2z8LAdcmkRMbh1
cZICtO8YdfLT86tvwHWMram1AihiTdU8ImzhBY0TO7+2t3tcWoC8imhI41+IHE3QZhN1O2xttro5
64Jv/Lq7RZzswPl8HKtldCZm/4Nm7Sr0gBIlgew0txTyEuQ0Jfk99eSpDE3qUMGcAaTn+8R+mwHE
tATF6d+ooVVIh7F6Ge5gSv5YdN002NcFgQdePkhxBgLuLCn66Yqc+6m6QG5+Fp5z3RaQCBTLeUDR
oFsmxLx2bIlCubShg1LCrrELSMjdLeTj9zbISW3wgpFem92teg+YsaAyZEVT9uieF+bbDABFG5Nv
ToCUuXM25q6SzvxxANKgN9ELdJI+BDF0hzN7U5VCNJu/HFzawmgcNvOHprpiZcyBP2pQDQ7zOf1Q
gIYF9S/UWot3v6YxLO1y+V6jJTt+AAVxXfHeymNt/vdoCxqxZnk5pOgigoQsvDLNz87jGfLAP/0M
/thSqnVqBdaVNbQVglWWMHauqtIRaV7qeWprhHWTu1kRM8SA0MJme3jv2+0FfaxN4a0diJfMNW5o
j4pvPYJaPqeGSlrL2k0grPhwXsWvtLqErFZdLJ8dQPJS0MHeG3ue2cdzn6XgcLHrKzk3jIFEmup1
6tYJ6VGo94gykKswuytZVfI0EXSvXFKGsyoEFdLR/JtdXMItnyWu5w5xuXuP+08Dr7jMBbQvt18O
gt1I7WM3ryp0joCbgHhK2k5UMsBgrwVvL5kASlCA7AGQ1lfh32Ng3OXhFVqDerplY7BVVENUi8Tz
N6Pk5lpoPFyvl1o+JC3Uztoyvmt9GTa5x2hfd37tjz/HbYbMR0wGzLV+WVLLNQq41qzqwaXkGopl
dvenIzdq1oHQl1B4WW935OQk7MBg07SUirDMYP2eqzKpTnlElIGftkQrEVrX98euePMag2w735o0
hhzBjfNKGVTyHwWDLbjyYx0ujVDceIAAKIXQhTYoSRB+FrD/6JxIwbUUxJT52SODRNx1fprTvhKM
ZwPQcqnslLN7gk7KlRH8pknrSYAUOQg/+2M2GcO3IfkYQWr/u3sUQydK+bru9j/trMW/sZLW490d
OIxAijvNHrfgjWuvGTuK4x6C+OhqUpJXKBm+9QERf7FIZC6r4LWNdC29eTMyIvcpgq84aI6nC4TX
U8oan2lbsRkVihV13YQxyqEUdnMe9qucRxE5JTsksIG2LLgIgSzrEQmCHkaNHwvQaebFdr+eSQR4
hKUzzlZwblQy7uTA+YSfaHpxgd4iQ7Res1rIBKACBE0VhNvnBb9IUij76VqEe6mH1baK6a/w0NPb
GPewYKXI5U34u89YyqfQ43ZrreM+rMzfUS3y/ZOW6s9o9HvGjGVuHaksT7HFN+g/5VgT1/U/ZY6U
yvvA8+oE2kbIJmPT2YAb3AcDNZaR2jzhEFWeERZHJ7tIG0rc/KvSZxVqQu0ipheeGb4d6drzEiPo
Fp/yr11XhVkNUYnUMyLn60g08y0vGw+RlAllbVP/LC8sVPU175riSS5m316/1ykX0/H7Nc/eSLge
KlRDiPVicrhg6h7UBa/qyHNeME2+Lw6TxOwuVlEoMI74CqatBRvBVUzb3DS0xjGJPU4lg8u0d64v
T/Tf6bfBTkAgUJ3K4ws2oF/t1IxNQegj8UMW+Wgp+XL36uHXXbuTlelCNEYYpvheLz0nrzcdAhek
WLhiCrmGjhKmw1okH1I8Yp0ylyVP7Uc56nbgrmCl7puvab2ZA4IdTBNwpfWMaknljsUznknMOXL3
5nwV4u0nFbQvZd1hFm6GXp0rtfKNmdB1DtOERk05A8q+cNIsS2wzSydY61NyzCCxpu9cxy9okeE/
v8N2N7bvMijzy8bpK9Ju2daxUYJ3Hk1Hm6Zt4gFtgRc4E7AzcERB2vwy4LSbNR/p+yMwMpd7rSpP
OdojgSSYuzwQQhXRkwKf1EJiZQJRDU46OwU0qThuhBkAxczQo4NEdFdNmzdARhPAT6J1VO0VvMvq
3hUileg+en5VbFNMTkPfMqhKMkqyXqI9NGHYQSpPO6MxIThm5FPC1TWAm3A7AtFa1M5LCuzPh+iK
CWRO4vUGWQY+PjrvVKGubAnF50TurYamhHroKo4E/eo/AGPmp4SXJYZA7/p9lQMXjin3KLmGShCe
OWcGB4Pw+orsxfEr8AGJlcWqs5LcyyM/xZuv+Cj8kHTp3g4qWhbTDfh+RYki/clq7aycZ9+faSds
4JbeJwRS/N4gv7tZa5DYtvJMxxJ8ihKGpBOmI7zHjpIwMOHJ4kY5twXTfycvN11BkD6aoJTClJjk
pmGwvAbn9DP9t5LJqgz5pXxFXqwLd0E5MVC1ZRhgHUd0TGVGmEivZ3ldfS2iUG/abodSUQ+HCx9A
QcGQ4w7RClStmZRNULbyb48XjxRVUmeyHp2t1hhNTwFuZthuJgXLc4qSdxfuKbx/7J7aUfB7/97W
6WW7HKypFL1OcWCBfsjquE/xqIVbev4kNTraSLSnWNu5C4K6+WrnxqEc8obI1QIrUjv3pu/yHokU
TEKe+Px4Gnaiz7U7yrIJhxKAd+7nboNWu2z0uOjPcV9ZHGGH5dei0X6eDzRR1npfN2ok6d59ckoY
JPJx4pqCdmARogpUqNt0hP/SOfrAgs8LF5WdpV35CwmxOHP3s5lK0IgjOmcP0eI/BB7eYRy1sWZ3
dmMkaRogRS9EBgl5bDdQGzoBrR0nVDUQ9cr9n/YhbdNB5HMocHdoUQm+8jV+kr0mHzN2ATZwRxo4
xuFw0Xf0VgJ/z938bT+4uQRxwnRjKmBlJLI6FlJjuxpsfV2Dn7DyoixcCt88uBaPVlLAg/Qon80C
Z6jHQB1xHbFRICff8nYiWlc/jt8qR7JudY2kaCAAAYrcvCthRT8L2y2Y6/A8B0ITnl4RpfvUjSxj
LoP9DreXIcjSq6TEAhr3rcmApIWLgYvWomxirN29PF7CHUgH1dWnouR48JjqCx7QjpcnDqJMerdg
7VTkD6psGXCv0itd2GhSd2hWvE8/oBNeGFVpFSSk+PstwOykQNPssT5ExYriMhK3UPnl6HNIvhbh
2g6CBj7Ulv0/24SbkISH11A4p2RbcUFxX7rryqbnWzunLRIxOcyk5wzIHJcW+CMlYCHB9W5JqOpB
vhO51BYvMZb0aol2lU7IXbk4mwafE27plsT5pImWWLHXWpEA6Ieoyl9zZnMQHJBNQyAMk3uMtTJs
uwUGt5WWaSzxY5i8Ip1WSum/jJew5WklGIbkEZ7YBLUbJscLzw7FEszd4FC06K8POkp+/rSlAlbr
g5zwqYHLGD7dkJEOaCPHelMTfVTJ4LCUnRbBlU7+8vogDAEj0qP7czLsmG9O/DAZWgnoch59kFcy
TrORF5TrHPFpAgsvNBL3ka04n/CXXFLdP94vwY7FrzarSXSB8p4zI7GFSZ0Jw34QwRnFD+yuwvmp
Wrqbyfyn0PnaN/OZDbZRwqvW3vWGO0LDc9O2wKiOi8ofRkKPIC+JdHRdG3cWKVsRRfUFnQiKWnI0
qhZhUjJHfTkGSIavMCb90yWku0R20vskmyQINO7bguMxsT11+OaRZq/J6aVS0NfmVjZocuQFP0LF
GnOGoaxSyn+QFiQSrBNxVX1WlTN2P2DRsqm6IpRdsNSAOeoAfXGRr3/m5MOF8MvE4xPJjQXLAT4C
iaqU723P7A1cxU1zmXOkIiCjpjuOI1Wc2DY8yrsBijjbsQCtlueovl1Vq5KPMFTN283WYuCgl4fe
lzDtOlLJF/QwbWxNQZHJ33gltmjQj7h4vkxIReZkYMIFUwy3VW5+/D6QNufUuCgG/D/BK7VmZ3Kq
7Kfdk0Rj87tvSoXFcu+UYKJ5PZ2zE9H3UKrm3vO099RmblfKenaXiU6Tc0l1uGMRSrcQbRa8eLAl
jVTOpvf3WNA0ZOWxrXgrEoSarZM8C+3eILYFCQ8nu426Ax5ehLG4wspBpg1L2DpCB6e6sT6IfcAO
WASGDQkV/OniEbboyu13DDb1PPrH8ZA2rSueFgHCsga7TUjJwyqmi40VmQftSntlrLIHOZAe819u
ashXFXGyJEhx9dUge1WfZqj5+99XnaEDP+c7itgkEhrV36wWh11G9K0guFlrKiIP6OEgJH4hdaP3
sEzN3WVQUrfkQE5XOQdMqBi7DuMB18+ZAOYA6/nqz8JG/PYCgZ55hvFc/UNOoMWTkrGbgQyw+CEW
6J+lmuCP6kYylscgDLBp3fE6RNmYQbtFXgePOwtvvPTscRnmEVPQVnlhgh0cUxKC3nz6obyFQV8y
VN8rkf1hdA72fqkjUsQ7ZTcStqvsBJfSuYa0UhVjFVaFNTaK7sx92cg/CZoPGIAe5Fn7c0QeXTO2
yQHipiyE7/YnRV+7vm8EE7qUy6C/O9PnK1jycRvd99TwPVRAidUXhWM3yqOQe1bP7ivtos6QZDAU
onxSz6GIt5o1BQK3v0FOaB6nJMmycvALwdnDW3ch8q2TbhwfeeKwnkoqc072Vhl9c8Ib3B7KIN4g
QJCp0DGprBXuJm0ylU8ZMVwqXpD5lrtrdDb3q6gvuFmHGay/6j4ZHeSvlWwRhzomwq+pHTBa8zYU
aKzE2k2UQNwf6CwSW5g9EGR4ucQPJePUILv1htnqGku47npx/teUtpuBQKR1cteP2cOytZvfcEi9
4XxptIYtcPfUdv9DS1k1duklOj3QztSGgysY1yhSRCeCXCwIJr5B3ksN2akp0ospJAogn4R0QwYl
Cov384ZczEBS1z7gdIQdj3isW94FcbF3KLdYLfqPuJ/BoypNxfvaom+MeDGGjtDVjEiPDHOzZMCh
0pSOcvJCOMtIzAqT85ibdoQN5ui72khdc8A6PwbdCUFmcqkFyGmXJffmQut9hZjpk9V0Y5WlGNz+
rw/goDb2uBc8ZfpDecZbbK99FTaG5gPCIaIfTQXji31iFYUc38m/qBKqzmU7pubDedAMtiA6dXiE
PeqlyozJrGI86blmvXtfGzBO/+6BrnbGVj8ExletQ2Lr/lhnLdTwbvU/sqS4vfo//Xc8ufmcNCTd
8HmVz0DP2BA1RJyPI/x8hbcSbVzgl9W59+RD9TRW2DlYV+ieJ/rHX48TZMr2Wu3Ne9yF2cxpBUO7
PZ+Zebwn4Xppuy7/T/olLSnp9AK0G83SOfbMVBV7PXhSInHwS4/u7vkfKCjUqS2hTg4vlCKn8mXO
NbWEpM0bXkRvQ/61Pd/vlyV8F4ENQQ5FrM66R/r4v4e9NYH46i+58l0LXrngNDlj69HplJv4ZIS+
QE9txv7cmO7XfJRgnjwhOg/lRDZxLKondZeHO/WlLgrB2hu+fVFIHmnXdMiewpEbRJZVze8nrMAn
JTc5iQ6Vy7rDPu/Pn9mHqQS7Dpm2X6IBd0lNWQbYTKDPeHHSDyMu32Dk+2XiRNWB1hG9A5Y7I5UV
LEsmeygIP/dT1eRK1LKWm8W6YNo6T7k5mFsraXk9g1Sv5mDzf6AFbImgB8hq4nv7D6t0qIJRv8wK
+n5DleWHlMZcG8R9dKEF2R9XB1X2D3SUwaBDhgzg0Uy+wNboGvJVhI4jVNgzbvTlyWQIWSmBoJHY
DuW3owJTVOxin4dLQp2HcSq3xcAqJku9Gavv5+pQZFJHhBawSYYh5w32b36C1Vdf4gRRJ21JW7TI
6bY5yexgrW50ggYhnt2EX0lYSp0kY7vyTN4FpGY8T9xT7dstsBBZw3x34dELdSGeot3gMjzNoz1l
NJ6CSGCBFYTeQema/5gb04YOgnlZ1JIR2xAasO1Y4IzIDXJ7zdkT9+7wXGYs70HLHWRXz6ZEiUnx
p7qJHmp4OLLIIg2YtvNDCejGqWEFZPHsJkTModc3KlesYARwEGD0Z1FJ7M6cqp12FZ5WQpsBDyVc
JH5bre4IS+/UhrlNZC0akbXLK/FI8u9WKwZ7Fyhb5Ow880u5bjhXv+KNTSoEYpLyEPYRXDTTfEn6
e/V2UaJ/OEcE8CtLTiU03RR03xEtsy1FA6Vevx6WC48QdTyMJnVJ1I/C2fvcX35ePyrJF8ipJz2x
+RuMm5NJ54qmAt/bkYOIU9Hi+O/viUEMsFAtf7hsGB7/naBBKTWcRaAjzJj/YZshBUlJw7aYFJSB
mx0g542mWBNmXY/OwFtDOpsjsxDvK6jL1+bOsilj9T7VfeMENYBxxihpSuLeyGd4XAbPtAkjBacq
6aiVsgdooegypwBuHqGanfFrd7E2Unmui7SwECib6S1a+c9b/dSvb/tYfr3zmHOn99qj8rvocqID
6PFsqqGkjze9FI7KEh1Nrhvr4WYLiKfH46sO2t0ShMzjagfF00xFa0aUtkmdD8XTw6ClCc95yEYL
la+w/gegCKg6CVIrDSz6zh1aeXh9VgMXni/g2ZWCocl3wwKAdF54A38cqRfdtx/4bhRJKD6MPN2C
XIe4AL19B9yrJE5exxDgkMryhoa2IyDoMzgJPBN1BtRkpDFXVH/aF9OFg7WeLQ9XZDFQ8H/o5L2L
j6OzJS/xkBmudvFAj0GaiW5G7AfJXW1sMwkRCUsaPygJVPv1zb4j0KqsfPuDrh3Vht1/vTTZulhK
aE+wsPH8lEiJ7TDOHMPPHeIeCO7JxzVo6v+bOk6IvfdIceP+XLUYhRTjrGFoQO+m0Ni5r8CAMlbl
77ucdN4V8NvePeLHvRFV/2MmBdt4b1+JwKz8dRMQA/4qyag9oqyrh8Z8g24v9HpNx0+rjOS9Gxm0
HfMXjWk0d2C2aPB6AA+qcLYOmpFQv4Tt038Wze+sylMjqrsutXnbNbEd7d5uNRyc/tsBvYF2kefi
czY8YvJxV98WAYyprH8wQL+sa4Km6GbpzHBwu35QavMhBPHZTQrGfvYNL3rAvkym5Px5P64w4ScW
fpqGZ0/fQuDUBGYdnbtAgnMGMrVYtngE1aSRKWexc9ZgWrkVy/DW11piWbUW1W8lVFq5PWJAmMeB
GQxHg72s8zfdTwc4QZD8m4U1S2cwh177gtrbcvfCnJub77Y45V4VVTlrd84LjMpfLmJQnguzdS9c
2/h4SWFTKd72S6DFsmMqffjn+/+H57iLFWeWH+TAnJa9lxAYAZB7As3jmoLgonCVPAXUSbEs60bc
cgjjsg8sUvJh70HsFskV+t8OCEmJy0aJmFZq5yXmcvrgGiBMnsRmAkyyYWnaXNPdLFXxFpAAAvAk
v+fV5hZksRghWJg+ZohqXi/HcStsa4Wmv7dis5Ny+MECe6Ec3K7YFDyMlL7djvD2LIXmRUM5Z7O/
J+XDS8m8ZWZPgZrsrYRyvxw4cwnwv4Ow6KTizUyIMZSk7Klj54b6zfD8b7JmyJSEMxc7m9uhqyx6
SnypngqS/GgslGMAONiJtrWxw7r77M/kRIUit+EikqOVyintRPgkJ/WTPGE6hPC8XA1Re3ypHkZR
Y7VoKGzDJqYPs5RgkucQngqaan81yqOtJqz7xoomGGfsQKo37SXjIzidJQ00aKidYhyA9+YcYdyi
k1TszrS+b4zv4BAYcTMBjg1GyukQcjoV7eoZP5qJ5iY6C7Gy5uQilfdqmba1N0I9/cERNCFf8Uk2
oFwyXlS4qZztat+W+V3PhA0baGhs745EZ62nUmfNzYW40BTTvalqg1vJSLmsHhR2L88A3+3WSyDe
cEHVTVGVOSia09+e1EH788h0yRCN2MgPZoXiQnp3uPHvCZbxzZTSGSyiAyeg6B5vWWrI9Jft2gPo
+D0gt8wASPgEcSzcfH9mMwZVn6YwojoXU0uxx5ywd3TgrNVzFGsgm7+Ql6XYj9oR77G9gF7xCIJ8
gihQLUlZBQSd6Kdl4DLs+iiIBEj5pfgp7vyIPVUNGdQeOL+mTfyXkYL/V3G+qz7JqCzZaURbvwOa
3K3WhIvT73FedsH4zMSC1ZAcpqK2SFjyodWH8a1wUOOoIvER4CIrhiKUGVc/7pwGLnexN1bTV25A
rE4Yt7C29Kg6m7ZZ6ql7SAVtAv1V0QYmJGf/gxAnMAKy17WLWDT5ti2dACaLLPPgilOARkfcvzXA
wIubn5La71kIJIjzJrB2vQNL4cT+2LCuQfDASFcn3MQa8Ci4a8tcebXbHEinknejqfyZxp9uyWGI
5cIdcSaAgENknV40RtUIhAm8gceJIRyNcYsZwr2DYBeI0B7rnKQg6Ut2goqQ2U7yvU6xLgdCe0S2
jFPfE8vB9A3yTvF6vnCs4BCaxpmKUmeaAggHj0agc11lac/t9/EXdkS8cJ92mzBjAlzyKbZYgncp
O1QB5etVd+i3iIGjHY8DQi+s+loEd5oFXx4IXEuVCg6NnBfNT4oShhFC256jhcU/dHc4Hom2blKy
v2KJ/YMZcOt6mWKXYsE0O2LdwBjxyl7r2rRa8wfQTtje+8QGEgtb6Z3eDDDr+IuSv2/YodvBAxQq
XX1nis8af6pXrt05MiS6KTb/svUtDhW6wJcNq6uGNdY+EeWDzD8UuSWIg/zyMLDeqULzhtzsvdNc
ppPjAXcOAT91Iub3JvMLR7UkIphLHMMDr8NU6s4VLd7XBkXYDEDzXmlX06J66A9LG3iFiUaNG0cq
cyfjCBAkss+1o2dC6r28SwDyJaM6UaiC1sXZqQe1XpfdPfIhMf/MO8KG5bxb+X8Gqgieg8QZuDPo
rFZMnGCzTcS2caxVDUiOHiyniD1dg2bzs2blNUELLq4b111BrMbZUxWmXXJd4HalG6mpq4+6cLpJ
QIjVxt5hN5u8cacbd6TVH477Tg4/uYFUUWb2Qr6ctyMRrG98w9e8JY7a8IV0hVeX1ql9A7npp7ox
z3umIipu/hJ2LoWaAbmNzzNha4l9ATlBcB4xKoQ1ekVFClV32BiZZnemZhwO5MQHSO8Ljerl+Txr
msLw/EdlNyEMlnPYgDamnZxYwFgkPkEtjiyuZYHioLLvtKK0PGowR3YgD0Nv3EEsk2zxT5tXs5P8
gkkUzrM32cgJbYOi9du4k4N373Dqk+2Ileb9kzaMaHt1nH1QdcZdI0wp6p3MNVoVCZECrsXIOaCt
jVpu0jngJgpE3e1jgdlp1rOU6aqfucqfhzyrxjiGGY7XxheG32l+N4A9fSYxoLM+1B2VhVgfwFsN
rUKS9PrMETB2nZKdQ0vI6vpsDttk8E9nvCXnV8pX1pX7utCIFE7ZuJdEuVBfnKCKC7bBu5alNGEv
FoVvdbqUEq6eOjFU/bKgw0SBlopyCv/HyMf6CxrAwjC9RwHhtdJDZFuMxKqpn3TJE8vdMDQwga6c
e/+/VE0OqzucAAdinVimyUayY8qIu0Djy4QDDqfEr8x49xoqINna4ePLiXrOwlP1oBxnfhnHu41j
7dKNYqgePzrH3vijDzbsSTd23uhdctA9Y/50L1TZck8trQp2zYfHghf6pRki197kLzgYEYl+mNMG
NJnxCvype2SW6j4VZyz++s2ceV+PYbRy6SVA6fTIxdJxdY3Ft5dQQvA8ttRWKGOqG5denb2yB+Z2
dCcovryPLZRddsLSu0WlNpxV6TzXFysoH8KP4n3FMlJVSihucn2EdWh28dqgyC/F+VR4IWl6I1/D
DJTjIRD6DW9/mwOiT4Hh3ex9dTs7rPAo6GH1yp2VyJgRBBdMUGhtenl+q2KEsHWb1gnGSK0h20ai
A897mP7j7tIahnDWidHIoSFIT05DyHXSw9PVblSiXqfwHAoPMM7+Ef7uiTQZ/wf/1ruAcVGIdiEU
IltQdNQZ9d2HSGxC8hkUxxIbWeorRjRoYf6OqfWoG5jF1hKNdPEU9+Q/+r0mYpOsM8YgSeYgrmuO
bEwy4TmrJ9FPpzzuGnIU2lERgy3fdG4jwEq2b7NbkxAcgMhOlvHRZsdsKHA0pdZij+H7ekTCzVdg
wg76Qh8TeAQ1BwQ4EYAjZF0t9vkPqQw7bH+lK7gjs4LXBYBDYENAkcJISRF4fcqhRyxMDJ183Dmc
5pbUsI+QM9b/prAfCEgkggsg4PM5rd0YI0mdLqzcVYainopDNRhxsI+AYM22ihl+njWowHmBW6nR
iiu2/VWXUWsv8YRDXW+zmUjOmrhl5XYe7NP9QGbrympl1H6ZUTRrHBBx9E3YSfCXdIoSDIMQwP9g
eV1dp2+1DpYz9W7c1AS2epwG85M69iGRviyhdboSNf5giMTtl6IpDClMuOOQGEsFBIuzOhvY9RbC
LIW81cdtkSz/unTllHwjxHWKk3F3CkoPbbk2OZeNPnc4aQqt9a9/SLzUlmKpXr5ycmpNyAxEGoxn
fhyul8Okp4WL5+/pTHbMTq3WrHjOa5EfXecvSA+4kGifjcOKmj/aC/5tvflDqNcgpRAkgA7XcVkW
aGfX6asUIWjthHitcaV0w8HRtouD+g16BxM3Um+w5wHHqETWDAx8Q2iMF+fNwn4S98KBERbES3Bj
8h5OSp00JjBxwbJ9QTvIRLHhZEaQx49+roJRCxPu9wNAaMvvqRyUVV7rE8l+vYpKu8LShE3Lnp0i
CXIcYyA+yc8Rh/7W7wGDRUStCYkLoQGsFe1bzfZU/IdbVrVmhyV7xKD/JM2qXMUeHMWmg3VCoztB
NnmdjWI1rEhsySXXBONwzdeolLCjSbZ+KstsZZesSx3ngg6HKFvxoZZcCkXfO5bWIBYhp8VYi9vb
k+dUsLruwbdh945xE/j/F0jUVkXDIk6ec8VvoFaCqkFvXFTPYeJbxkj+PDTOtz0F401b7Eqz4NxC
srkR51jzXMRxNVs673V7/p7fc1GChjdPaFFwcT62o7WhKi4sKYqqiymOVZPz10YxVC3aySsNZ+X1
VEj1AfziZg4MuLDjdsGiEOxV6dhwJCID5UyEuStB3cV8tLw+ynnbNKDFREsZbiS22eRj6F4jff3s
ADnkNx/emkRl3In9Oi+1pnioFg+43SAWT0M1naJ2D4Sed1aBPuyGVMPUJ5/HEDBvN2kshWJBefuP
M3/x0Blgk93yHeVhQ8Ff1fdRpibTGzNiACeTCRsm2UsuHh23fCCx8j66wCcVctv5Z3PMlCW8lpAB
KRjtdPc1AgNtqA4qOw3hZvNApMvvjolCvBZNOFGdgM0Vgu0Z49EPHrpkw6SfL8dqFR6CiNHSClGf
unoPo3m+QQupXFDqCuQgEnShnM76/qlyQuzySs4KTTW/WDZpZSWR8jZ50LhQxTMxDrWiIbml5iNs
zWInZNzXc8kHNOXR+gWaJ+FRRzvvCaOwpEzr9/v4ycTf8i55RoNfdulJcynJwzUuH4qPiG4+AHvi
5EkAuTiB/iibOw+O59NbKpSl/Zu0S6FoNSsIb0aO+il6nOT3d5hck6wX43q+6TbXzH8gkv3Ominw
wFWboJO3BUDnSoOkmxNyswNDnx9XsIlWvKghdQlRjXSofZoOswTNUVBk2kRMmSMzHb4Llb+nJ7R0
vkAwzTi7AfNsd9asGO+u7rv1gdDmJwymdSQKMiz7m+iBjpaaKOKrUOr20+2HulfS6fiiGLyFDAfz
A5k7kYDXZekedHcMWtINrPN/iPa58nFe1Ai7lwCUrqxo84R9KEXysBiZ049p4F0rd5WOTb5Ferrq
pfAlu3OdJvo1G+5Y7HYOoAPt0o0qyJJsYI/xBrdQMMu4Q/76zSMZYMgSTaccWdQZwY37WZh7KhBn
gFeMtnwsWWym9WUsQ7QB/Ulq03XtJx8REDs96Uv2QRhHtRbiLttvFrr4KL4eGLEzBUQXm5jij2CB
+jVybYjXxAdJhCPHkUwUP+UsINk3IBX9jSFM7vXqTn5Ig3P20cYCvvGUMQG5YW/sGre7NABUGQY8
EBdq+5V6JiqmNV6VdQzGHaQVrwD5N5+zuOtSRTtUoWt7y8CDHwNU4okXaBeV+QP91dYow6XQzcAF
fnJRxtLQeqZVU8w/4kLCqzWy10U5VbDX4f/0MbGDr52e+Yde5sUQT7WFmMaSHuqKsvYNlOKAOU6H
54JzUJXrWigsnQRIJARTJgYWbbHABsHEsNUwfTHl+cBm2NXkiyRqkx9/TjYD5BPKjiql1T720HK6
fIy+dgygk0vmo4Pky+s98/OJ458aVPC+uGqTLb80V4xC1bhWyWAzzSUA2x6iTvPd20OKv77kBgPK
ZUXVCOaj16NEjcuWPLNZM5C3wNncYFtrDhFIAVTJFcyBiwZFF+1J4DpB3ZC6zAaKCOhhCEbe36bK
sF7bXe3+O5lGvPg9rAKYnieAhOrU8fhomFpVz4c+J+NXOCdVeQwyirj7Xjm/1xKBSUs66QUDw2oO
+xazJNmgHK6A3JqYzLtITuVCPapWEuhvYsOnYrthsrCwNJJyE91Xe8/tFNafQSKbWCIoDwIPCgvp
ruoX9cnt7JVtjZt2LV4zyQaIJd0skamBL5b9FdY0mQI4eNlisILKyODEaVNEY/NDH8nfPItuwLnS
rSr4CuEdW+quD4laLFjOsWUFlMbDrMSwr/MaJuNCD3zB6ibB1eHliM6+o7DSQeLy7/xuivzoZ4tq
cZMXUXuL72VVRIrckJZbiKDCjLe11HwgCzTJzew1V80BZOHYSLObRuuItEHQMDaafZq04ZFhffbp
73MlKIJIQ6r4ysLbPT2Vit2a5WLTywIDokieD6Jmo//Km1bQXqvihmfgleAJFdkZkFXDb6HdbW3A
v+6B9b6u/gr/meX+k4zD1cEeIhTUHxkGe+KRUV0NiNi5yyA+yrFklTxZmt45K+c/fC+zbnW1s4R7
Lm7KOucvdXQ/CXqYC3kVoUGd18o3VofP0ujGuImXE+CtLkgE9X9C+6yOAqjWWIlnKVev57ExJl0/
qgW63VxSVT7kjmYrfIla0Jtj+o9Sk/1fgKYCnjChLM4pHlhztNRCUg3d0xFRqz5UzanVJzoTYtY2
bbKyRgMg7y0CXIjG4grL97l5XDx53YX0cjz4+K6eqj9qQN6WdBzL4fMbbrLhEGyKVn1lIYvB9r+4
qMG3DjKuX5nWBoYYYrGJImxCqCytCW4WLMjdn/v3P4t6/wB/y4923Nu0nDJANxZvf6UDVJwwlgGL
yug+mNKVm3bEAe/gxJH1fHFduJ3E34xO4eM/TMlvQUjuaV+GdMLKB5kGYRHv/AGUIbrdkVrjy+Ri
Pxv3Vt3q+EpfUegqpRsqK8kwsygdpwxN4yHP6z+uGojBt4Tz0DFjiddtAv/qYRTIWWy66tYhtG33
KvgmEbH5oPzwpm+VCS+46o2p4J+y8qrHVsDztNLpAc/00ju21Vpn3jlKD2IqP6IcVE/kN8GZG/9n
KQwdlxx440eM57ZmNVWxx2iECJ/PMLcPt8Lnvt2aR4me2JaWC0XeeOeoQuEk9ggMyIvVIQVOAcbW
Ut8cpMEasygCNJkurNVXocZ168Y/Y43tekY8EmMzRHTyGB7XMPqyq39CpU5erYjWHGLCabKUrAar
SzLd1uj0YPtKF40qVIN2GTiyFTCPBbypmgX5BM91VMvrShbePbO0YhjUKFWcg5+Za7JrRZd8Li1o
381tRXDYBxbQYZ6fNOzP6x5Q7/2pk53qOUvJrc6S8LGJwmvYwOCqrvFPubur/j+TuD2dy/OD2urJ
boxxx0fkD7ruSGR0x6SBiHEeZz7qVajuK34D12VV39HfqtSpK3+pw4NcA4mwFwdv1WhXTdt2+oki
YavjnBBe/sF42xOIbeeOG/510KmUaNh6W7+zNC8RtOuLegbm/HhnzwctG3JTFTtdqeE4eCmue3Mh
OtB5HH3tupuDcuKyJNqBUmLRPNI+ToRg5g8r/vekuCkXXwIGfibl7Uceg9Zf/+VNaIz873Tjmgk8
jhhJsEsE5kW2GIn+GUWSbO65AqvxWa+6s8FXSmhge9gl/NdKRRAdC9cEeQhLDdv4sImAb/H/sBnw
g9FVPHWGFxsgVI60kSQwABRraX5tMOerYjbqcYumrr6XfXuefdmAxN6O+GauqNzfhtZRvA2Qf8d+
4FOzJGxo1KmqmqsqCLa7GRVeX7XyqRrggt6vdEWWn4n5oMEKI7nIwmG2WMfWgkziMWzq3d4MGcIt
TgvKHamE43AaNcIeEa3Gh9c3+TEe/mU42XW+A1ldRYlyAaTy1dL5FinrzFCgDMU+t+7tZlL+uQWE
FYe7OWuLco9upcENSDRQ5Wtcg0VHD4tGKMt2mWb7KFGOnYUcTOk6fWR4VJX97/FZNuVzv+w+qY1q
AumJrpQsxWK2jYA2LHaRVdw5Ck8hIT51E3o1lTapu+/Xb+qXchV+1Ng2DWe1NIIwFKgVHXpwTcnv
hXpurXGK2uZkrPn9eC4Iyjh6lhvYbB7iv4zGPCDKvfnXb76DE0Sm6bUTcvsB4yVMWKeYDzsXgm/U
Ptl5Uj2M6Pkns7rKTMC2CYJfaPfI3yVVZiwc8kx7U+PwA5y1mVOJ0oJ3XjKcX0oDQTNfDnky/UVQ
Hz5Qq3imYLu9UeBLopZ08v84QudiiEQV5qv7xG76sRy7Rgmd0Eeh7OEC06y2Ua009wphEPLrxbtN
fKSvJF5oStQTyet2GHDDArjrfZQSR+Sc54SReqlPpc+Ee/00OBNsL4lX9Qi7BXVNE9rx1WJGnO0m
baDPM1aXHWguHbpql1FQesAtt5moHY157j2wE/+GaBciRrIUFFTTT4LTkVRJ64TYHFoHFYnwPtgV
YgVF1TFwi6Kz0a26uCmta0qQIeoDMVX2yQGRrSJEGNjXZtClW6Hq8ES+BAwv6IyQcO+YQDwW4lGh
2mkenTntlaX3k3qji92QYmKPwoj3zAWfFnVs3yvpNvY5goqbqroy4EFlp2prIX5DpT3y9mu2wInl
s78JqQnzQsqd5s8qZr7M7yengfYxCwk/luVUPRJiFMs0E9SyaBDKl3ZEboT45x33bE14kYvLjewv
IFr8XqXyAGpqvbSxQZHES0vI5E0r1YEqxTTDozkHAIgXc8ZOv7i5Vpa2CjLPEXZKA+8xZmvXWDRV
dBCAOYOpt8FLerAJMHjEdUDwyCZejFSxG7vIqBgrMe503xZH2IfiN4Bw13c78IcyWr+4eA+ZIDXB
SLCz7FQEqdbwNb8RQ1AsaJOIL2NYB2iUQ4LOA/BHTT9GUfl3GMc7bMONgD0xmWCOqQniUozYwwF6
1FPSGCK0PO6qHX7CNd7tn0914Yh/W+nVY5IE8l7iZYTV4qpndCXh+6DszVw4xcS2BQfYNaZWBqQl
z2qrAjFIO59hysYQX7rSA2agleORA7AohRW2MK6jepW2g1o7oC8j2G7BHrBQdMbx+h+LkY2vxIS4
37ofe09XLBPvbPAjeY5jNxnRyCJ0nZS83nF0+pH/nuArS7to/L/SUX5nNeEkF1q7jNUpYYI4vjX4
0vvIJLKbeVlmYcWzCe2lkoKMxsXthHFxRAFWLGy7LffBpMTstljL9y4jAVA7vfpTBfb6V4S/Iu52
Vm4MjA2n/Dt+oy78Tjy2RQ5DI3rBFMNDkBRQVBolQftbkpLu7QdRb3AAi8GUk0sOg38qMZtLt6zT
SMC0OPRIfoRqsTsKvgojUXd+d6OxSLzGZBMKVvxLfz3Q+SG6+qfT9jr0dfGwWdUjAEyYMJkAMUqt
5k+w18KcVEB9YPkKvT2o03DPykpnvcwfqKdSp8ojfn2s+o8Wola5bGutCpwM8BomqNkDaUvsIJN4
XOsH2gN9Fps91g7+T3qzs0lXdDcKOrn3NVIG8E88QQI78zBgqiBPqS1mgnCT8y1WJW5I3jUEd4sl
tTV13tABR1Rf2oD1UgNpZ/Yxfl5L2F+AVwtrhHv8Uy1Rj6jDaBrsN0syoFa2dFgM6BFo8gg/S7Dx
fEx6AfwZjBS6rnwW8azWLZ2fjf04hDlzO4O0N5K8yprrYnL17VlWvY6v8061PQPzaCsqThJ8dOsb
yefsKmFVSIEo9O07pu2S/B5oufmnF60uoya5IU0YoidyaIE2uKo9KnSpoDatDpJak5Tp4ggO5zWd
gPwYDHi/hsKhdklM1fp1phjULocF9CsU3Bh/xeeNwBPeZFmyKfIzbcs+96CYqgfI58O9++vz9qgr
4l+e19+kPHUnLNVH6LQmm1XXTtRso+cU9s0UjQE/Jbu6QFWRQb04ejCQcaRRDSoJDNWQPstkt4vM
o67CHvh3Eo9mM5im4EY6leHC73H7ugy9SwSdE+qwx7oDV6nxsNnMg43zYdf8+V/7xRMwoAufDgrL
SQ5HIZAk8vOlFnegvS53Fa+OcauBaK0Z+CDdPpg2Uw1ipQkAMNeV1iDPHt62y1VEme8wSsaPcsgN
0Htec3OiCucaq/cE2zjXK4B4dJ7xbvSZUJc9OLp8nrAlxLHi0h5qH536PwOLQvuRRTMvmWek2exU
ICYXyUqEPyDJwiaoquM4jy1uGnleqBUU9vYYRJP2WBzWngNpXWkt33IYwkgJbVH1KDXVh4htUD1t
8QP9Qcnox6vO6TpGqMW1ldbC0noDn5KYAUrLBblAvc5TNWrIWHvrpiznrFQcz4zIHf5iJssll15R
rGDlDjRgkJECiNf6Q+wSadO9G+objHSFq03EMYV1NsaJhc7UB/4jJmQH3X16xp2N2dLcZOZZy2L0
sF6fqMhHUTqrFKVEtPcc7k4WGQ/dTxeJ78Gl7FtpBRf9pTkqocEv4RVA3wPZ/GwimyRRLG3JZ6qt
sgi9eq7uI78I18DFY1IMrJ5TzKOMqc9I/UYYyAJQLSkmDBwSyQdTeUoDyhgcu+FpNy39tauGosDn
dZj9YB2MWrRh6TjHNf9cCavKxnW4BOv81vHnRZlSQfX9sRuTPSZcx3zIWsswrCrrFRkp9QmclMjj
eT4zIYrHw1EMjhn2VqMHxNvtFtDHFa5zblMBPYB9Q7yxME3uMCU6R0lldJsTD92JnkOBz4S6b2Aq
Ye2ZqfCwPm14EvC1iYu+Q/KL2eOXtH7lP1y7yDzGwHgEtfLnTymG8gtRJSR9E1dn0cTmYd9KiGTD
4CmKOK3Ujw8aIWO/d5GEpycf/2puk1SJwdG8xfJlWbQALXU4Yt+4Dp881b/BEp/s5H4cKDGFF7E4
pxT/iv3Den+FjLdr77iL0XP5Cu+L0c99LDovISvBz3zZBlmEO+4Pp8J1KM7CBZIABraYo5NeKyBq
YXiroPAS2Wl6QPrn5WD41Lnj325F4PkMcL/s2Xf9ByA5iGTniBcZouBhmQOxKHgBZs67u5ruKl3S
Ca4RxYXaN6aWNByq4Cjuj30OHnBA+rs4N49woGwpNeK70Akjd1ZsxeKiUVS3MX+YjYaCYwG4w/Ns
aSSsgKUAagv7SgqoO1X5Mo+ZuIOOeXK1mreo6Ly9sCsLCbFlH3qAsnOG2yyfDyP6btZ0T5MytzHf
9m0tjfrfc+HncRqrXggjZtA7GjbOyGfpD0zYqybtUW8yzibj6ME4VP20szKNVhpubqYIz77tWmNz
T5pHnOETSlVvzuQb5/bndMpsxHeArA5QGc/Q3pyaVVRJzuSSyInso62Ks3ZZv9e6/obfkAMZEtCn
zMT68m+0Z5VYu6H9oN0XWxVeB8C1q1DNKpsND897Um+gGujep6DHnAV8f4isSIbfPxvYGJ874LOD
9/5XJS0WhMQ0mMZVBJZGMNBnBiRFk6ncQWRyp7Pf1XJh84EspH3L9H89JcMZSnGfrZMN9GbdZ0Yw
3nWt9hIkvkNte7/u/hfO/QSpPFtzy5G1fPBMuG6U3ORlz1RcYLKYItk3ad7QptK9a9UOlNhlnZIv
DH8933/7QCDa4SG/1TkcrJbNMkb6lF9cCrUJN9fclE9vlZV/vAx+ODR/Pe4xfb0vlSiCWE2GB2C+
fH8y5pe2UadUqFKQ6awp8nHyOvsRkE+vMOKb7V9a1mV/8Slc7DztoZi7T5wamEcP23BAshT0+OAQ
4pwelcaHNOoOUXy9g20nzcWrlZGQx8Zpu8iv7aNLWgyCHUYMC4tMG3wjPj1xpK5nIFpREMEicIIW
H31WZ8+TEfO/8r4XmIRNns0Q4GIadyLV/ISuPqI45aYWM2OmgDEoGu6hvkdHQkcHBkQlADpfZ2+V
M/18BS1vru0ai0dKKrTqc/ElO8Vu8l+q1NsvwQa8521DRI5t+w/+toEzwcvdEAOE/A7p4WdujMA7
nPhKqz3f1CkFZWBfkCtJqIt2m4UYczFk9G3Hwqpr8RuoXuoEzw8a2Hm1ZT579+tWlCc8M1Zr356Y
CoTnPKwnPAZqxDiFGOl2aJhLJezrqlGZh1r7dSUORz0KGQ4SkTSHyVOxWiw83QivKTZOrJB3DY6A
aRAHlbL0kuX2duLnWt8YDoy/nXTHxbA4TisKP8hlBUXpZWWFPVnglZQ90IqhqIiuaer6Jf3SHlq5
eXfwh4Dl7XjCOok0x6ES5G8pnl7k+/aJuwOvTdMNlG8LM24HURRxErzl37EUKj+T7TA38GHJzDIU
IxlVwEVIGOY/2UvwSGeKpHFdqw+bNBLhYhZ5b1sGmaqLq3rHFsvjUTz1am+jc4lazSF1xLfpgffr
mQWLwF/KwiSX4AuaX9kWIKKYltc6hTdQelKv6OwVVJtXmOr/PrCI7lPsfCqJ+QdhonB1hhXMaaRx
W02Ji4nwKNoSRQz8NMqK9wpEc4/4UghO+l1zqY+WOLNpeqn0bCxDz3Kf/iIUuJCTpVtXP2gk+rjV
ZmK4ADVp+zDOMvpVw5EBnmXN9IoQga5alqzOEauAsKuQ2gUyR1z2tQ+zqhCqCogDDifvsjMrQIbH
NOnyazZpqDjuqhqkyhEG+KbTxFGwt0JsfI/XosOqCtv33ILuKg0gMV5o8/VqwLriIlx7nct6WsAC
w14VVptfC97+OViBZs7Ot+hKo5LnPU4LHHbVBNIzj1gf/r1D2dDeo8JNGK65KhomBH82hrtOfbEz
yZ11AJOR4BkWZYldRweZGzKmhSPGgKP8RKqepUSbIVFrQCTxyAPrxNEJEy6DLYYegVo0f59hSzIY
2t2cyWjACVEoRzWtsdK9ZdaNa9tY3ZzRt0ys0yNfjaGEbjHcoLQkYyO/dbSfgo4FILbT3JPKD2MU
Lm5zsnrJc2jaPMMBygnOQLaoGgWAtPnYnGM1wG+x61IFlp3gxwZSaeZ3xIDqGGREeUWueNXWdLUp
gUvoF+WB6vQTNy9bhCvbq05IyOa/LTrkM98jE+DLdJW/CEkp4u4qr2mAdrtv1kSs+wWbYaAt4ksq
9Ix4euSFHgDypxr9jQLKgOX/dJhH7ud+jB8bracIMZ8/F/noeDkhwHUgTtez2HYmDIz61UfUrgBq
5HDj692vmR4FPQYHC+dL2lVRr/Uqtu4BRTIhhPS4IFC+pgh6DzpOr/dhmrdMrIQSmQa3zyDLTHiP
pcZ3qexVmfbcFsEQIGpkezz28yAvYrUtyZen+alXPaXKGJlpvNJEP220cUWzDUAdcDdk1xn0ERaS
HdCefa/z4CTxcKjWqc4qAUUzM7+1rah3c55/n9zRm/bPiCAIKdxtnr56MNeWzny9+RI5KMgjPDeb
VHMjgvON2KUsSEhEzMXp5PfHMxcdFQE4ZBwVB/5W2pnMuJwfsgbRxMqTbrVHwcNKaPZJWs2YogTL
BCPJV6TVABQ8LW+WvJr2zL9/DnshGHo8Tlax3JRu7gOPE6TQCconKrio0tDdpnUJQPm3K8mFXBxd
4AzHiAHwRdIoIGGpw05AehaQRMMlycLPYhc5oLjXAUfdd50CQjvyyr7UqTcjwcoqBLj849mm+Z/5
h0y66DZQDbzipnsAvVtYcGWskQM6UJrXodx5+Rojxs6MOmK05fAt4DhFWj9hl2J+6VwRdyfEkpkG
vv6VzI5ovVHkMHUZoDdkN7/esI3s7zBZ0TbKcVLfULUMtqjNhjuWMQWcElIAPsUqSyKpyoNH4/2l
1fV1XkP8AGpkdYivKdZy0CMbgfmi4l3XNK+BLc5qCyuWglTRBzZ+KcOthxsAlTjmLMhGRXxemwQa
/uH/o+F76ooxKNJaYsqVPxkdjo9Ll5tRyPProILraBjSFCZlZI1ymUtxSgb+/QkhNa2WFM7QUPUJ
p3kIxk4kHO1IR/MNiqoGNA9aCR1eoa7RLIOHEoDJZ6zHyZUq4wS8WxSgH2zy6VeP5d/T99fm74qc
fo8Ux5zRqYh4EubEo2TLzZknUFy47qHVuhth2ozxW+9YavZT+5UWchx9tJcWH/5XbPe1pzeIU0QB
j6GaP0jElSNSI5vMlRC8i9RCVRhDPcWDqu9KKVO1NK4E7dPsRktpFmCln7zFz9Fqo3oZwQZPqfHb
p3YI8jrPwlLfuQqeLFnKKUbEtsNzqTisEjSYzygMRNu603f5TpLoAJOVWFK4zxbgVCc9c6gHfTbR
7exdidTMlx+MmkAgYcsGdNU+cJu3MsA1DmWfhzIX755ke36tebZSW3nYtypoR2H1bXJZ1HD91+0e
SlrlR0p5sb+AuKfcnxESxVUEo1m0GkjP9cn6XFL5Of271DAHs1+7b7sZd78nu76LrOdUsY6yCzgw
JcJ1sVpJHyQfG0RLKYCcwMlhGa5dKo5ysHfGkhRR/FQMQkfyktZ6lkwL2PvcoTohYbyl8Yc12ofx
cNaL4ce1Os4Cy9CC1C1oA+tUSLUKM+rj0dr4xGePz/FCtsIWFp1JbhVgUO4TIMPONzi8Fx1UutYo
d/ubLN1eINQIuqKCbWDr0xnLDfmDFhR3dJK2Elk6ZV2YKmu89/cd/ssXCtEIZneHLYEGM37CN0Wm
oW4IlbcPgi8wPUZfpCW7jj5n2QpDzo+j2IftFbN+nP6UdM8m3GIm5Bkf+DMsAsTiCwTLqKWUYj50
yOZc8Ys8aPXNa9xOm4P6kWU8PlSNVZLrzIEc7HFnJ3Rk8MscEPy5eSeEHjdM0H3fLxYMAnTFdiUq
CVzlzrEswVnOqLbebOclzQQfWgHAMiqAqBLRnMEZfoSI7UUz8eVyx2dnNIgTgATbLERyOW5XZ+x4
1ThbHfhq3SLpsRTgG9Ovnv+l7/OFbTJ2g98Ynz5HqcvDz1q1Ky5q89UAY6kqtoZQsNMXCsOmEDBs
5nqM7Q1Fbn4cd0ts90amnEtr7jDho5mZxfyJe+z9j6ZcvgFd061eRO3GqsAiB0LK6SvukrDunZyB
7Nu3JiJM4naAIV9JKYMrQsY8gWLSdqPChOhY3+Fi3e1KvyJGW/UlXXKoZ+ghTMOioTvVotM9JhfQ
Jb1GpjPSG87bbPU7bsyNQmjsd9fgtAXcE5AfA1YgIk3iHtjDwbYZAPwWD49/BKEwGxFbnSK6dJYi
kILicTJ3UxE0bhn1ek6lnSvxxNglBFLzaowzIvGsAGE+UFAcYEGKSXIueE2H6eEiNkFe/5wra0G0
H4lHmb8CGje/CNGzvUIdWTs31+I4g3g2Hj0RQvfAqjKRb9clOw3pnQ216sDu96SWLF+KP6qwNX67
cL1HoNvZWy+PPaujUVpP3xqLiTZBO/yN3kywRRw6B7cRO6dzK/i8lPNECiesi7XwYTh3EiysG0qg
9zs5XKcEzC5fWEjASCe2HItG8DLh1ccu0LX+omOCGPAjwwGS0gKG128bcl49a6FW34+SkInIDpK2
AZG0NISzG4Ls7uQqBQrcwMLWGWTVa5UFfS+OfJCaUwJbmHtEm5HnLhQJvFxV+mpuGGt9lA9PS3sn
u3UzKk/gCbvBnlZXNs0Beu66FjoIXFm6EVrnLnAKkNSflFZzxNWIBgLX4829L2O8fb1z9EaVnZdG
l/cUuCEqf01pmzwZJ/Eo80PB+1dzj05D21nN+qcYywkNSfW63etnT9RnJS3As0xznP0luqht2XKm
xvCaxuaJlIxlLEg2rmUaXra1bogtNoH0nytqqqsguuqIfI8FlFPvo0RaBkQeuQOFurWDZJO9CyIm
mSSVGi/4nIMWAgjQS2QKrAxnujjVv5oBtt8KZQKyc+48z+WSqPLqXWKkxt/uWzAG6JRlPOmILZED
988dPN1lghi4623zPN+Xt3kO5VXzWlL5zG9Gf/qdNlHwkzA7k+pbddNZwRMTgr+bIVAJFs4ShhMJ
d5Xm6syi/Biu4f5T/TrvFLGYHfNUkxK9m9DcwJ2w4GKF9mgRoBj9CJhesHzE9WEXYN/fTVkvusCY
UfGUvcLb2ynInE0nGp6WNijvGRb3IcR3fbkVWxUvR2v6YR1SpvZR6AjIP111XYF8D6PJOM3rrP3f
DY4Z5csLtGnJ74rYPf459gbovU5GjcUzPgeNklvo+bYPirmSxXMbqv5TM+YRKRxLGV32Qn92kpJC
K4XCl8WI8xsCPejo5KE7iZ28y1D6xqbxw92yN6klCsc+c26Epd6XBRrUKwXP7hSwNFsbQ0jBpa2J
zggvqIXpt4jXtSmLDkEDD/lAD85F3b2eVu7GN8Y9ou8zki9AmUQc1V7uIgwaVKLvuG1OfEDycwo0
QAfZzkD6zPNvEorgXvQmOpICgN/iEZTHKpqTomnNY0GHfz/iH4912cs2dCxsjYs6sW46gMrjLYME
E+6vmcH7xm1Mc2FK6HIl1b3tonLZaNkkBDlp6iGiO0TMUlhwiBfxfOnaInLYISrVlnPaHK1fau3I
63WVageWTy3FqJhPKbRRux1fyzF+4LY7ZT63VTBjauyo0DIcbbrq6xRw7aSbsfTGDMeBiHbVHb/B
otDASaCKzx6JqMaXCAzBDZn0ypOcD7TcTcKp+UF1AuaX4VgbwqwP27FYkXuwVp0++PXJLj7Hs+PD
Ex7yWGXuonqe9V5vQsQbpUNt6zwIIYKSx9JatGaObBip6UJMcGABVWqUOZ5kQxfuwtTGYu9qCzKN
+hMMhZ84FLcYfRcMd7LSzWXHmuK/en0J3+JwPAlXOeK85hVZP5Od2Tnx8xQC65YgoaLQDumyg4sA
5LNFKEbDmFOuK1tCl2Tsc0ariHttTL0z9MvOtYgfMjyzQS/dPGni/5JCtgHtFcfBE+kZsqFk6L/6
r1XxuchYkpzCQLOdgEE+vt+2LXVAmSIEK5agg3yteA9kdunYl5jRsk8npXSgT9OiWmJ33lS+PDHT
lz0eIxtqpTFkvxLXlvtfXwcWL0dFz7T7xCBZjRxCh+kj1G7sAdeFiy53sRx9FEEE0TLKwAnow1OB
GUzFOTyHFECksBsvp4tDnGd34HkGIn6bIo/TZB+3GimVRI5Xgc/TkE0TPhpUXKTdg3IRi/r+9DSM
n+5tvi0UpZeo+Wm1fUvhDklXrGjpW1SEdZ7ginm1KB0P03fycULKeHYSjqReR88P44mRMUW7qkLS
oMd7aeK3Gs9aNTepvrAtMfHVz+l8YSu1iZoYPeYc3O2m4LWfEzgJXFjuP8mpwlCblGEInzxNhhWe
eSiCiHw1oezK55sXArE6Zo7NXAy6tflarP8GNbCW6dDCmznmKVVC+QOQo/Ap3eXe5bpYoHMONOHr
7rsAu64EAq/t1EiUl6yUokWZTlt/lGlZOVyXnmbRcnZizO39cOQ0amRrAOnda7JhNTvcX3iHXeno
PE7zLvyYonP6HyfW83hDEHkn87Ct+dZhBhsXvzR8chLjo5rYyrgeXN36hAINNNj5KSl7ReDyscOB
zPRLvIaBuBZTFFTFOHtUinuWFlhxygdvTNYf0M+HRLu6yEo1hthOjaTuEPBIXya/m2YIIV0i2LN7
DKYQ7v/c2sSBgIq1US4iq0dtUElMAXRl1cqmC3OZq8hrEPfIBbSmtf6Pncfmeo7+2Xy7Z7NkUx0b
VI1l6ifHf1bHt/zLDBRkf2Y6/+a6uxZtRaLwcCAQP+Bs3ExnK0VcEqD0eMB9y3xIJyCSaSDi0niO
Edi/vOaDrB+FIE9TcFBKbPR0QFCmYaEWSZdwHtNeZJuvHR4Zrg7U9rPWqSd4DauGGOYnia5WgMZd
cyHT9Lg/BHNxX+gryoVZnNTxveOWvJN1q80v62NDjAbwC4xTqMiHILeFuZuGZC49lOx8sNkq0fiD
/4wjEptj/IpN6XagLIyTUb/9GRG2Rj0oS773gLaL5J199wuDiRsqqu4UbtuZQyr10Z87lvQsEp8k
B7ti9AYwzvRBMXsxHRhc9EhQ+E90AVWWr5mVjT1BpKCEASY5c/9AUmt8aScXDd8uU/enfDdkNjoU
iWDceJGQaxaLT1UaWXQBqQoqS4eCfQr8wxv18eBngeNFuv+PqA/CkRCqXEEzuR8FR0Dr5VwFsTmu
Nz1+GD3zFV82VH+e0fTGRX/comA70MvhCRkwwsa8RJ+yLHTG00wC4YVDahRqZnNJkp1HPvC7wqcF
u7s9xX5gVC9sfTMa5mzuUg3n86auYOVDGHr+nOHRS15runwo0gBJn3+pdUiieeZeCnkwUe6t8kcx
gaB9Zf6QxlXvT33+5jvKFE1RH2wgVqWkgvwATy5lJfJe/qyUTImArtoQ85oUBwVw9Wi0S2oLX7tg
MgLfN9imgkXttAa3AGuxTHe5He8K/06k8ylRCk6jqf2anxTDI+ghnXycsx0EJLDTBhJsJppNOIhm
/I5jb0wbnwjimk4SmctLv3lK8V3Yuro/NbgisXWDeZdTlsy+QSdRZXI96G++nxQog/nQ7npH4fxX
w2bktJ5NyzoVLsm3ACIUoO8sV66CwR18bla2+ufFpfsBh3NTblt0oNx29dQwezdrzXCV/8dakdCc
/SWCETQcL5/N9/7lPPlQz96lRthD18LP11Sl9kV8XSq5usM8pFK38OqJDRGlNCAkUJgmxIPi7+6O
wFAAt2XGVTBFqlmxIhzb5hMsTsxxp8w8+VJavyv56aUp/X1kd1NrtvI+zUY2UttopIXoF2eIV7RL
J+2MMcTH06cBL5/wM0BFvw4wOcRNhO17X+9M9vmStkmFJttRYsqFJSwZhnS1g845/eiGDYX1RpEE
IhDnZxDB6CuoEHWSnEDmFD/iR2RkvTx69L84VYNkMhr9NY/rUNIIbh/5Mvoqg+3pu93S6K8WvN52
AoyUBTZXcO5SPIlItdCawwrGkATnvQz4DtJHUhKhNaE5eVWf6dgCfzWh+nKDbApC2aQFipFKwlG0
2xH/64JyKVgWpU1hCXK7Xhyq24IaqMyBoyIm3Mrd30LkVhO+hyuHYKdqr7OA9xwLkKbqBnodBA7R
YQXCtCeFJT2aaT6pOBemCVGpjm9xPvoanxDIY9uN9jLdKJe3/Av5v4bNDpFg48uJjP6c+9eGAS+W
soGUIV0iKFz2XkYLIYqvrfNXn0UY3R45e8hUrXcaVdCXUu3q72h/P2u0HgLg2vzxyaP7HKnmQBxN
Zo5jCkVjWOB1Wkn1EqxnBUGKrL/VWPxv/Xck04Pfpq8tL5q60cuC8CKnHaCV7DtcbQgWGlfV1Jyh
viI/Q+DgGP4aynK9A77IMUOd2a/PFuwJxcHCztWR+vfRVRwMF4WCbMbhR+weGgxICKG9QwlnP4dA
F89lxx9muWan91bjxNdPaWONRPfbFd19nswHOaDw++TMD+TRTkQ1kVVT147ksVwweGrD6TMPvf+1
Y3ZJujxSy0geWbNJu8adTkaDiSbu4qZoxiPKAdFnuSn7QaUQfzQwPL7TeI8E8O9iNLna8BWUzoA5
fWbTzsv0aejJYw2Y0ANlGA2ksV9fVofLj2Aj+uMQRIOL58fJwYXUTFTnu9KV1OqPDdmRvn+RfDVE
v1tgqmqV5euWNoHDDhLYkcCgrMQx33SqZf1ShuIKD9AduHINSd6HTE+QrSj7TRIuBg5dVIjbj8xO
p17IF/5sW44VtXxJOOx10MxGiGU0kaVrvj9F1LnLEeteDiSYL8LoefCNZlu4dv3y2KbXlRqQJtbr
9S+h2l+zOPJVFyDL1Eg292Pqo8lwoeVIVxdMaVU+32egz0YHwoorWXmdnVXWPK1nOaKjU32CvvDu
Fy81rwLbkM2jh7pEkDTeczngzjNMdzEclNUDLGXDjFyZo7yWod+AGhpSOICMpgtA6IEi6qtse3aO
jb+oNi/DN7u+AQum+7ZA7AoRNnR/MdT0bjw8+CnvN/tgQjwweq+Lhs+PeLzM7AQNIDyW9JheXGy+
WVSotbsPSWPcwDwYC1zutWlq6iWbcwT5S3WbxCTQdroux//jiwcH7xrNeYuq7E3Pp8tUJwl4hhYU
gAnXMEs/GdwbvZZauiPSRHmu6pdBPHYrJfhNFRuhTAEsZ19w8kwisYkCLHc8oTcS4hxz8D5sKr0D
wBoAxq9V0f7FgQv5R9kYIOqAd3/NjqWKtKEldUb3afhTo9Nq+BcVxkld/q5yD1IGC3n7NLejuH2T
kZ96gslV7rE5qwjKDoishzVWM/dhhuzdPKDrztKB+w4N/hOEDL5N/C6AIwuco7VdvjbzllqhdHnU
qnCsUioCtHHBNhzR5fWqa8u0TOQtztkef1NoUP2/RCGz1lYlGspeh//p04MSXcIH82BlPhxm8HH9
RhuWHjs+0kcvjy1F0heU5o1QwcYen/Y7G0qbtU7yv2fb9NCzLhO3H9ATIkISN3zjkZOOJYsltNjO
+64K6UHaiXic5PUlOlOM6ZLaZaG+gibgt9Eofq/ssKvBuMsm8pclVBtcBtveqqxezmXNk7zRWJuU
dU6Ii0nEsWdEDtiZmGtvViqC8B+R+MxFcQrG9jAQhV/jiQzVolFz+pmmpQZ48LUxbtOHMl0ezVto
zsN1/I3JqxOzMOPhH/aXrOwB+Zx+5w8wJKmlnzUHxhoeHKnfscon3BYY5O7izZvT8SAm1BOsxnhm
2fOa6mmL7a+Rztsenfdfn0DSPbpFO3XzVHWmNaBSfWenYOtuS5juA231D3/kHgoXuLKQLRPyZW3k
Wf4qz2MdqRTcYrYyUPSjSLJRmFO3nIR3qaVHPZ081RfOtXyhruLxMLY9New0srlvv+q4+glrLlZa
AKxwcIPuLugHiCekBC0cGNQFvJ0avqxxcxjBgWavDo14rs0kd4a7LZdYpLpw9GNP9L0JjD3ggF60
nW8UVCLIeRE2yNRiadDsFjw2r3hcmBKPigXPqc9Mz9BUW0nvx5Xkg5YcNAw6kK8LGfQDE/zzbjS1
AkMfbdQjOmTG7CI8NZcfIBDSoau6e4FpRYbqwGL5dCRknsN3kZG5Q99PWnurXyK0+VXmrAZfZUpT
fy5t+EhfZd/mgSEh7CKzj71UzjHz/uIGsGWDvGQF8EFrOjq4yl7dTcdPT9HUrMGYExS8YGPQuGMD
iE/nEsy1GpRECg8FOvSjSBQJJq8C1Bl8qkBLuea97HQke+9SdE2YGMC0AC8zRaeTozDOHZ1Bsymo
rCj8+m8NQhJDyUDlj3Q24549g6hcfLAya3P9M5/IbA6iNk2jVUKOVabCz1qvPqmKtjGAAlnmDBYn
yCphlKDhWFn+yx8GXsoEr82okF31ZkScUsS6v5AcepmtrrPjtRuXppPXKh8HOj1wc4ZmPTMmCW8J
rqFtLU6zJ12gjEtcSgNQ34mRt+rbVpDJIJWRxo6YadGXfD8jTfFgkWuzv+wIMkjd58+QNyekJ3kU
0y0Pr+ixJ7KX3pLrlsR8PuK+s5WVqV49MYrXedZ4sFPDOoc8FFMQFEzHd0SEs4Yyk5JWRHH7Zlez
UrrDthY1B0yNIenkk8IY428vBOuVpK558wEY3KyBx2L1OCnQfx8+5/99gr+kY79MIkGhEKJP116w
LRXGKQ0UsiGgmyRIzzGnKje+LvTQlZXttg60IjtMO00+cxzERIQmmjEwTeppdJM4ZgRll9QE1vNw
Q7AFLkriPRSc84vVcZgl2ru2fPhk4WJOCpkmI7fyqoCl1/6Sh2daBeuhn2qDjgd06xwI0DX5st8Y
T0yf0Nn9PiGI41DWUTvu004FxkSuzEgw4B2A7vmwUGbt3iZVWENeYTtxSsfH4KyrWUsZO0ft1voo
RKRPGaiwzoamXkEfDLoInK/ScjMnNuJMGBtOLZih34ZWJ6UfNkidvgWzG9qek5JUzKJV2pf14BS2
GW4+0zRWFfBMSUcn+GL/5pVChZPDdF2abuUTylyVxKxjWGOkCM3rEWN069gvi+ovR+5tLkaorxhJ
4SOCkOr4awA4bbhk3iMvtICqRjdMyn/ZxwpYZ6/Trh2nUz4qeJLPGFBwRcMhUV0+UMu7MLPH4P5p
rx/N5IigkoDjmlCbz0Q+IA3VGGz+8mNjAOhKZsDyw4D24ZSDq5Uy2DMEszQaFWufGwjyNg0u1OiD
xA5Lia/IDhHJNDbvfqlNuNFql/OMmTtmzTAbEeKIAXtz7uix/x7wRuRNIcJN0qgTmsIaWjB070jc
coEkB7rUM9Pq9hODTx0E9OgrxGX9Au6Cg6p4qnepome7rBPVDUfWpFHnqRXmnNxOQGWxH0yszqpZ
5sUCdLwYT2GyjYnB/NR1arMoN3/5+toD8OqjjFALgh7KhCVtRCeRNCXKMlTE+ijFzbbkxW7eEwtP
YTydD0LUH6KUrgBpQIsD+c7+8gk/sAt0TAKi/OdTu9JN7nkswuW8r3xQksyeFbzfLnUwIi+ISPmq
TfdF2SNVAIgWgvuQsKJGx/HAUjrRufa1h8Ek20ofUBDDfCWHjZgIS7KrtD7QlO3KZn5F0CiGjKb7
S2dGzZUl1qhp5SAIXm8GFhpGhMvWiG7VTU78PK0QSaoPBjvETM+Z6X+GmGtQXOHqxEXjZTU0BvJt
AorX6B1UCPVG4Y90rmV7rpspuwqcQxN9nFpWR3ymygh7dHJGN5w/AlDQdHL51ToMj6rHTO7OPLiF
Jp18RM0rl4qtAx5R7TryHn8EU4Y6kNaSe08VEH9TcuRDUCFHnE+ePHYlZLn22ZheyBKI+wMOibfo
mSAjC+AbhJfzvw+7gOhPGaVdokzmD/Wc1l1hXn4OIrm0BDbWWS4ZCA0DUU/Aq1403vgMMdKY7nbG
iRNo/j393oO9GNV5YehKFsDcCfhj2ZjI/2IK73gipMkukt8KzHm+vL2Q8VDgX8shyV7biCmjLIzI
CCGPOrRRyi3oMLHYummOJcs7Wr8o7j8RE5yZ3FHbZnGF1WLPx2LhMLQsB4K8bhqIcsprOmbQ/Bq8
xXm3QSk/gr6XlP6UFA5jFMvkyKo8LZ2fLeoH8zhRc5mE54EBRhaZli4k4uOqiychFrD4CKkD40yy
AoZaitKZ133FlIRRrDG8TEGEO9+0lT9SsSMNBcxYz1MP+KkI9KFQGqoQgqbczxyF3p1QDhp8XFx8
aqV9X018jSfUO/I/uNLpekaLYbtYfclkGb4ttKmt3fq1/jjOsh8bYNHniZUr7aCkj8xVvi2E6X5Z
jqcAyoGBqqpLj5QMMyHvHrHSngF2JVNWbNUjIbSCKYP38vfrSW9UkiNdS/6KIX441eu2QspdCuJe
mWqF6QsBw0aW4G43zvz2FTtgJBFwgT6scttPvWaUOSkJHQEXk7h8IR2gFhHN+cZzItOeMW2ZmI6o
xANt627dlOtGmuMuNg6vkofD4APdjBGo2MTE5eDyGAPrvzfUBA/BRhWxS1cIU3XswY3VABQHX4zg
AoE+6dwfkBJn7kPz4WIb8iQeXg+okUk5z63LhWAopXqR+qScJn6N9Of85s/xLxxgdr0KB/FHRhPu
rmHseJYwqPaddUDOOeIRLJNj1ZGLeP/e592m13t9PcjtDFnaikNwDZkg+lvBUyg2aD8H/8NbYsP6
sjIE8gDj8z1SZrqUssuy6cz0kBjjjbnCkpLGcoFzVbxLLA/bx8qzkaqyttF63ZZ07NbqM9wtVXJe
d6zMExmhAANjZdHjhgR+fgMAKxguufw5VAGWNLlh/fekuzIb/O2RvTwcAS+3dsHH5JKTySNji6cq
H3of/4+KsWJab4udBujvPa2/J0zSRgdn0LYO/VLW3vTEW7skgVdDrNzAldXJlNgxES7MUro7QSWR
O8RUqGBh8cpLb/mXWx9qOsziCRIbimCN9MwSe2Ujzu8ERFIzYyQeLnvJUDA65WhuafwyXonGZ1Ol
OCG3acRuqg2tX9XnU9aot4NmePIDxfKevqzdkUy4Si+eDonATwCPZAmL6M5BUqjO4OIHhD/dHLUr
RIRRf7Ly0gR0+CecbYBI2yo4qWWHKudVZWDuOnsDzaHOK5WfdNTsa0j7n3LbaOaueoQi1a96OUeZ
jGcEL/SGVdq2rNwpWqUAwAX+svlykHMgrPd/Gi7r9OnA6PEJGxVH9MhIHkZWEKwveTamB4y1TRSa
M3Z2YmVWUVGnJFv0Z7hFH000C3HciqFaQw8mWhrbM0djlteGXN6/hoCnuCZPyQubJPoVrfW8kxr+
o0ro7915YTMSudqywv0lZ26/Weg6aO+U3yxB6hv9oL+2js2wu4nJaoySzlJ/IitA1xani14NMEAb
4CcnFqxDexJDh76fWWSUI1E1T06l4B5lhzfnLMFQ9r2iTQQ6bUdGJtS/WW9llIcBg5HY1CtZiutM
Tb/BssLmNDKjvoFBXSM0m0CFSPCWM+bbZXRvb1KIgKUT2PVkdDjev66rvyKaYQ8nbicbKsU6N3SR
XRrPsBOP3U7V5xc6lVrNqH5xAYExFHAy0vFwvAHMhunlqHOehXkCkYOQQSZvLeIkbWPx1C078uuS
PnZ/c9Tv5LqA2qgszchS3J9OdSqPpBkpr/oAPOEVV+93c00SS6lFB4lP59ANJKwU+LjJuFHOxHUz
o1yFchP5P80LQ9/onGPtJpVyqIGXKOkjDH9pPDBi45m6/cH3Aoix2cNpyK/8J7Xob4s4o4dgHvoE
+uiUE8ENb3TdM4qUZJdxYmYQ6vWu/+/w7/qgOBCbQdLA4q60RVABcj6Q4FoWXrXXh+um3yXzx4DK
hKk0Sefk/7tgRC5Run1vJ/pOrzW5MOutSmq37KTDImH7fkK3Xfy22zI2xZCtPIBWvQBa78ePSoEd
PzNVq34TTJEReO+cTvGnLPLz46dFEgj0uZRZshJSgDEfsP9NSiPcm6t2DUro9yIshakHJgAc8Iif
aTSMbXQRD6Dy3yiCPIOC+j30iEDRZ0TRavFeDIQULZfSOnXI+4MZKqKZNcCfWetXAUlTZYSfAcoL
wkhYo+kEipaNPVL8JZb7aEo00/vCB3LcB2NYfJfPVGSGRtUis2TcH/A7LGqsvJYxw4ajBJueYkGo
igM8NcbWMNcIfcXy2Qz7l6OLshvvZwWsfyFlwEmHb5Vwrhd5DMEh7DEjPIGESw/yrGC70yt3Yu37
xnFSikRA6nk6tnNLlfIoCkmSrO98lYYinulfkooYiPgmOtnr3ATsZ3vccIPXeA/6wNnwQVZPgUEO
bxJuk/vejkwEGGXPocp/2e1mX7ZxPkRn1nNKEDFhgEVbcLnUJ5xS6iz4RdaAdd844W/5lL83aYvs
bjIrTObGv2CPl6yL/Ub5skl+p30ROnE/wg0Z30BtVd/zW5JAJeYSMDDSTbTsZmK5Psxs4q8PxauM
mCVRH5N6jUU4cwwkwbHn0sR+1K5F7UYKqR4ByJAPBwdtSCfzn+T8N3lLJzIWjH2hEAkOhKt06qYE
szgv7JG5pzz7jGR9yiJEcAi3Ef6rqgLXnURmfmV54YOWenlgaB04qMpcwTqZitFB+34u3J3SNNg2
y5UmceefpnF2gXa6ceHGH6RSfsWO2JvJL2cKFMLMko44U6XasdOnp5SUUuaWHPpR5vC0TqssAMiE
gWy0kxnz7zymrK/ib0iDyDGB2EOhcZcYQYFfAr8XX6yMh4VjtyzZhz6lRrfDoL2U8PdeuQEjZRLt
5TDfYeZMxgsitLQgXKO+lWQe9yYop58l6spkgiatTLS5APtorm+YgpbJxm9YLu9Kxk8T52rsWJMH
kFCwAhtOinbu+TSDbr5LVrK07QYyezHK30ojk3MgaoPE7I3pKLfOuvTGF01sVfHh418RuV0wpOtK
zE/6wDiglAfc+rY7kLDWZRs8qhDuhJyz6Rn9A8XqzqWi0s8wI8rmvL2+mnKDvfBLCLdje2GaDTmC
lMT8sh89KRMwWUKgmfObrFgVHU8J4hajub3pRLvyq4lOgZfzrgMSsrf2JhxpVyHk3qnsyDtL9H2n
74cwKbOoMtQbdbJfqUIjZxTFRAlS0GIEj7VhjpROWlhkEBATXc1YEDBE2tlzsDTxF1JQG6WFtvL8
jaKP6v0kgYeKKX0xXFYp/7vZTK26Xp484x8nghB2NZPsLmbgbFFs8Tk2r2X//QGJ8kwBUnVbu8uq
vGRqx7Uyi7zeZqpjYaLGW6WMRD6Ere0Sgftk22kS87pgFZpd2olaaeNOxGW/KkWtqhiRf35Xx4IT
JiZKvvKfE6wLJRxvamTlbT1ObLvR2qxeo0ClziOujatT0kn0RlOUPZGQqnFdMvbBk6+sifST0ZJ8
evqfsZHvG9kS3f+kqjmxPbAbpanzF2QIg8ICSNpE5qQYrG5qi7+vFdQStCHvQdisZW8qJKZ1vWEx
vfUqisiYvYmJrK0r46pukLWKyjCjRD1W5bHy7649la5tZgf8V+s1EHpplDOemK0Uw9Cp1GKMsyqo
lPyNA/FoDROqQd40uPE+o99QjN9wHHUmDYM1rL+QyYSTXtQe6NGhTC94MaeBgFUz/lUqN2Kq8oYy
ZyeQJvQ0qYnhwqn9bQ4p5+4NeD9hlxqG1osxuvwW5exeB9UNoZwfEabmM/bpbSK19ywPWgcNCkO0
FlHrxWAMNhltm/eZG62NSgQd9Yk6vvLeuBkvCkaQGAimKrfuyG1frGY6z9MBSxxLoeFnBXAhvz5+
HhFPM0vNU1AVk2DWT7mNkrE1UJlqMEKxHbiGBv+PcFU2vHO3yiLFZq+OdwkRr069T5tWwAC/LFZq
HX/fz8KOLA7ORSuaO6yHoplx+Ng2cp7BISS1lP7nm34NocbBQ2/5Dvi7cRIz4s5iTJX45hwoqVH4
RkFuivcYM9fDZMwlbB83NatMKYSTIIHmNlSaUxQgMISbI6U1+ZE/hX30eKPVrdbohS8rT1uAXVVM
8X9Ab8EiVZszfyIlShmSGH4EjuDdsA6WlgEA6oZWmUMS6kXMZnvTsmRVXSvph5l4aSDN96qoZUHH
qpYUjPOVZgoFfyEspcX/bX8PGK418u2nVX9AKk21rbLSQrWg22loRlVM84uMkWTurb9EAgqxEPnx
QNAigam33b3BhzIco2wFOPfb2K2vuAElOGNnyhkwazfhiD1cq6phldkZdStppVk/Obn/YbG+8zJw
hVY/D10VmtreR9Sat7szm40ICICkJDPoL0T2LO9kssXKs95Guvqs6PmGBD1eHbp6WnJHLc2OZzom
JVK0z6csd6ZX0uNsddM62oFgkisn3Hz+BajEE4Sztn4t06aCM5nXjYyh4Yfw0emRvYYi2mlNrgms
hy1ekO7wRHjWaFfPo/4lNTiSMzGhagZuvC369xxccohzOoOAxrBvced87W7UG5PbitNpKgOkkx5J
v1BciZUmkX4A9it7diGSBRrPjAfqrPLKOw+KlnkHGnldxFHem3Tht+seZlt9DIO6eZncVrMx7nUk
6/O3nE7kO+WCc4v88so2+uT97ymnGHfMXKOhJ2n1Ol57Sohrpz1KMxqk/OSSNB5azGBnp1eLtxW0
8FlJiFdSLkfdlGLItB7hcS9zOAcewcTAWVlEM6u/68f1Ipw1WyGoOVMighP0Ur0zEEbGetaRrG9k
t6v8O6H1n7na1qv2dHPH9FUnV/VuKGZwEXrmo8uVuSPMLDcYPqgQYEhnSjfn7yaCJ0rPuD3sQtan
3rl/1h3HdWb7+stmvF0GFi4iUE8596S41I9lfpFaMg/40/ARKT23ypApsn85OB0qSln5bffkCW8m
GOTywooYzSStOZj8Zdllti4apjCQq3DArzsOT7DqhUf4oQfhnwP/1Kd15zUjfOb6J1c17tCeVNJn
wSofDHYDi5vGzH9UiVSrJO75pmoi4vUNRr6TM2G/iRcCtoe7MFIwgbMvajqOD9DaCyMplyZ04pAz
RIPjOLjHyhlnOtdljjQ4BfaXWO+HNuVCnxjLCJwIszm4UGZJVpZs5I01h0qse2fnz80XxppwFeBR
yPN3HdycIe0BYLYTYgDiJ2mTRUBuHcEEJXJkV0TEy6ECi75QqzfDxlpeenTHQfkGWtqZbApVL7uj
5uCvNCmToarXSWkW6iNmdE206tSkUdpu83sM28Mclgm3eHXXSlY6R9vTT9GfS7ZWJ9BqZucbx/hK
SkM6C8EstiwTz/dERy3rQCrHUodKYfIGONrIwVLqn78M1JDTzljWkFllY0abr0zNAlXHC9/1KbLF
OR2EVxnYLmz6Z9gtesAT+51/VMR5hTZrVud1+rvUwdWHvdMmd8/CEMf2A+zV10NEuuON3BvwxN27
Z26HmJjMYQMW5uLB2Imc0zi9qZbDPp6invU87FwTokzn6ndrQt0xJld/5fUpAsaQo6CCVqnnnfHD
Rg6D8NZ1jsXBAR109LUWDWSnkhilM5BLirQZlQ2GaPb/Bz6taZ/5+Tu1imobaozl6ff3+a6g5GH4
6GeSYkBaRYTzCOiaMfK5MljqMyde6jzRsESoG6bw2JMAGnS2Kjzzs2em6UEpZAIycg0xZXRz8Yd/
1lc7ai45r4IYi60+LlRm894CGa/Eu4sFGZzQgJb056arvUMEMNAnGnE/3j/0dtysI36aan1+64+k
ja+af4mRsyHrDYFCjcAPDVH9wg86CysiSRR4eHIDFovpv+0AG7lNeao3Tk5gmHUhHBumAdg87Usx
BENIAijJjdt2OfMVF2o9oNiD6gTvx5b1IAUz0GffdZH5/FjBIw8oRquJqa0BXiC4dulUU3jGD243
Ptmx8OPuT3oChJQOrBJBEa+Z1Ul6wuxq4moRoKUAdUlTHcjVyGM0H72LhytMZD6yEeeDA3lFJ92D
3G92QDaBDgd8+rMxYhR+Xj0xhE+RQVopdBdq3cbOtfz8Eb9awhsXmEJJBkQUkPllq8YL8Q2mfBXl
AL8QxzBW0fr+N8Vhmwy2HYwBmamP8Pza9ZeI5f8wULd/fK8vxJDrBSBm+Hke0Tp3aBhkRGFvN0uH
CQ6U6EW3FRlunATi2Nex8wbLI22iLUaXtVUawsGsVl0PecKuFl+dKOY1tesIsQTsZoqLen7FsQJt
1nXmVg+M6OyuiRwGj01wmoqArfBgOb5ACvg88Fl7nRcRpARfYehaaYOzofFpyC+P2HrTXCgroln9
Mj2np2azmdteaDFsb9rLh83v4IrRILvIsizHQAHcvX7qZOdmOHp/fcDIw02kRz7gllwWBrEizsaH
2yAiJoszjNupPnv1Fc94eqwWrTCyl/a8RbWCo4ruvvso5X9lJUDLX+BWnWtU5WFWjYn+OGsBjnYS
Kaeto4Pl/lYCjDW55iKes/6zJmEJHZJiNGTBz3QcXwYUhRePHSRorG+ZAIoQOz6Wd6l4TrCXD/B4
wBiVTCCfq6CO0eCLZzFGfDi6yrnygPwHXnX/vqJ8D2u7+cy23moJ6Rm9z1lyY5N+HTgo5vp7JTru
l4JM/HmRpeHqpL4ITX7w97oQpts7gfuBYM4nMYtNDXduOxAba6isHFsEB2xKKJNnIG38vVynHiFy
A5+6CGmznN1nkf6yoma2uJVah5HwXMmIAGR8U/34U/UEtJEYrknp3LjJxqFwolJdW0AsysahJfkf
JGnbiu/aR9HXZM6GhBKBZltZSFB5wh1nb3FbBhXrhBcQMqNG7UIcf+1tL1nzGr6p4SPvYStqUQDm
wUYfmvYbJUGjA17T1rWP5VyctSx1Cx3bh6BDL3nTCJh0x9oVQOnmqyL+8XVzjqDZTxU+USGOB8Pi
Tb1W7ZY76ZxjiS/g9olo4DFZt5wsXMh/D7B8iokiU9JN3/UpxkOkLoDlyLgcYHwNLcUMv3R7mPEx
PaQeFhhF76Zrg3zxm75DGiOEDH2FOZ9dHBFqmfjbQHRVVDtHZbvyfCaoYHAtFDJTy2unqd3Tf6Cp
BfI1CUbTwxuHeL94KPQMp4G7UMann2ZsBTzxW1s7m4zXRAlHxmnPyXvVUew79WdgaORjkJGpqAdb
fchrgp2qWbOY3XMzdKKhZhmNxKxQK+yGIthxFwqXiwDB4ycSwrU/OKwaq0D0aJ2jIOvrh3PhDmmV
jn+Yn2XNl7Q4SQGO/86rhZLEAyorIv3mpP2jlIcfBl6qH1AoReUdYEtKK42O+Pvj/tFjd1CXRldf
lx9mHLfv/8/0joEx9t1eSP5H0t3CIvDPJBxacwPsSrqLFVWLI+4BxD/la51Lj0+LILUo5ucfSw5f
9xRjy9vjLiMUOLLw0GZqgMQgieJ4T8GMCpF6aPX6xVJEaynkbDZfGc7NncqMQiRtOnnO6XLTz39L
NQPckJnbEhtS9aidIXJ8ODD5Bm1IsVU+IEHVf6fdlxo19b75z6wQn2Jg5bBvRfBAbEzuT0EGHL3D
CAb8JNC6PM5CedBYQl2uO3REtCCodTSYVWnAZlNGE9wlIb5Th1Itl5yd9XUwhpvJ9VXH/FFYJuEo
wQfLpG8Lq2OGnz1ZWBThgFM99TseIjLjGDD/CejdPWP8ihGF53/JXm2VGKBinR5nrgduI1dK1feC
5HwQMEV3Xrym1U2Qr46dXJzSBQv5Fi7lLbXlDa5IHNoIWOqXb2UShS5ji6VTraxDENImwEm/hm2S
i/py/3L+JR33T7sepISegZiEyLrz/V5SzLlnEWORihmCFqXD9ZYHUgcQAY0hW/opT9U26efjO6A8
I+eMq8pGCZw0UvuHOWzTbIuKKVyZX3CFL/t7aQzoGWjBMRsDX9RoOYoLS7RDWVePKlFI0rwWuwIl
sMEliRi+KCimbanUphtAOa2RAAa24+z144pOeRcm6f1Of9uOwrhzxyzIbDy+JoXvhWDK69K99h1Y
h8ALdeO6+xeJ6NE1a0rhWNUGGTaxGNJW5gKUC9LQXQ7tUlrE3ocq6nbWzDWdFnT3Zdttn5O5jgBP
2zLDrfidpj1UPU9xyBAXGIpPykJrr6PhnnPE308cl84WuYVAqcalIg+Ly42V910Z1kcQMfSbsfnf
+OCwfU8PnrpUbqNRuVbIdgyocn9Ix0USasM2yuxB/pDhYfZLWCXhWXgxC4XonxaT0BfeLpSgaq38
v7qpiwSroaAtsMRnDYYZ4HfQ2oSwmxfWN+6jqS0F4JaNZhpiy2iPT7bcJuXZNw6Xb0bPOUoEyg9d
rl6jspbK5BQsPdgHuBAbCWbzwKvP9e0iyGdp8LvBsCMZDuBTMZFShcz4s3OqSePGumYtgQpWk4VV
Y1vARZLUMSV454phCnG32+vufCHTwQg2WdQIMOoEgubmGHdiPDDXxKxbhXRIm7Rpdf/11rqxNZzi
UJfk901gsm+Oq8qKXpluxO0Jx5NgexE8ffTc5dhhu7F5sEJNSixs1I3oDLAE4YDDvSVOsNnGkJcY
VLFKbGNWSv407eIw48homD9mRamL2ruiqlGbpGYhAjpmwnnLDwFjrnDXEh4pme7FhgVbIEWEqXPH
/TyqN6Yx4evW49ILO5wJrPofU+f5XbcIVjMb5FV5yB+Yw6EgQ7TWAuzj1B+45EXWSiMZykDqki2d
HxUW+uxztFNVGU2hr4VPmhspkEcCXhzU9yshu5cGvvFACjLedqdBGW9KwGJv0PHD7z9TWQhU0Dkh
rGapxUH1LABgVIn9WeL7JalXHqBLKRhvg1s0y85vR/lMvh10xuAs5khlP+XCU6mKSBQHIQi/oVW2
FtrV8SQgsk09CIL0zpWxQZruT3QV7i4zNOg847sjiUPL7kvnh2aXRinrIf4E/bSu4JVuhbJzXCcT
rXrhGZHCMhAP0Ymg6H0rfMTEWKl6vRi7sJCE7YK6KEUbzmf7mJB9+HnXyNhFzwjAV3toMrDmgig/
YVFcnNIaCgE89pjUr424R1WbyFUIG3Omb40m4S8PSfYdImVd8+9tfB/dJ0Pp90o6wlh3fyRz/Ss3
xQlbvQDLn9Y0ebW/MjpnBmsTy2kea8WF6XUYJiM5EsMCYdfm5h4t3nlbBHeErJNth+pQPIbumfZb
EtVcu0qYNFYvwXVdijewkfxO4wQ+ueuo1LRt8JqgumvlNE+WVqsKUFAMdxgcCtF86fObpNK0VLgC
IFFGz69z4soSIV7fKXKpYu8RRBlYQSgvieaJNz1dDHLI8o1R2BKGy0TmDvghlq4HbC45MYvzhI/k
yM0dXLig381N6a78sIGAW5eJhQjeyDhNYaWgOtRJG6BsR7d/dassT1QPlrH+lZTVg+IwIPU5NHzS
WblNWg8BaAMTRYftLwK6h7wM3rvHo6l1leGxrPXV1m1iNkixbxudTH6ItKxT7IUTP+rTwVLo42YM
CG5nxTtqg6asCKdC0MFyZRImT7bvvbqsyfWSr1msoIK3lonIp2jWFc+uKbwxbuxlxofZ8b0lz+tI
k5d5V1BaCsSUyZzK9m/1jDe7w0VRE5v6mx+RYt8M/TH+e5sv7nWS+8kxO8THh4Lo/FCkpr50Ju1l
kqQCDd3ZHEYXeCcXO+A9GAvBjJ4HkFgLQ0sh9GNcmQHSGWfYyS5v/X8+9b3HOKfSaR9ZypaT/g4k
jI94FvGWhXIRCkvAvDPLWykWJV9OaesiSajSwYrPvkq3qF5JFQg/xY/XS46vyElK4hV6vxVzXQ+S
0PHzaRAsKNDOMFpj1rosmhJb9r5e7B4LIBIf7KevdR+7TWN5XDmoauIZJqZjEzdf93SSeJNHnruG
rebbZCGVGRPGck3PXmxbc2gOxBlsim3CYuZv87ILG3S7TitMrhtn9SC7R9MySAmJBqhoHHTzQ/Ti
UC27hWIUt2EtkQ4th74wwfBpTecXIR6v+WcpZrCYefh58rCR84n7ReE8QkuNFixKX3GpZHbyRjN6
MTUfG55F11+ATGVG9gY+OcdLcW0wInomDQGLdccRkMmPqAcFvLr8rBPap9HMXga1Cp4359LBiLEd
Zs4ZTSvODA+ZR10840d3Uqni/1NXdcmSGRIqdZzQvRUasiqmboMQ4Lx+dj/2HuPArb1U+v18ZIe9
V+TAt7ppq0Mo/uWfhDFU1ixOT27fnwBbhoLhB6z+I+ima+PEB6/Y3dHoEvVygTkqix+pg1Towjh3
1YRkTc3qJCL7Dph99plC29+9OtcEd4AEbvWrIJCPabNjxlukX3uhGrY1CNj2EpQD75u85TNwmPOj
v/LoCTcBl+PIgunJkmq8cjInScucTnVF5YSDPMrApFxhHYaJDpz9vJkski8pgsUT5EWc/8ovS2Fw
GHelJvl8dszaLk9X2b9iq65pViGwu0Tgxpl1JbUnjzHLhhjfkHiufQX7fqznMi5LR0IPiIVw88+a
RuePjPl5jb3B2S8fJ/Bw1Hb4hA3x8Q3W0n3+Y5ELS1bv3jxU0zq2T7MhhSmYiRL/9tFrxx/+lA7/
CUpUC70ehqNEY9SlHijXgP9cSLU5zaTGWOI2oPQmlDkKlMmSVX9hiRBByvtWZqLy7cJEebkYFA37
spsiyxWolIIrUQJIwd+7VWAO2L/whLukoTttEzQm9CRUvQrIC+sf2Q8Mibk19mSa03ZHKo/PaSJA
RxSkfr3GIXxEVjw1zzNU5gArutfrb8yazcqxght5e9nsMamf/DtRiY9HuWMjGHeV4HJmPuqxS4U9
Mdlw3jV/3nFAuHK9rshGFJYh29tclZwmw3GVKS++HpRvFqiiw7MqwQjl7tJSBwMl/bLGM/Qj9KiO
Ia96IRWxvmbUJ6a2/kA2v3vtxy4mMvE+JBnEHcL7XaMZ9EIcNO3t5RF7sIzqjgzCnexxCevD00M3
Odw4NfPCpLx3Lpwiglc5QncOsB7Wvx2c3ZDejpclZII5/EU2c8+t8+Wr4X5+AzbL+AiLiQiiEoXZ
cCH4k1729BVrYx463l+B3x0IrfntFyI04eCuIBHKjgKxxocAUQylBim/F2KM6hdSNxwWbFClbhyB
m+GcVFssJaPqbNOB1Y2nga68p391GOV1cTozSMjlT1k7SExQ4AWkQuub4Gt7i/vTV4Xz/FrEOWM2
b1yH/2sgJRv7RmDiY8RPkVoMwG52c6M+JsuW11z5AMAm/NlGmTNPBs4O/ELgVvE3Pzs3vz8YZ5Hw
b8DEGVS1diYwzml7dSA1XJLtdGx7XJqJc7oTM8sVqa7IpcGZjNTqHb5NKdqQ20sgXdUFzT8CBBq5
ewOEwJnVWBO+IVnMKjaG203Glji/6pXOsQFHmegB4t1w3TzBOmBy8Xcu68p+kthmxJLbJ/bVZLss
lhLYmqLMX3uTsi/jE3kFzFl3nFaj9252BwBlpaYyK4s/X3wDP7d3sJuxclfvzgcltzdR7/PBCC8L
krz1uoxHdSNur8tnpwpEKP3aXpM+GzAzsjBSGnuC9FS/cK7SCmrRkKNRVPv7QATS1SsA/K2N8HOL
pER4tLvnwM/+NUDOgBa+afmQmlEVSmI3aRZZYDyYwmT3I07FpvStxnOmOusWBOx/4gwQrSP448td
xHD4Nzqu97Jl7XzHYdYID/rJOZp+hmr/atsGf0OC/tStdxzxjyVH08lrpiAHwYEtzadHdqV0qZ6r
IitQMKnsF84eXzk0RGBBNoVpO1JDAf8kyOIuhYQRkVVw0EibOGPeonvntQ19eMPuWbJH/+d/o9NA
wv/A0O5Pf+T87Gwdgr+UXSKyGshJx7tryi0QbcYKPtKFPsEbBTGSz2aS+IZcvZw2BJ3LgaMkuEYC
NGdkj22wHxmYL9b3HQhv0odnvWkQ0nIWAkE1DpOZdAAbSs5j6xYZTUQo92e5R8eHZsgZpsN1ptd0
lBMO1Nk2lBm3/sitsS0Ad5/q9WBbYHdknijZuHQs8TqFmZJurUL8UD+MWS2fNghciXBXL8mwxE9H
LkKLg5OB/HXD7JVJcbbnXwZ8RRWmhbCWey+OVbkbpxuOJH/jmxXJDlGor9DEdqJc3CWpMBqza0u5
Z9a9ChUszQtZY9LCViHsm3wu7xkJhi937N7mMrGXuWs47z5vG2bIovdiGHx2niE05aWhUcfGYqLn
Py/TPTnxGxvmsHeEEt894TNVHb6kDh3k7nAOVWYBPkhBNQ+zyX8t9TLK7nEJoiQHhpYGXLQ58yTt
1dzGY+QW5kDmpWuKJHWB1+rSpSXoy9B6JXO/6RHvFl1DghdoD//b6cUJRldG4rNMnWqEHQiWiZK0
ifA9BJob32TGs1eBV9NN0MQgw1doR9LkwTURQ06FK6PH2OVVuKpzxU0dr+uXu2O0JhmLeJ2M5KRO
31Aj71BiFNvjkO8MMTeRHj76gYZfzWV7Bo3hdNgFIl9bNMcNdmXfUpPB7XS88KUSveR5ibJ8vdgZ
xyc5Zq1SruDf5zyG1HT4D1tdGWoU96r/WocZ0lJBWlW91H165CPsZBmlOxM4HFbop4k1H5J9U32C
jP1P8Q4Z1BHx5uz4Ol13ru2vbmLR7CpFZRGFC5coGCmVpvC+FPziFZCkHItxKzgbiB8VJxZF4/jE
ujD+3k+I8MhGYBRUOhS5Yimfec2d7KCL6jAphjPttKhxhbIQIEG8oclg3I+kf7+rXFfRKqO0Phq6
2VREIIjDm20aWRzlM1o3SEs/Ha30Z7BoGMOLkMx3bMHqjUGcPxgPLKxWHpddBOdWCS7CohyOQ722
viiyUDcjsgZm2KuMUNtqnns8787wBaTKqJC6hiGvJ2gTi7Go4iUWeTDa8r+74hhZiFlVPkp4hpdn
JrZNVLW+/zVT1tsAKsNb6rbi6GPRCWx+rrP0dx2RhxbVxlob/cEbnjf397/+KYCw4sCoUMdm8uU0
WqEWNpJ567tKqoCWNtNlYsLSNAid+ODngjO8yKKYhodOTx1ObSW4W+s1bhHh9UlYxuHAVZHuDJum
Z0lZI4LCCObeKfhq2T5dFZWsgshKzq4oeAaaeurPPT+EuhFl7WL4CjLdDvpGreL5hxBtjICEbtll
WXb1ytPWDAoB4rNtYFSrB0GcjOc7czYHtxBHysdKT7zloxZvM1Yaa0nf/XD6IvrOgIcM/b499VA9
VCtwKM7jTVjJs3h04nTg68PYPmIGRqEbIxmjnJTlszRWzUZmtKqg0QyVv5yaq50k94MTmq2BDXkb
D8rbk5evn70krbqUwJsrfro/cln0gKwGJAo1KMLLLKaGEY10PtIYD7Rwy4xq3Sj7BiqXD1CNy0qR
5JpDZOCURqz2/AMC5KySwQgXFH4otdiub2RUAgTQ1SIZ74qFpoq8/JbQYukewyNPodTJXz/rgLDD
hz23RMvcw8BJ7fZJ68gQ/NCxGEeNEvqFWZgEit41e/WcKctbULaAx1+kDwsLSV4bvRUPAOTHN6NM
k8r0M8BUexOWGBe1anZBmGUUd+PnmsYR6R7IDWUBxYQxb+/+GKQcz+vXFcUqLkOwJIYYDx8yca9F
b1Y9h9vbI++9awzyjLwxgdnMBovpYTMkHIn1j1MZNIo4haL5tSGJdalD69zWJlO9voJIykgwiwdr
Tad/Hfpbc62QpTK5RqbXRmblmFdWHO8XS5oHksHA5X8QudF37MFQ65oTBo1+rhwPBCwAHUp4MXtz
65zuGHcnagXlbFX95X1JC5r/T5WHHGSw2O3cu9XQzeY9NResJG2GQmohju+yC0ivJliyN97wUY3j
rf/bWVTRwSsmK5w1N9kK4QV/RPhRmAbl/RRLwfeiDB2wXGHp2u0vmITEIG3ffu0WePYMxtATGdIa
Ef6RJ1v8vcZC0lWPRwlYM6HI3pSCyMkc4LAK0bm7k3eIK97Paixa9BAQbR6Fnhaz2MPEvTLRwxO0
Dcw2KFx3tUgvJ4xdMPf94u+e+dNRvEnT2Kp6EvLWn9HC3v+BP1Vwu+6a3W2AFY83gPuk2DmjFDAY
SzLq0GMWZStbFHPGKBR4+CLRfgHc5a2nzZkCl0OGePsP58cCFJX3eDwSTWr+Uuruhhq2QYHYlFC7
5G474BTIOZj/8WLfswEhSBWFDc4nngsI5xomwPQqNJu9xVgOBmCnm5eDt58MSIeagLoYj9obRcuo
SMKx97cv14hfGNUBtLWzkTWqAuVSXVgOyR4IlasjMjN4s4f+cUHYw2oSAr0dPCuNlhZhdNzqSH8f
pGPUYoES32uxyi7vgE0UqxGOUUYn3V4NN0LWsB1a62EdWmoIVnxuKeRiu4sVl+Rd2macq5l9+4ES
0d2v9q1gK7nMTB80W2VrrpgSpEdI26Kwl1eK2roUutFBNLtYXAMBM7l+DWCWKV7tTecuWH3xR77N
1XWCE31hTtbwMAqWZFXwouDxaFnE/hemsH6vKXXf+w5/J1b8FUbZwBe4RyJwWAaz5oFMVqT5TNYk
olzQVdV9N3Jt6v0p1B5prbXc30/tQzVYqx1OMk35iztzUJK1Rj5qzW46AWFCyjOVjfPG0yer9G2c
h19U4PqHPJfq7RceDUyXifxgXcLz7Uic9cN/x/1is2FUpnO1iZLEO1FfHevq3Ti1kWfg68U1wSdx
0us+7jZodXeABAYSaHLC0BlTbqGKe++38zPaKG7ugIEvWVqX4oG/snMuKpzYu8d7aRMKiEuYE/Ho
a4FyzJia5A46CKYpC/qvuzCSj04aJgDJzgtqP+z48bv2JSXanUrqGYvrCIsXPH7YVvrpgdpuajFC
HVZrtSMBtdbGTIV7+a8jCk+d4ZX+J/cmjYjAFahLU8k44e7RuYkScGh5xsDQ9AEszxLfF/ejRaSH
O8hs7cPQCKSQqWnOFe7HM7/qpW52oZaVWMFtx/eyHDcYQ4nfcw36MhdQFfU8OkyfvQ/8XmpZkrmc
X/l9fY0TLXRNtWgtHUw3Y+BppskjNH8ny/GYlQn8g3xOk++tdTkUuxU17NAppczc7aw7CarznL4C
Du0nzPWA9i/EtwTUBl1jre3feAT2ug11kmPaRmFEnlbrFzcuURV69jemPt3vi8uS81GXUhCEoDCf
/uKb9zj+Gz+G5bY34EY9BmI1zashvORv6VJYdbJRsEGkAoTxzbjxOe6bz8CLE3L8p48L0hloJfD9
RZ4otTsBgkDMZtlGtARZZhcfqm62LOfXwAyp0xVwc0zRBiIY2fJhTVYlafR3wI97f5kwUflrReOX
IWJKMANzi0oQfhgHxCUQ3PSQpm9ADXuv+3L5Oeq9rKo6eqSWvRQCCurb+/t4QWVHr9YRzqRL9Wr6
7BTL1E1rOUFpvyVNPPrGwJ7xGQY447mr8BWf3kuhPZfNusOybCyT4KcX31OzukUNeyi3HBS8f0rV
KA7Vy+vwDRK0rmE50S7sSL6fLTI9v7O0CmF+PDpPbJPAThKJLPOaKLY2tJCVhqxUkAI3roCSJal2
sseqF/yhNXodDa73Daq3xGFrokxwSB5V7O5Hp5rMpKmzNBd6RDugc16aHcA4lZqFBrpLt9RzT3Q5
BJ13ky+njeu6JdHG6pSTMysRUr+PMKHLdP3zwx2rKf7NB5EKAJi0TlZzSyz9j7BLxsTTosJSSs34
sIf6MSw6MrNiPz1Og3paWULUsvU/zoUVXSfjRw5/FOEPpFAuw1LVtQz6w4lYFK3rUK1sTofTGKBB
tGS3N/vnNhGMyyF8RiAMdVHM2fl8vfap/iLlIMq+Oi07QZ20J3QPG5atIA4VmmeOn+XdprXxm11/
nq3FqZ5oBvv0qKYnlNxnX09oz1VuG0qPsPP/nz2qcYxZIv5cxNuNll+Nh40pxiDQXA6rsHdMytae
gQAzCBjd1X0r1wakGgNbvriyhT22u5NmpkeemyykLC+1qmYLKkQxPCvUy5gy9lI08LYz/mNT/G4J
4XSEvM2kZfkoFFhKT07ScSGeetthk36gONsM0ZZstoI7F+kqEj1tVqIR/a72MRCqenG1Gs/rq69H
aFYb/ptPxSSSDIkhx3xOe0RFOWM+rShrPb7e2Rj9C6VTcuBGHhaSGOBQpJmXRpAxeDPgb6vJor71
unSLIN04U16GLlO8tkwD0Xa64HO3YxwD7aCpiv2GAgIVZON3MqjoH8HI5O1ayJXc5kUJVB9rq0Tf
5a5bKfPripf48gI3adRBTdNn/9J7U1wZJ9KCvBB4wMtZ5n9mwa/M21rtcYzecFoZ2WUf0lHT6cbV
5j4XIPprz9KkRH1DsU7cnmdw83LqaeSUK8quzdrN9Xf/4dtIZcvap8KWrsXZ2/v86L126ZxIUvDZ
Y1RTf5og3P6Uk6S3tuaKrbNdYlc1gP9+U0+Xn/TtgTg5ZxS0kLMWRWWHs4/R2UiDTXvHjq672pfi
ug09HwPoNOp1ZEduY/cbAsxWOV7EygShwRJTFyIYjTHEmQkfgjPMWnGT8Z4B3hDHJN1IL6/LGgz4
fRZlCRH+W2Nrimzf3eEl8klwlO/s4CiJrVlyfS91L6BgFERlsfv1tfZ0lpdsmyKdIPzWOQOGpTUE
GJQk306/Ag3anZF2IqGUZVOD/QRUonkj9U5rpnE0LVtjd3CUJ/Slt5c+rejcgKy7G1JIqXfKCGVw
AHh+rP7rGTuNB9PdB8nmfeR5dXlYVoWJWSmpF9JAbsEpt2nqUK14OIFqgGAUIiVxxvurkJ+ZqR3p
ztNlv0nUaS0oTKmzObUQkvXbMnslQXWQf3ZhYZzca+lnQoIfaugjgp5Do7ZWgRA15xieWyr5wb9O
FMAabpPrxVCuKM5MNUvU6BvqYrJeutidwIMN2UpHSsTv2xPZpVMguqOWQ68e03SguwCFWOvaM7cR
jxtDW535o2ZDJE33Lrrp5bliiUDO0Nus1dPtXII6OBDwMip3VCFJxF3St0TDmJzR7myyjF7ryaoL
Ddq2WhvlKCiUXhSsb5uodbHBFfXpuoqXdEInz41W+bWkgkaUxAwPiev5LELu7QSGyR1RMXGV1pOF
wyEdpi7qbEgSSzVWLxF71zFO0rYDAw3GTo9ABKvowy/tknuEVwVqnf4XAZV5NvZCHYS532uT7WUy
X2IHf1rgPK7kffajWw5bpJMrff3bWdfrdSBFL7XK6cSXCzpVG6OytgEWibbKP6nR+qf89tvcpqu4
NzRUoK0OhTtWkYwO57vHAN9YGtUG8+paAOiWyYdjv4NghCtMMl/lIKKO5YmtVG03K77lEtiVTYHo
A+lNg+VhyL2r0Jpy3fFKlFgu3A37XNzZCS8okbDPN/FyJNAROdMYiZcFPUqvU6agG0VL1tBqWFpu
+aPa/9KNC/7g5E5U/GBdloaKUKmlZzDdbsC0mqXJRhOOgMIFcaY2jeG4qH35B/LvTDcYdbNqMgxk
+oLJDUC+KIsxwh5sidYEoZQiGApy6A02VluwnPn/Olb8CIT/Z2+yL/w05str4TcjpH88C74RxRY1
+QVyVWBJ41KOHQExDabirrmIG3g4OKQY5NKZeExt/ur7FB4UNIOvMRb/ZGyS8tB+vkxE2Ytkkz3V
claUWtBGHXX6d1/7iB5nUbFiiXql8WT9cJqW4DYwaLsBDi5YMAMZ1UA++CRHFgOp9GJCSBYaEvlX
or03ZfSvmfc71RKrpw463qbH4VtNni4rrxPWuwTQ+6eizzZB6J+w5wUnP8HhChKOqNg6wtIaGQ+A
WWec0gT4NHWj4EMJlfRt3m9/LVN3yXU8wNEcgAtOsR3sHArb3YGWyfwO3yJryQLQwGIdyo8vboZG
4etXCUAGlJp58cIR4HYk8+2cO8cNybe6pJhHTTDLUA2ttR1iFHUdwuwlAHhNXI36DTNQSw6TG7M2
FrNnUHY5I+UCiW8Kk+39bYfFDiFt2jAZ48B/JS0RTa/85L8ZYkbuoKPRVPIo9GAqlW8T7dXgyfRa
/KJH9OYASnXFUCB4t8kQh9TUz1YyuuqiTi9vUps2XoA426MtRt00kZ4K6+xNp89/45k+bvnY06z7
LgOEJTXWgTwzr6W9/t16T/jk7qYBo8qMBcC8atL/F/ES9zSHQ5LcP2vgTyTGE16sDQL/MrvRhPBQ
5wfM9lLSuOteoEm/P7wgCa1rmaUKcsXc53S+PWhGXRAH2yBvQDoOWaD9sichPeBJJGvvJwD95Lzz
NxtkjHV+LP2XoV03Gfp4TtpDl8GDn8AeLVntQm3AIu6ZQ4UzD+CST/aaAz26MCftX++NXQ6GHRRp
1TbX+s6+OejkOvlBg4MpQGdJoLub4axMGIGxncZ2b5JEjOM0cqJsveMpXRFPB1dlgD8jv6cYG9Q6
cIItVlffjEfqpH2j4n3jrtE8qQ3brMeTrSmJyio6H4UlQSJK5QKiTSzzEA8wJ2ViVsG5Dp0D157t
4c/RaVbmpX2IKAnYUIng41qLZm4xZsaOdnWYmozcOeUoshZEIf/k73DKATmbXEn48GePca9tZMJF
oQAFcan2fn8hYITLupD1bzL42LI3WPgUZ2ZdD3GJm2MR+H0m02+XoZNgNrcY8Tlwtdtj5MV35Rd9
r+7pqyxkROpWYhL7n1yP/mlumTZC7oWpNmVu3SoYgzcJGLNQXwCSiAsa+UBMpXvGUTLL6eBuOGyp
A+kwJx/MbiRPonJCqaOqZ7CRh0ub08vC7bWeQ8FjQdbWeozsZ6fJarHtof3bqtAXLv6inmhiHe9H
9aoRIGL0hjzfmCW7bVpeIDNP7zhiXm0gHJk7l3aTte1lZOGOvWTAChcHQEX+6T6rhJfcjVAaN4E8
zfDIeylP9xRwa4RA+99h9Oe+2A00P8eIaelnIFBbikLizE7IoOB87P7mbrhjOWKQ0LViVB1qB/wN
5XaIjvdPSUJsN6I4LMBCDVhsBHojoLn4NDCnfy3TBmnEUItDKx9NBkaZWlHESIkQfQvCE8s0wY+5
RXjrmsz7Ns0Cpan6ym6GPwOaY91wGkT4Kp8K/axfdy8RwAJX4FWiUK4iULdwCnMFoBlPPYUXT/tA
r/zu4CGnLLARSjiqVBaRw4G/CIwVxeVeFR9JVUZI6kd3MzAEvt6E70t59lNXNHcz/YU8OflrU4ai
nt09WBrq1RD7Km67dcWdyGvRanxGQ40TwbLjOK1QxmGDhKt+rVxILlRAR0ZlIka7EUxWgV9pazdB
pA7RSAdo39Y08jM8l7y8EWu1FAZqReppHvVZsefY9xb7RduyMoTAs9NbG293dlzmhtdNIMBlY16o
TgTiGlZCC4llDya7APn5Ph3JgggpellyqrbDfbLuj9XgFIH7niHdKGv2eCGAmabtUcjiSjqSyqQu
Q42FezF8+aJQ3LOML+N1v1mC/elHdZaTLY4Z1q2gkuNX/yj+r7PRoZ+xaVrkhkdkN2sw1CTXC+WK
J9aLD29dPV/mMseL6q42NJ0tizR5AQjYSRupO5xcE91lO74nqilebwcUvgeGQtcTlN1BFNw0UYGW
deskkghdxZjuF+lGdTahboXklKXixPbrGG7lgTmy/YXXXDyRZHRCW1nrkBbHRvKINd7Ef3GffoCT
ODwpVwjiNabgI7+Zq3CFcUBWcI6px69tNN/hY59B0fvMMc1PKAF7CUxIEU6ZpnLkRu5jmR6vS2JE
iYSWa3Z17xus+Znm/BOVIOr+nNEa+XO6YHC8EksqGXA+3DdAi49KW55dcFX5vw1MXPW1mxq48Cuz
V3EJj2FtgTtXjTlbmj60RraaVPCMMLzPO0AptjbDbFHPdfsYHJDdO8XU76m1HQRaIckfw9ViauiQ
xI6UxkD1rz8C0/zt9L4c+nqknbbvA5MlAW4s52u8zHaw4QiUS7PExQOGoaCRARb/Z811e6YbIKTz
0JqhjVJLqccwHc5E5zC61wfqOK1nC63iIHh2oi5rk7HBaOwqDhGRIbEoHfFkM3sLqy2Ncw+F/XJJ
1aknWxg/VDb/xyj/LXfq+e8ErRikx4iZdlEwgiXxkGsYk78dnTypvBlndzoOYLOqFnpD0EwjNBBA
IGHatlHOVRyoxPfs4Q2x0gXs65Z0RHg6Tzl/LNpi1mUIe9QpJRCTXDBKlCFWmXOL8+dbUn/eRWTp
noAxHLbPBo/nf1ctjoOTWzcU8jN2sS7S3YoRL2msa9UnXPNVSOBpJddOrkn/1/fuy0UuAfpn0crL
TLI/SKpMLCk/8Tmyas8w/i/3cZDd8+SYsYhCCosAVgRxVfd0WpDS4qCxjKY578IzzSMWLN2jazf/
n6+SbC33UVOobK4AksC2k5Ezu3/AscNfuyqZtdGX6pPJxSf2ROLyXvF9C4POjeXyu9JXku0egpbY
qmEAisKk8Jg54QCldDVNMII4PQjcSssooyg1D7EF2LGbgbnYqV1f3T1leEMcAMi8kA0xMtzCTIJs
BqQpTpq4tVqAo4K9+o9Swrn3iZ+3vt5LCb9H5CVyCl2IU2xKEIbnV336UX3S0PwKFkkCsofr4Ezo
trrBZioiMfOKyaAMugCqe+DYe18u9HTfHMHmthRYpHQIloBvYW8Q6BuMUV8/QK+nr1C46a0ABcCo
wr1CFrcpKQHKT1ci+/Nq0PQKLL64SXU8bbDtZg+Hh2LONCwqahfFN4IsgvuYnxJ3tBD9YxOk6K1Y
WnvR0YEPhibrNg32CHQ1bwAmCrKFQeWbU07DFyfFRUK9OIPlrowPJR+iugHLpqxbs9BZROGC5v3y
xFEOXtptrOO3WAqCiyFyV+Y8gNKjM15Op5kjqns3XWLOplYt8uBBpaHqkXb+4WWhjfHYlULcnON6
MgbZei/JCUO7Vu2W1alqnjK1dFjr4w1ODJKzbCLudR0vPCMbyQ/iQxb+Fm47xU/oG/ew6T6xarMi
Hr3VkuOM+0qj4upBdNgtqdQAAtjibCZt5xB9Io+PGxg8rfb8Y4zC7SC1fa5/JMp+bBs7nFF7oQBf
VWpVRedgbWZRVkythBZkCgXbLF1kpbjzPbXueu7GpQEYpJYAj+71KeUwK9YRKjzXWPTo1rb5JAEw
ZtOZQgJKX8zXosSKxlngV3OAkTY1mafYm06JTeYM2JORVLkKZfEP/iuPHNOSahhYkLe+Qm1aKiTJ
QRk0hDdgOw+5Fud7ABYhdMS8M/A0tfh3jkm3Q6/DX3B//1RpQClKMuzglhd6G0IC0rEqxkvsGST7
33WEtWYc88K2ivWzyIYLymb6rXmOxuedHMW8l0V9HKm5uqEeCE1ksKW8SUDP57TpDVpZzHTOyG34
x08DLVS9DMLXKgUEEU+IEP18EoKXJOkWcMc7Y/cvsd+esJIon5mpdUMmV/wFOVF6+04wo+67WqqN
MDXaod74OB5h5L9sTpLLjbmG3/h7sxvrwtIPr1boxGKeuFq8bfbZ/jRq/Bi8WQHuIWxaKkA21ZsA
EmhmhJluCLS7PzDhdxQiB26tIqXV48sR/LUbEVRLHiWF/QAcV+0ATX5jclbkyZrQGP7tPpLF8SF4
yifHjBkG9nVOs7DafL1gVMbTsHzZQw0FMVxGB8yvd9zta1vfrtuazxb9drtkFmm/P5Q8RCqPcUXx
iwK6pktaiL4zas/q2blJMsCtT9qrv0qL5C3qqrUtIhjBrEyyBAu30F7hnNz0bxbym6D3pO6lW0FB
/fexFy5cbBoaJMXpkt+C7s8t11ZXRAD5DjvTqCFz5awXhbyyUDI73XZSOi0S87SbtqvTq+7cXABn
Yp2bcOK6VZ7ZbJIDmdoJMgb2nBu0MyjJtlMT1WTsyO7Ag34qoLWD2A2g5FPpbz0moSms92G/y7mh
759Inh0ZwLKab9uZQXXKSzfB0Ir5kLvEZ3HnOJVNbUOGrtVpgcaNBGhg698pnpTajLZzjTI9XX7j
VKmN6u2X0hK8vPv5Mks7g8YQzc16uGuJUwgOEMwm8PIwZ22W9GvXXLzxiaePbpMQYpSoVb5ZmPWi
owWpaC0tWnaXCB65vT8oeD069GJF2KPn/kmwvB00nBhR4vQjoOhaWyOOR3rJLZ4jccFcIjHj54If
Z3gZvGXxlHZz6ljDygmU7R1xSj9lE4ipOTUUjVoFbBTwsfwvWuN/2Rj29FW2yu9/TIE10whTkfds
bkuJcZbD0j5oKaCfqjsPK9719EXp/9xXB9LHiDoZgxmycu8AXtuDKUZhnJZHzDoVB5UdosofW9bA
wRtzO17kM5Qsx9ZuhRdH/YL2yhNj6Z+d407nv+AxVJQn7tOATVLlTCLpUPRk0v/Bb4CevD1NywQw
GDWJD6CNzdcjT2udTMauLAeTBBUBcxdgVSUZdLTE67RZvHofEqOg+1mZ+RSa4n0lw+A0mczWKDCb
wEi2o7h5vg2m3Ja0PmxDk9i+5ITFf12d0ltYEkfrfAErJQ9w8p7GaobeVTc2hNZ4q9BHUblH67Ai
a6RlTLWcI7qPUQm4ReKpGDRXLrCzSJ+RlQULj0Hpd060QlmmpYTimEp6Vv2hA2bIZWdZELz5nhb2
UKhgTbPU5DhOLppK0CurgFZwoPOHmTbw7DhJgFGrDzNhlKNJd86S63aRahZVTozJfhnrSZngG74I
01yjHe+6L9SfkOXmcD/91LHjwjQRdUbNAkyrD5C0Eps5yIxsH4NLwIltJXkGRpSacNZC9+fB10Ic
fDqeSq9zJMmMnvgrt/U5m/p9RU7hmey/VyeWbci1FgNVtGlW/qZ5ogMxWy2w5sHFIV8gsal/GBjf
2M9ew5+OBPIUr4RreU4xrQRpNESQocfFL3h2/2r1Bp255uAaj9ppQTcfs+odEddLJCE3AeCTBpSz
c/EkE1p1R5eCzJolmLAdRFmJJ9mmow+FhqrVIvC+aQ1CsWmRzADncaiFrXu/dITpa9frLBC+OzxO
AF5E9kKFI3XKCLSmoU0ucBKyxZHPR2xZIHcgcTBiE56z5RNUtogwM3MIFiJGW7rQP5rF7cIVmu2W
Iu3GmNI/gSdakAVvO+064yTmsqblE+4W/MEkB0w4DhmWGCmFnCh9lROB/+lA8PajjlQf/qHdO8Go
GuCLIlxwyZe/9noRSeh2eiY3kcjFJnYoEf5DYceyDpfp2S2OylU5BfzDAHY+yoY+sNg5ijnvRbn7
WCYMio53N1ap/1tgsaXrSCCqq4UTNyW7Cc7Ts2Ba7t6/80CCGJWLUgLLUXrDBU802bymcpBM2x2q
H+NyhKmvZ+kv2n4VxFGi15LVpdHn5q1QpPvMq0AmKrHTLRxZOr4ev0f7UPfhIpm0fs9lNsGaCnZO
22b508lUK+stY4giVPv7ScalvW8YcJVM6HfNjwFrGn+ytMxjdLriIJkeNBAH+RFR+NniW1oATKVh
sr2Zu0lgl8Dkl/xB8/Cvm0bAO/KEKlK3uLB7wj2sdl41II16mm7w34yUNfU2xV5EMY07FmCJigz8
6fbx/qNq36oSUV8gXFJRnB2aHD5k3YQMqYF2PvSADGtmhSGE/DG92vUqq3cJVXPQ1QrCZ+1WJ9Ny
MoSweu1YjsK5fQy1WCWbTtVB8PZRbaTAEpO/No6cCIE63wxxFdLctjizklAICQ25kWYwRnxIjBdM
cTzo/Jk6p+gjJjyboFZLlV1/2W10RlVaWWu50+cbLDPSEWj+KhxUI3qmeZmgRBghJ9vq+UMmNyBV
MfMj/CQzzeuMMc0JgNyCeU8utYXzMdpHivRquw37jexLIsH7ZbwyinzTCHuVLWAK6ypKCvLEkqQT
8/G96w9260CK6HyFawr7gqDrHuoTZEX3jA2GqNb88fXuj6wuP+NkuE91ffNFrKI357aUbcG+gPXg
A/rpMuI4jkjwYtJxsYOxpYN8PsBgK5uT451U2hbC/t1TUA+a9kN8fm+yW8UawfshV/NjFsDpt/od
DzLFBA3mCLrU+NzV5omb6UHZBFsiXRyHT3bE9EaYYDvJQAKK1NDZHJem/kQmh678TD8NG9YsxMUh
Uavdk19DqG2ghGKfReW91CtysBuJdlapmwLaM+NJypCjDPXuKH1f/dN/qNhGy6vyMHNNvEtx0dso
MgmkbJ9E9FXY87uQzZK+er02j/SEYG/r5EWL14Bys0/aqvF9BWh5SVzEvrL2PCAQnzwpM3Pw1qWl
qHjCflW5wDPgAfEZV+NflTFM8lkIlz+sCCQq1OD7fYIXZQYfm+QKuqKffHq9ITd+WCqHXkgZYuCy
UHi7Kux0B11FJ0IHgoDBlYb3REXVAE/7Dl48QViMVZX64i1/AIArz4IjzUxzmem5w99HEA7BkV/r
YO0oU7zV2u9b3E7rOqzmhWx4Ig2NDK2aTsPIhj1sMaE2ytxISprPzmYIrCJeYgDwkZ7RrQMCbsdj
9GxMDrcCXmoVvevLuF0De3fZOiodd0ZCGr2DUitXKu4lHC2iFfp06AFA1clIj6zhQe5/tLKYMrfV
nto62KeBeS3zzHRazr3KCe68s5FDQoiQbOZgmJyI5ORd1Ab4vAc+cl2U3eCfDOIvyDVKHrdRQWmX
SDG6bChDJIYFPWMLcNvXD4qyJax6gNVFl0iBP2IrRwsSZ7NIRJfk6u+A3XcQ03rcBOSvHv4lb42m
Iav8EjFUfguK2mZXUlNV/vrrxvuqX/GL+QBsDXAduaTQi+HcbIqhzEKptMDt56b38v87NzP9CZBT
G4xRD4LUScXtnIIgwnp9AUt8N/8uHxkzlPzBZZQ/ULQm2AbjvmTo9OXB0ucPOygDjoYfwOXJOQ8n
0dh0Pj5KTCOQ9A5ERQfaBcIkhrc/yjsW/nOSsdxEcwrmIfY5hLXjyOI110NoHCKf4VNpGJVOr/7B
2GTY3BZsIPKi2udv1Ov5dTEmzJTur0+enTbepCc0u+8dJ6qimkdibkl1qOuBB8q6lsGV6HyK1nOJ
HqwKarY2CCo4JRyF3pmfZZTPgcwMBhNYTgOmLbUFKQY+PJnBbsDBOb06IkmgtV1aiw5XbxX791tw
6Yraeckvj8Qa8Ct+kAoOU+pFvTsONZ/NOsa1q1/c+WI5iqi4qisQaUxqcvKnfEPIS9xs1sw5vcU7
5x2x9w63A4CxDmHykz/hJ1U00/iiu8WYlXOrnVXs/jdINFrwtM26e2aVZR3bqqvreWf7EXtExw5+
lSfdvJ0tWCOykwL17ddGcWuWAm9RMr3rwOfIPmBAj6AscKrfBxco0h7nxQVuArOcVRepySFBvFvf
SNfARKO+i8cUF+i2ejcOFrO8i+5ABSB+FSsJ5VISVSuOer2o0nqZ2xzqweafInuEfEGt0SUe9pEY
gGdMR3QNmiLHwuavOkOxSl4t5R/G7kBnp8LDQuKotz5FxblbkvDZwMZZ+CTYLXVBs1/fblpdSqvs
Ma6UoMA6TCvK94h4Tdw+CCwydWPiZHPXjBsrVgc/65kWdYqasGB7HCYQtEBTXjOMWYpk5rTUmdsO
mLRpqHUop0B9jat8MBw8hqSFtuoK8WEh57KDRGZOLhXyXVXhmGOHUbuUcsQkm55uJXhpnIWabkx6
5326QSoztXC9KI1TM8a3YPoB0LfHNDW0gfqosU/pjeFTXJiPs9fl5GqMOxR0t7zqQxTIIKZSXsJ9
yp7/T9YTUqG2kyDJ3xGEhX/5dvwz/ELoAUGlyqMPg0jOnSzeNu4iaYeTMDoQndouUuzBJWj248JX
4elqpuZb1w6+yGWlZqyTpUdQy3NaJNmZ+ocOKPLntlRfpq6+ILJYSZQhc7Q7GnnwmnRN9jSsaydQ
JiL7DcdPs9TLzIURk/1Ov1z/dmEMNJ2npM3BByzJ98CE+Vwe5DU8/2KKQC3m4fOUJXGcS8hOwJFp
qOmArbwqpQz93tBjMFCSEWCNBvCh0CPAAfUoKUYI0SKmvuPWDpdAfFOjfiYkrV17R6dFwzmX/C47
idYo9930pCSSsNxYww6J5ZQAsVLdHt9iQyojkxm6WQYNGx8GvI3B5dVeh8DYD3ryFog6ddwhSlyt
Ka3ECumtlRNlJL5U4uihWKGHmO7xPRu2hMyoVrPTovJxSCVB6Q9Iphui8qfoTk+7penwx6QX5ynR
HgOkL47WQQQQWBQj/Ihx90z/fIML/P6tsKAoIL/yo/5/LNDlv9d8E9pfh8HTlemyqPiYsOuRLOsu
UcuYqOjGXq5wROTp2bgB1MMT6wXZhYiZDuaOyQqrkde4mIIB24kN5AcnJ20EWUoAnaSHAc9xaD9k
vBMLL9UMMNfzxdbqtAIOaWHRgTlK/Im8rtAYz1BpaEuenBtJd0i0hQuHIXwVDPz6d9K5sptC2bSK
OqDGFY4ZB1/A9o3+zrYe8A3T/FO7OnNYyaZjHciieb6+qsGjbGe10afEPgPdjpKeAC1cwiu0AegO
KUhMOeW3CTsY0+uSfnaTHbiGmlUOnnbfOEqMnzk+N6G90bSGRg2BQgq6WpANKjPBzTGDIMBag/J6
jNtmvBfQQ7IZ3xrmQMTNoKvbczOvzrzdT0FPpd9r8YkLsS5h32eFooxJTWlSRD5IpABeiyAn4zFn
2B9/wPwZZ51+5q73WoLKgUNblRU8U+PYSaF6g13P9X9EKZXAhPaeCvLfxO3ok/A3C2amkuUTrQfJ
qc2itmGSJRiw5d+hX/PVu/oJMQBPQ8ULSSIGflimo1wyIl2MS+zeMQNL+dsnrGkOejsCnOZTGTUI
LPLDYtDYVI4BqyS7ByX2/j2yr9+QCA7dFDH4SC90zP4D/8+zXZhhdJl5gi53867/85qY10C1oYNN
zWgsMHDjFIZtOhChLB6YIj/yjgitlT2x/QQ7d6JKsHBnkp5YZvMKMgIVMhUXiw5RQfqgByt42IF+
KKg1si1vNuOCHY/FqJfsP5rT16P4KNRD07US6H4ovkqyn3KKd6G1yCKinBcVg+sWKJKKesqJur1L
YufyFJI5qyABozNdrmKBPXvsTNE10oPA3WwNfq09AS7S9/QoQxFx59B2SgaZ3PFA05TBvp8txQi6
gMsxFVRtnAUxzO+adADAOMcqCkLT+yw6xNiSVOy+95ZIry87EEF44LaBfK93v01lmAQutsKhMc02
xy2qvOj4Xbsz97tosOXTsGfmP2bMtbOLVtZYzk/9+u/slxuMe4rTW5p6xy0QSb4F9fAjDPPQBmgN
PrUbzywRmOH+idttAoBfv0bMbZBvA/wOcKit0ewNgq5iQDy5hIp9buGZFe+db2AtVKRQMJokbNUF
QUAAoj2iZeENe01A3YW17Gh1HQHfRHX3tKplHbritNlpWrb5mHvgj7wW7Yt6QOMZPg+GFbprL2nr
2dQkFSYQJMOms3cz9N09BMsci3bAEa26qs4V7a4ulPM3SDupVvJ0WL3PKcDFRqoPE+vt4/guACsm
29JNGDdpguSWrTyCLh5nv435tWHG8O/O8xo7uTbH2nIRUx/kaXsHAADmv3SNI9mrVF/1KhKnpKix
9FF0wjFQWu78VPVqEkCveoNFblVfyL7dDeZEd2lIyR+WV5rqXjPCqY4cqjYjwlg/p3Zgy/iWl9j0
0KXM738l8CCn0UNeBj56R86sxNjDen1V0xSZQQv/p0ZNNycYXkBpFx49VNC6Cc6Mi5KlYbTqEm1r
mgCqy65fT5aimp03Bb9JR2Nlk32zsLBMuO2ZXWEUpAAQIWPbOjz9XoOAblnAif1SeOfJl/+kc1oR
/CsfbN/DF8nzAeE6kPbGcSUcW0zFyHAaiNyhJ5hrpYOJ4vIYVh0CylSS/h+qnib/2Nps+1BFGd//
+OEIpVhs1DgSgHNrGF++9ndvTq0QrsrkBZDy53Pd5t+lfLlIuPwrmE7b11fNb0SzkYRYzBCcoMEu
TqIwiMCdzCN3w1sTCnvEGr9Gvu1AIINp1SyYHApyriPWtG8+jpoLkzucCVvAMKRW2LxEcraJsiKc
GNjZV1V2TUL9jjKGFtAGw2rs072wGcP06laoZ1YMww+kU16pK2lyTRE9gNlE3iVzyAVoWjwDrdKZ
kvmeUuoTZMTFzKO4SZ4Y62cO7wj9FyWH0q23CTSV4UFU3CdvbX9se6SaP32lfN4CGPOWyYjbDVRj
2+NnfQZk9uAzB3GncVUmVHadGK2DvThPpBR9ptputbx1DrXGUWep4BGYINO0vOccDGbTRaS5mArB
YGRd67RAvojmhjs0+vOXgdURxNUUKnidmxsVrMkbzuw5nOJHseFSXieaJh0yefA7ck7zbGhkQvHL
IP6MrBZBn+gGLpw8izfVRZbKSm1R1eJXcdT79M882vFNpUFREzb02Y0rTIUxiEBMVJb0NKizo9Lj
gZ/gtqrd/M7OIb/ayRUg/qH77XI1dNGGL1Qa9C0j25EUdo/A0hjgLHMGflOPO/E4o/eoRpzaTx8y
QKAI2eUJ2QLAM1gKYjFAuF+hQ7UH+2Uno8puK2KnpoZYugEc3aCg/DlMkg6Pe0Ck/cIViXX/bTXE
zMtXqN9KIPSXlGRRbmdPWfwlwG9T6BxEiGJg7W85sOjz0+YqCS8WEBEmHGs7Hl4Nuxbd4EoggKZw
hlyfA3IFkf/H6I/LI/phuCat0NV6G/4U5oupxm3buX6lewrBk7a5SPXpQEnlcuX/hykF/1AHQOPO
FFER3EC3TxC4mjtKSxpvvdYod2aO8YnHEKw1//5UXKqXxVfbt0hV83qmqM2eCsyM/ywFcMaAlav4
C9p7JVHpe/RrNMQvPrH+vmOnlfl8MZcrBKmotttPDMwqRpNI8pA11s3a3o3PkbA7TwzC0vlcT8on
AlRMFbDHx7NUfva9MLPgWC7vWmFIQALao2zMGhvxrd8Q3pcX0pIVaLDjO/aZRq8F9rOPGKYJTVza
xdPUChfLxtWBJlphSfDwHNLsDCoWKDUjmMKi5s1KsMfEwAlmJFIBtBdOP4JD3Gp/oeS+8wVeixXP
EqeW94YZVlugWS5aNw9p5IQMWR3pdTthu/PJWCUc/xqI76yxT4vncmDM/8g5ryfRfSmb3iKMVSIF
DHYquaHQ83VXlJTKH/DW5e7X/mQj2oqWHvECw23PYKvad/6/yPJ779q/dweaAY5zMO3O+2wS5LRr
Rk2xcGTzLmms4LiceNm9ugXV0/wqdEuEFEZB+dXDhc75ODRbjC5GPzgqicbCyGOYHur3z72rjQVG
XpHZ46WOmOU0fvCdmmyun8gd15dkj+HXuCUYaoJLVtdi+YURxRWskNo0HY/LDdeHRJRbtQ94uZta
H2ETvThV6EbiJzwThIbrf6lsOp7FHF6VaxdgvjKlTcK+ZK2qyTQwaF66hdxejIHKfqG2jdoghwkf
dP+VRu+6H5MqNvkyQcpDNkRVMqS5LtIHpGiyW4X+GCYGFiRo2744/rPyQC7ndVMreRdJFndOSF0e
2k0yid9BDCLl3CY6UV+MubGMf1RYAMNqPOdwhxi+AlD9II9qFT0jU9Wn7+rsfvD1fDAxqmjyTuA7
2ud5U/jzksTmukQ8wGDaX9w0+nMgfRkuiBYtuTxWAXrPxGgEwd42CPZIEHDVqDikdookdfx6zpE7
/FelNtg9E1xQtOqVG4So8tF+A7d3jeqaSDuVlEfAxQD2HY/QTQ0ek6VWl+ru3c69oiQarN4W9Xf+
Mmlq9xrw756ov9chEayBwbIRH80jJytwTyT5lwLuDWFfj//U7RxpJpFqNZCyEAzHIoPOcH6zx14A
XTwp20PqUfSwrG9MCt3K18bj2Q01qGSat1iNql7uC1jL0lkyZf/hzgVrlVt5GHyrL5Uo0PEg1w7x
2us7I80hZd/lZ1Yr9XP2wtMoHPGT/FrUdMNS0wziO69VAvKcX8vzStmFXIw/rQVTUN8naz8shb7b
hknbHMXj+wIIQcQdyNeQ+89CAHInPiuW4ESmPfYuFsse2YBkh9TT1FFfoATRvzRmKYTT99Mh4f4I
sJszD45zHZ6NsMuggio+vt7QPD5WFVwEBxzB8fNZSS6ZGVRBAoCBfO4JCGJspynVHpEoN3Pk38p2
+Zecuk4hBmn5iqcxGsb/knos8RtTk8AliwmofyLlJNnThUd53LKX5M4IzH7FatDxahzZ75qBD13j
RklBLVFvIAcP9avTRiU7LhGdTHBeP58XLa3zMF/NC/BXGRa0nqCQEczMdr9095fPWAooJ3jJLSwo
NuC0FKfdy1nf+234cwnHP13tDM9MGhnfjPjqZex65xpOhBlFySS3LpWMaQM/XEld4j7fwkrNKQXH
cZlWpjWb+AP781/JRRQdggEQ7MNkilHGeVuGdxtpeN/QMpS8UBBatBUSARrbJ3Nf4rXg9iUzH2ve
eBvRCtynZKIQeGZOOvgtBQ+I2ez2goraoAu1esXokiS6gzQ1MAXzakiyfZxc14gXjw7m1DpqNien
UfVeTTTXW+0aRIPjf8oPqrJ3QqYpdLQ0DVCzewAK//LFNChwBNvYrYMtS8T0CfAkXWcDKi7mpJbE
2UfqQH7yuNdtWMbwVjlQdFZn300iVQSbGN/3erdiPE3aLmBMoYUumDfO7Ytt1zfIm1MNisDZhOiE
4ARUNX2o27jLmWFVDPhRbgt5h2md4j28zFm5COaQk4NjcUUA6XqKFikfBf/7wOB07TI/F4+igoFa
4iJP0LPdKwSK9ystyjVvS+1jN7olMVJW/aQI2SIOGrjpl22TxZBek/PZLyztjMMsvyCfC93AdJMr
0AkrMxlCEN3+QnFchkWlQDgMy/ZA3oOmoAzmxdrJjKpX1rOAZFRZpiLlyJmMXOP4VG5JFbQsv3AI
BUSCIQ864kE0ivuBOtFLp+7c0EiYjrYGm6o74otIfW3v6znx1HO72oxNsfSP2P6VK/SRVqF+lFqE
1utmB8YTf/wzrlzJosRn2RAyd1KsaDH6NPYcJY4DgN2PvEv1xf4LQOFBPI6FiMPaA7tG2ZRvcwEH
nMuO0/DvVe4l7B4tpANvqWZkvMWoTp9ex7PwPufGGNC+OS/jt6EEXqgQz9ORJZTWctsOZF85O8vd
tk9hKpHYQlyI2y4L75zoCHPfhRJn4+4V7S5k9LfZmKWklFpxM20+Ab8hS4PrZbKqtu5OeDpVe1hI
yg6hwXngzvkCqSuh9mbLv9nJW/6H0TdIDrJbMRFoB36GpYRPi5woisPwAd4LHyj5wx4NXOX7uqih
I28KcbRmBnS+8gjVkxDMkf481H9S+Q4hjww+EekVKIJBm7sfy0Ua3UaPUcp2GmqI6WCDt7yxceWd
Nbu5forUwkpFE/dbpt76HWWqjeH8kjhKUJsgvrlZlD2Ul730YKeuSQawn9IAXWuKh3GHTyEo0xO8
omzOS3r6YGDZgErSvZkBt3fSP7FvnalKK4EiOkBftuQCHFWImZjrDJDFR+wKieRQUkcFOM14GseH
zSgXU5bQElFfxCEmMboFpHYDOCYlaLnYU9AI+iexxWai/H1T0G6kEuchdNKyBVnCjl0rg3cvVM3f
kjmY640Cs+aqpaW7xrbOx+SPvSTnpZUX5/xl4XJng5OZp9VwoAaGp+vc2U6Pe4rUR66Xt6UISxG5
e6hkuBX8TgGmz9Jes3OdzbnwmH+z397n6di0BeUQOdW9gpzBgXJcdfN7e4ovbx8I70fi7MTjns9e
SUwXozuXpOgoLudqgxexJ2chjhq4+e9fIDVN40L19mAzSmvB+ZZ2peuYuG5yZBFbhCPsCD5D25wG
q7UqzEtb6aujXLJtvvlLlNAuQ/bgRPmBsQTUur9BQMScXO8ykUQKuBpHB78+0zwL7paoXeabvPsC
7hayrsUpvRq3rllwrtxx863ooniyhakgPtJdLxtrjWxRqesbJT1QKZIeCley/QncU9DpIMvj0oav
LR39mp9Q8hV/I+Wsz1AoV5usWMWXkXgN1pQcji54yoYywLEIoj/8Al+gYvwDyVn9ZBTpbXOla72V
0LmAnl+tqoi7z0rxSZQUZsqjPcszRu6giKKIwGC/CKG1HreQ9hNvZbWwkrzpfOQbjF51oY8tKOOG
ANYs8gip6+e+qhmlhc19i3pKctOO9xw2FW+HPJ3dq2WlnBRoIZ0NxKkE+C8CEusX7aZC1bByB5Zf
3tPJFbwuxt5IoATkuj+CdYqlxU7VRgHOZZgeaXWKGN/r/6+7n112LgA6l6vZvTMXqctpkl1aVQp2
8P3tqnqmCscx+tp+fRabMdrnOiHtsHy9RCc8Zn1h+EJ28hqUIATwH8eApYJX/iSJsok/bx06ZesO
yuvuATh1LQcGe4XiviVribPtP2NcqlBG/sRwZw9fa41B3oCJsbgXEGcr24D8tFKCCn/EsY22kMph
vgyEbjufzFRXpaSU7htnSm883D/xl5WMGKMYxz5XsRZLk89KwpizsLaZjEzyZ/iNCpRhvuAnT+r5
4AkfV/nPWmhPGJJGOf0Jb5u+ZoWeQw6XgrMkxRiZjQ+4BYU2Y+E71nCcfw2B66Os7wW3LdKzuJSp
m3ZVQavgDLy0SwHn2xYnjFf3t/s5kYEWxuevJ07BhIrYePmgXdbEkpdIrGG65rn/EB+IbLVelZjL
dkgn9l0t5upF5d4T/WVKXBRqjQjtrbTA/tLd0ZqYXUbWun5oxu4XaJ5nZ3sQdwyeq0rnPB506E0+
VWAuPuVyugZ3xDeckSbbw+IyfaUGK345SjqS0qx8uyy8nWWUt+yWbwoGPHbRq8igMOzXAU5+l11t
SenRaWqkoC6jXIDp9pdfQcCyQ/kWBMM/Ts2zF1LY0rgCrSY0sd0llj21AKHQV/Ub4WoogR2kRGpE
8kDI5jzSA44NXtLhCN853u7Yv5Cpl96wPlONdh0dw62JiweBaWK/4adCkJYqtoE5xLQWLtBqVqcC
rKXeUghpJ+LtX74AdYLpkFINr7veHw9cxoi65FndnWPmtuvEeIlrZOXZbYQfNw5EUOo8D7lm3mAM
2Vr+oLcp3aWd4jlgWSMJRfW9J45Xn/4WxEePGfcDPpJaOQjE9jCUfAMoVehiq/IpggAd54PT0GY2
vDGZhpPU3opT83D2oSLL22O1C38UBbWl8F4L6KEGZ5TM2qC/ksr6umIC33vDbDECTFJ2NVCQ+kYh
0QNjBZNaLEoDOt6EIBCvZMK01DufGy/X8ydt0teQJopgfXO3rJqJMaZkj08mESWHfqhweKWbl/US
e9oXfXdCqqQRQyr5dsya5K0/gN4sR4JcfeuZ4XLjAtAAcpb66pNbbeI+OAxNZ1s4xZfZjQHe4XCJ
IKk2TuHI6p89XhWH5OYg/yeim70lytW3rBpfD394aDHF/IJN9tyQnMQVRPNOd8Wo+JPpVXy2phzn
b7RYVv+xGA2Pj8+sjhFL5Z8blFhz3lFF7LZ1LoxGnryovCmCd/WIHKcEC9uyvThEALc/pW9/fixU
2MsLW6LpUhWBP1jzbIt8IVyBhKkV8IT0UGEapk8ogG/sta6Vi6jbENIFubDJ6sI6v9erI+Kcru2/
I6o0eiOR2DLAdT8j3kO8B5v5cPbho0ymEcbCR7YizGU2N1CrWC1YOCY7Aax+w6k8OTMroiZrDBHs
9KTDwEhNsOElUzWRnqgS5GYB9WHjbd7aEFrnSfLv4G0XavR7uloo80xtgofzI/oPCF++voikMBtG
QuOlCWIV9qqTqHL9N179y7PjZI4O4n2SbvRSFz8gblQxyXYgp3BA+NHzzLVSrPCCgdLkH46inBFJ
JTL+9RLsqLsp3Vqfrt0uspIVahIQHrqlP5LmuZMZZ1Db/pCVSjQ+H4+u5PRjLR4BFk4LzlGjJO77
pO/7B3839A795fZNnImuiLTlvlRK4Fj7U5LqLD6HZ4UdtyJXI+noVSIXC6aqfeu8G6HkqLdYaVjA
xz4iAhpZLhIPvcnrqUMZ0xTky4isRaHjq/j6Ba7/NvbsDmTrFfnrfx0s1llskTr3cQ6Ziy6UCRwF
pSgoLSSKKYzZNNxXKPYYXE0bmmP7W6cNBLs56Dv8uNQmmn67so5g/ZKYy1OtZoKG3UhdCh6zrOyv
SvpMaouDRLBma+zGzLkGAEJT1lzSasrIa0jDDsQceMjY5q0vcKV7nt5H6ASCENtmu+mxEJl26eaS
E9t8i62EW0kQev83NbO269DfWsMbgtHtmlivCanIUkxazWgabQUNnYQUFJda2nCKy4ORcXLFUg4j
m7n6pM/pxIudRYGoY0S/eW7VAT5SveQSB4a7Hz3Unmoxz5J4aYgfTEWrMxlYMCr6iFbwK8kUTTKw
/0zZWPjGppGo6D1GOg9mcB1wljqHhMDuj6thMUzHqJFD/CmzM32vuuS8J62maNas4OMI4pqM5UuC
jYCQ9t7YX5kFt0s/RLJFXFrYqnErP9jDg1Ft7LQBuFn3b+fbfgOKUHl2l5e2YgRdiaxSiYB/hQWp
P46G731Pu3fMwCGjOj1A0wo5S5vfcxKUT9x7Ew8eMvyZcYH43d8Xw1RRjUllAVOu1PPnYS+SyjS1
XeHt+ZeYyLmwOeNZ6yNfLzdjWnf6dyJ0s0moZIXZAIj5M21Rd9loW8ld9nBPUbiD0QFh8XmJYGTQ
TxHFyzsNsEph1CUUlcgwBRdEP8tb+xMuIEl6vh8jqtc03cExtdUfIzd5eU1mxHsYu10+cq15nK12
EcR/PYC7MFiLHWbYUFSrZQRayaSIPN4wl6nIHmjHX4ms6Mygc5YqcolD/vKRBaMJrKLt3ntkUrsm
xdVrHRE0LhSVpfRq8F3dwl4bGOjTMrTYK4EMCUbAM2l1Z1LgAZy9cfuBqCHv36zJ2s2KPcqn+HmT
x3QUQiu4jg55ZE4fA6OgmMe9SG8jHutCsiVFEysqHHB3sMhDdxzXyJElV1okYz3H5SkumL3Bgzef
8THYnDYLUjNMH5nqeMnJDUEnUqRgVLMVe4aGVFz4PFtUb5SlVRZHACLQrJ8ACHGDyE9/m8AwoxeK
w/H471R3cbSTtg3fLYvLnTQgKpBWaBJ/vojiXtvbSaSdRHWcm09raLv6a2++OW5e2asks5fcpXjy
+73WSFlKvGquiBF6zNdWvF/iyrQwM5fZ8WfM3AUYGmKwOuyQH8/aSRc7LqyP4M6vqz0OAp/IfT2/
llYdL4IEHPI7tlZN4J5Cos/Ic+BsEFXVPOOAezvMvZWsr/sgOUv8pO4z+WjLFRehZxKIfR82oafW
YJN8WPeyKCSCaygc7eDHRY0EO1Jql0xpGgYAFO0vhGy2jkwT1dXuBpjKtH7FFmS5lQjwsp2ixbG3
0CxyrCem49TlmbfGpFt5h9b1kn4xzQXSD+YrYOLDGILLR8sfwABGticXIfP7fwmLcf0eZDq+p8MR
WNF1T4BnPjUHMmaZFE+wSpXM3IPQqEQLx7K3Wn9EIDSUyPKLVNQaxXEG1xeLkp9dx/+R3DtA9oj1
wtrGvBCe3FE6YF6xYTWl6SIf7zUoNV/kLbAxse8td3/Hvf4ayjJU535bD0xkPglgmOLSd9qD3jRA
EQsSP+FQL6XIZ+1EQq4ZFKK4jt81WXMqA4Y8saUP9DOZqprE7UICXHJILU1mvBT65mwf9Hjg96At
Dt0pAgd5CFCJ6KcFhsJi8DKF8XoupoKaPZ2f+oicDOJLjXXcCCK51ZMhXsQyYhsAWkbuc4wwjpGn
eb1LP75wo+yJWZypyTlgSuO9PuCyBGQMYmTlW0UrPz6hdZy+q7f0kfeDCBxtF72Cq1qy7F1D1Kbi
er5UPdKzSlyjargPiFljF7ZzmXKBxzRCIHyzFXskYEZh43bzOGZpzkfbsnZR1yWVcMBQVCAQ1aC8
qvrmX8Dx4ZqB9M6A9n/GIiFQo4VwiEU7i2g83F7nbBSN8chkgbIyvTY/quhvoKCzlg1Z0lPyT5t+
+FAh2ievUTGEXBbBLta/7cB10z1z16G4V1m5VCt67aVlII2rvp3aYSrxg0BAYEyDRUwVCXICF6I/
aiIsfjpRG/BJtAymqSYL9brhOiyVyl1yn7TAZOKlANiEuV+cmuu62Y5TMm/FYTdNP+HmWOl6J9P+
OA1GjIg/xXQbQJuy4rTeSmH0y0fl9FZk+ZOLD/dRbC09CB01gUEO9uy/9nmR6P1pnrm5vpu10KxR
39OzgaBDLkv6aIF4PxPak5FyUCqiCODhrGOeL60vkbbSNoYVUAuG0W2uyO4Cm4GzX5DOhWG022C7
tE/U1UXxIcg5ZFG9dVUuOMY0D6F1QenEWDbvDezdJ/WnkhgRYnKpp0V5ggN52fLTGBKcz2/OfZMX
KOyRz7/dXYKtbMIRk8mNdtMw/HqJdkGbtWFuOg9Lz+2XegBdyjWxRFx83rwg1p4VobFrO/pgsgmR
/EfC4mIiV7Zg6TplHyoyJnMMQdi50m3yHebUtYHeB6MM1/YmwiXO2xsZX8RxfmrUqJ0rHh6xfK/b
49WS1bqLav7rDbsYV/ydLQ+F/oPT4XS8RWiLkkTWSFHFhkl2jnVXUI4oge6wSjxBheXPPdWmktXg
wz9IXaDR2ux0uRf4zYm8ijnj7Ch7xh3LSewDlTXInAQRE0o4v8NkoFxT0MC6DfkF6s0J/Cm1DAb0
KY2svDjOxcnpXlONnir2svVj9ZMp6g3wX2I3ka8b8eZ+oOcGeolhQE24Vqmp995qrc2Ml+92uJTt
KmEH/FZ2IKNweWh18eb+P+Lc8hWncAYt0vr7m308pWAbDSJq5+aM51nMCi/zPL8ztLRzwObMo7Hz
0X4ncT+fWaX2KzBYWWWuAETUo0N36hCbM29spNLbAb+mw7mGs3ZtIELqvWA+dPqYN1BsLm12xIYe
//QL8VmiIEeWy7SmwLOiXVIlGwFQS7pjObvu1ABnersTL5tO8xlmMH+t+da8sKVTR4xo6TwTx4F/
YhWswCxmLMBoaFGor0Q6H5DbDPJLNnwH+Kf0pSmgHxo0duNd6fmx0nqP0Sp1uRaEX1yGy1wem3Oy
iT/nVEVsDd8PusahnoTroWk0op4EXKi/mwS6w0n6Az8DP2h8qIrWeeA24lzsweewAhWTkJaLdqYo
jY36ticSZcISuA+D7zIJHHHm2HlNFET1triilDT/Pb16JrES8uzut2AqnvAwC9AAoY3A5kBISqsa
7yaM5AyJ7dBWm9p/iPKXl8qtQCzvPAkFagZuRFmh9Fues/JPGc92k5GWrG6ihAJXiGVsa+K2qg6M
caywtKS090DhSnfFWz5FxCfeRKn07Q6YyOgL/zJoOe5WdLF/ti0lVPubD1r2TPtjyUifchxE8B47
2+a904L7TQIl+eD6HaO+D7afy5ExiA50tosYDJnVlF1JFi7GhJnIXci1uGkteN5Kq93qOIDregAp
g+z12G3GEh1DCk11ugWdRFoJY4RWUe4NLxODFskKvi99huKMh4mfLUo44uf0+fS51Ti75/zqnP07
TGOMuUfkVCW5OJc/4kh3vAHmmQAD/HBm8ou2YUhN1yn04SQMNNG4po6jOmZ/jLuVNSkG4qTj6HKR
MQEFx0oNKjA1epANjUx+jEjYsyYwkzqIz8xs3RKk8r1KR5yGV4PeexO5vk0rU+AZh6mwL/l6Ai8H
LWP5hzci0fve/6qHNSFuQ4d138FuIaq2nl03HG5VfT4iAP41LBuYp4LIM24Xyn7CGPaPDJLVF41I
aY4lpAh06bdk7A3L/DuJZMb5djYRYAmZZ4LxjyvtA9ocDN8cWsEPftgfBqV7txh5S5lFwaQGTV6l
Z1xCBP9EhJHP1/tE72cc7Qq8Xz5lJhvnBqGJ7Ib2TXKtGUZkuxqDZ2rSz8NkmfqmkWPkPwf2M9DW
jhvyigX3akuRiBPgRxhwQLk0avQS7TtM52YJCqrSqcBMgInHD4NwSYbWblmRfsX+o07HSm1MyLWd
mlBZnh1kEpRQMoWX9uM9KRTMFwM96RY5Gvcfg7ke2uDSM6qHxFSIg+ZmoFMkdR25AYOBXVp50QLD
H8FBlbq14Vq+cCgse6IuLmTGMIUK17A5SItAAQZbIaQJatAiYA/S/nIgH/bC1NZNoN2T5AxGcoTV
dSLD9Kn6DpWEWSy2lKLEz0y3+vAweRwWEaeepu3fQ/M0GQt8FRCyUGFu1jsDRKQ9hDWAnXZfsSwl
5p62kXpn9MCUGdxoDmvp4J9D/agJ+uHUPbMf3MLl4z/IAt4NrgioFeeWEWIt674IfjqXENLub7tn
JFMNy0U+7BQzVOPSjOq+8vvjCzT8NDKCnzRfueprIsF/Z18bGKPd7D8Rxq+ZCQ7m5Vu3mUOXeLmp
s7HOvSqBJGe9Bjo9265LpDXId2HMETU7lP2xJSbiumoloebYhZJbMeI08zwLS4tefvlerHbyExSA
GY0j/SOKvDhjoVY/yyMXgP14dkH940GBCKO7xsHCxaOVZbUE+DMWRMc2ibBwwQ5PX+8qguS1uXr1
lu95eWuZSFI+G1C0ybbsC6v7b1hpsDpa/cSBB7L7tpDiG4VmyLpHmbzM98UYgOv0MCNoLlGQqbpI
kWL2BSju+s0HwBnEzmd7RjwBu6IXMXcmK7lteLpF8zmEZphg8sqw4D86BFzp+cjjQgPAwaH05WIS
6lVCaV2ehRcuMrnfDCBs7lBNSHsnhoXKiQmi15q/R6Ue8CQtDceJvdx05TJ2zZJOcDeu4MoZbBqv
Dvx0HPH4qIA0dqApW6YpG958aSVDYTOihN9U2NInxAFBSkxR8Rak+Lr9BeV//HFFz9aB02mkGHBh
qB1WH9HvQICVMS0zUnR9VKJZqoU66CvWraM5WxQyLBwp595YLrG6LFrN9riF9wzzkC+l14NgMbsb
CPuvNLSYROzVCAP56pWDbM2tZ3d4o2eiE0NgXxCpXTwhrMbaRBkV4cmfI7MWDupIP9YWGiAR0o1v
IlJtT3cA+ssVp5ntS0TQzx4eNNX2aaW1PGYgr183FCZDnY8WgFFTrYoNr1AhTndHkVrYTjwVUE0k
ugkzqlKyUnUgLtWkRtQR9SJtohGG3i93tE4UsvldOt8nSLwk35iNYw2zUpTDHl2uEYopXm4AGyka
jKeKEG2orheGwOkB2bPQZczrnehVI4/W+6fZOa3fBWO+PwhmOtL0/KTg3juM1ma9HUmAuzx5Mwzl
jO8r23HRObxTAc8hdXKE15I/pZE40vuzWC7+EEc33Y3V5H2EvurLtmL0z3q/GQgqz+8jupz+ULjy
Q+4mignfBu1mSrJiq8PYwGxp66gf6Si+PLAfB7jS1UqJ0buDsNEVbpXZxyCELdUUtMncb0sk/FMs
YA2nwiHEJJHZBpRQq+jrgP36MD0j5oXz09us5Z+BX+xuFHr+AyBMp72oKmXcdyBKVx1IcyHo4JIm
1/8T75Ql6HXxn9ZuPlLh1bgay7ANwMTWucIYX7yRDpGDKdRabAD/+LhvSx7/2m9MtHKVXwlpS2eu
WMmWuBa0BZzbjrjb4Adkgdc5Jn4G/dnZcPYkO9e34KmE7qyDwnJapX7KIHF4iks/HB7ovyOoicdW
HoLsnhvoM7lVkJpoqMZYdlMkxcMOlhVb+S5CMgW0/VJlF3OBF/paSjav/20/uDRrI5qGwLIgAEbS
2fVgQjKV33PAJ6+ply1Pq8jShkas9v/EuWjhVkjadDN293GpymdLoobofEqVmVUqDP4v8esfImdH
e/l+o4RERGMDgQPzAOm8hJ8rHiZKECULQDMLCU1ItpR41+ST4fPGDYK9iwBnEIvTYSv/i5U9Klu9
njgtoxSJVIBCS+U07QYTFJGwhsbzXyVDB7gKTBEh0V29nm0FZF5rUkoPsWC5W2tfj1zPzM62h93z
+68zRQx7kNE0OTHgFaNikPer9zYjQkhVrD3yr6bkRX9oNtpA5vzWnrKMfNCKoGowlVtq8xR6C3bs
iYlUg2+DVyZ2vdABGGLOaraho+67SXE2eYQc7fLK+HglIWVwnIhO2t61oeQvhisH8NDolihuffgZ
pweoqnaTH6XEhlK7RWVFdlYqIfgOwxF77r98nbZyHNbTqaFFzKJN735YPOZO3xfHFH9ZKP+w0VwK
libMTZt+XETbuzyUfmWorag7pIC2RYfGgaSU0rOS9fhCF+V0LI+svDq1jOyw++1GBeudJrx8O+xO
s6EdhD8q1fYBQYyazdkjRcK9v2uTI1HyBvv20LId1Ti4lA0sChXdX+ANGDLoGIuou5ViGPx0qLSF
EMJY3ibJKhqGVc0XT1F/KPbmqS5oCDsrzUlRaXyfCO1XRqeL5BOLKD9BGa2or5LryZeSeGbXOVb9
VKxpWgRDqAHI7oR7YwXEcZnzXAen26E2jaSjXbRChecygT9h+++78CCJmiabjvAZIEBhbVEFnllb
/e1cEvpUpn4bWWcWnAwbMU+DQJhOV48CQhB6/K9fe8Q8kUDncfbALUTvh0FNpiD7i2kTjvWpDRET
DQyjaAV2ayyIVHM+JRsDa7wFCovJd1EsDqoYjM7yjtfCHhU2Ypz/tSE5FVLCD/YDr37em0fVrYbg
iUYUgY96NkefQLtbyd4OejlTDGUFqyLmk6RjklBNSOqGWruKghZCo1j1+WhMtV4C5j9+Dz7t21va
iSSXQaURHq6SpUPnOhtBIBIABqlc6keQL8vbb1szSJEQwb7O03yIyM9u6vTYJeofeObxJg9WVEYe
4Mlb96G7no0yKCGBRGaH/cLjJoqj8Tli9oJyHpX0BRgP+Hd9nfZNlOP+TQEDXjn8TYa6QZ4tva5F
+ricPTOzYEj6gPvy59uv7fWuOAi9k7JCPjBlCNdhXBjWp+3YEDkZ1rKs237uNCobMnKZe1r4uHWf
x3XJVwTyJ+PJ1YRxHFe/XBWL3lDi13IudQUpMaSFa0O78Vx5E39CgDItkq6On4eRIeerR3f4wuQS
9JUpY4ddRn3juEsin0GJpB4DhpvAbyOR1z3EDYNydp2wC1omyQr3T1EnyRnwrM1P88VBgLL3Ly82
htBs9orm/rQW5WNYo8/F0wnfZi5CwF9T8j41ahQoHJ1WrycyU8ur1bNNh6EhFC7Mt1Dkefo8gFBM
oxoexWInMroe+Vp9qmwmMdru9ug+dwkd5nir2ZbicR3XGbzKOy7GGHRLikSAnI+uRB/yMuMreU9i
Sgx9bwkGqiVZp9aOyebLC+OiF2AF4/tfNeM+0VOiB6I/MR4zK1vM8uT7Wzkn/kCtn1wKFb7DnDhD
jvUYv1iVjyY78MyGYFVNkTx/+myZpRvUbe1E8o+oSMdtDzgbOzJkOLS9cVvKiAQnjuhzB3wJfxkA
3aafobNlDMahgYbRCOziOKp+JFpktFy1Hp/AJQPSbtAiwO8hXIL8ridVVH+v7lbYhaHHQb5GArT0
spD3DeZTjpwDRNuGE2MoSDevaN3eKJNRFkdunOb7iWmn88cmOEJGorNs3SdwRAofT+8xQx9Omrcr
9c+GKyMT9C4J8DBInt9hGWtyQ0Ba1O425Q6AU6MfvOSgmQneIaTPzgL//pd79vq57iPKoks2cRoE
NC4PkuE+NFa0Jp5wg9j8RxXaEdZWLiJWmz0KO2s+UdKL1kZX9QXnZTemds9HLVmjxvAo2mGuJJIm
7EboUhsPkJAn8PCt/G8s53tY+ZUH1tkf4VwohBop/dzOgLd7464c/6Xa1h73WXOP48VYJTQVdjGj
YeAErdSB2IZoG0PZuwEPHLIsay+BN5FySBwA0VhIMj62O32FSxs+dw7gRpyAh3Wif2Fu/Fgnmh2a
YPqvX6smE0gkQXwdk7G9mdHhwV//F5VOtot2GXJtEdSQS7pJTczMB346xaTjVC0o7oGlAJvgeguV
g7GCgigaKkvHEo82EY+JwA0368I8clKlEMbfrDBLV1DJMTqirRlolMRS/eA8GkQVBtvDq5XVoyAK
J1HxMtiY9cUZDPuJ5xH72+iptmIFfezdJv+tbBPA8u98iZ8e4yWsuRnVhW45HdnXq8nn7FM/LB92
lazD8UlwNFs6+sh5zhFOIr2jcP3QKLpzubSWnaIiFC8yUc+RZW8yMOBh0LE7fm4iUoKMNP0HA+Ej
RsXRy5RzNHXh5bv7s8URSmDUXwfZ+jiW8YYpAxxFEikFBz7pIJS03EGgGEgamNhkvG5/m74dzDU6
8qM3YGzmgf/3ITmDaj7i6Ux425eT24Tz0rmEoyaTC22fjsvX2s4gvU4daddVoz96/eH7sKFOU3+9
z876hJNvSPgeBguIgGr5fxTZFZyQUxYoBkg7l0lqUuhMIePgfa95Dsp8jhfQdCZPR1DahhatQ05T
ODQjnxRY15teaj6VAXUk2T8TdVKLzfwJYQDJXgcZlmGe3MNiloTUhk0+1k1SZVPpFXXzNqp1pjQ8
HzWjQZNPN0beuPvY3zr8Vpr64WrTO/dgaxX3GcezqD/XMM7q3bnLk5VCZ/h6B1rqsfxjAqi0xrik
vZXBeZa9sqcXlsv8xodSM8FA4B7ahuKHK0LqaS8nnAhDYrUB0aN8CNO0D3yGNDWgNLGjnfQPlAIC
84tFVb/qgdYqCNwwpb25hdyU6S/o5Dw4q1fJA54MtQ1I+KIIlj/drZGboYZJjk/NUdY1YfrMu3LW
Hn0ccpHr8DrWbcc+yrS6A9KmYSsVt5PiFoT7tiRuimYH/RnSDae4rSVyCKnY+dr9lKHWDmtl15j8
U4QTKFPsBzlTG5HnTUMMvLmagMzWhCTFEiRkl7Z06lO/LX5qfXJ9YOKbeZC27lg2ptDXNXRptC4L
CBJEHldMera/QvgZhIFy2swsgEWkCgCBWuNRh40WpQe5cLq3xBa5OIM9GanTJNGc5UcryzdcLKiL
Q6rICkyxFkaLrdnm3dIMEkcJDVZesCcXv52XBGQUQBWMWz1l/Etn/p026w9EIELRP56nBfejOcvo
pYrcL4MrEs/Mm7/8FyW2AMyJ32UVAyVH17/NnBOTKoiJJdsLPe8ATec5xS0ut8xHXNo4mDyTbU5A
OcpwShCErWEQzdd7IAvDrTChj2CgQGTQIvGhXbiHX8q9lxkHDN08xu9nynktqU8dnnpYmCg+EKFZ
L3A4bK9DSBKynkTcFzVjzcwJ5KU/azW6TBvwywwU7eiPpSz2J4MvgCkVw0g7MaAwHisSUriE7irN
jDv693dGd9LRNzvRNwSp5Z6HrdN7hbkSZim/QCkpokQrQKED8vEQK2YqrEzjKmvMy5L4WXIS2Pdv
7nBOYp80LKuS5NsBbjjB/OAsto3KjY6IWmb53CZsAKX3cvRoRcEF4MRWsld+GOIftcBXp1k6O5Ry
wTItgZEAj4rha+VuPLNawdIxD7zo/XyRGzgEvNXUh3yVOait3/6cWCh6tuJy8joM8zpjY+LzK0Oa
8j8mWZ4Ds5K5z9StANGlTDw0jGQij9gSwQRfc1ewKJ6g9p/w+VaRuVVJ1wtccwu4w17kyP9U4VQP
i+41jKhD+9a6hgHLafzDR9pGM9rjJb2TO99t5PKcogWwtZuPUl4tg5EwdqQBbAZzqVfq4WTxGKJe
/YL3uBnzWEnoH/LQcu+2n/lFDZvyvtW3hxVKif3AKbjkLBhhcclNaKZFwC5tVfs/MqwV63PI0FCT
3bqzhaHd5kQ5rb7TSK37YSxYQAGjKG6LUtVZ2wQeJHzmgWZxp9vextnCnMam9uYfC8/3YbdwEd5B
n1UJ1Jh0b47hEXOjavacNWU02frjGkHXdSaQzuhPCvKm3NcrCfVKqbBp7ZI9cvog8IIsLz9rUpR6
WyQTH9++ATs4WHGttho2cw4CrkE76m+O8MSwxNR/GqEhiW0sdq5Qg8xHAfylnoGFPL40CR4nv14t
A0HnN5zm2N6uY9edYL+ind/clQNcw8E8wymJ9lyuYvTz/1FCLTZ98ekWmXLdnvu1pGHoRx9VLnwp
PbfPQ4+LAMropdtAQXvqkxOmD05nfSmodLA7AQFl/KzgGA65A4g6E+QoN6M1cOwTydenSEhf+N8U
lX3o+vf4oimMJMdviLCVs99N0P9qXEk67UAn1cRKZemf55Mb8tVJX70dopb+Wb0vSy+P1utS17fQ
4BlzCymhVRS5r+l3OdrUotrTodKMFN/tlO6JIEkXvpcOImKctovEYyJQGIBGUEbc8AJyC1gjzSnR
t7HcASHtsVT1sj4FNUlv+2pjJjbP636EmuEgduyehaTKrNJjxPlGYgOxOw62QEorBIZn9+1+S441
pRvh0JoVYjonhuReZqDi734Imt3uplD8ldMxpvx9WokHFtX3aWqA7B/W/KDDbNkHx087LBBiNr/6
6lFZp8j8onsAaAgNmf5JC9k6wm+TCRNnKYcAXVU+w1URKUnz6zh2yaZA2HGdM4Vu4f+hERnHNjea
n8qMoTz45dkCrxBNiDT+Dvu8kh2pxmoxBsZvpCedRWzSs7+dMI7Och2HdmsjwWETyrlBvdm0MCLC
nT6vDoldPRPcHj8TOG2c3v3OW6bCKLKHUNgN/Da4c7f/9HqHnXi0NdtYRwtZ9MQLJps+RHv8rtTz
UM35HwEempfNkPVHLpuHjcLYzXDos3KJ7NbwrSwgSIdTtKs8ISQS4ZUpvtxGw+gykIyUXyPFAkUK
yDB9Z8kvb1s3uedgj2JuBhUElh2qZ7e8kuyMwWAhL0cTf8U0wg1drm9CVwqNT5CWG7qXiVPw0FZ4
VrbSITKy3GBTVOfRtiJ+vPWgOi11TVsIAb+gSO+/mw8xKz+9RxYbasEeG6BuikOrhQh3uJE0WpA5
mvvHBnB6LGTGcazcIUSz53jaSGmdc4Cgqh4HATlelN8p2zRwOpAlnSSTrLrl4yFKx6UAMv361ISP
ylE68bjjeHU51QcuUdeek5uqHowax9t7zqAcfSSFtToOvEROadA8HSG1+ywNyznVHAwjFwJnAsbJ
3FIi24KdyIXmcqbWcIdjvbbmvyDsgU80IqRnnxKUpht0Jo8MGRKmaqoncMy/+rIONWkqclE+1VgB
fMJD6yLPEDARXT38a8obrwTrI+LIv8ZXXarMRZtmzfyOphfkW0xnDF+NMGXHDE6lZCluKa5reO8j
UAX2N0MNF5r+tD4/RR6auKGVY4ebw6I3blFl9WzHC7lfGgkNQn8Yja07WyerCjET7Veh0A+2oBKV
HYk+VBO/sB6S6N6rcW+KKHa/PTcnnAch0YL5oArXmipchk4c0N1XV3flKS9SUR+rj9MvLF3It8jd
qxQFaT0+TEU+EczRgZzVMk3JRVZrwZ1j8MnpeWJMHfIXBZBIW5/hSLJyzBvCgesUWBOWlT2z9GuR
180PXTE5aqFkZuRfGQAlJlv2XpdZLWOI1+/lpEWrzxfE/3DJ402LQovnPI4eJppLiwzEf3w2FZY8
AdPeAcCn4zdvH+VXnZNgbErtTg0LsbMzyLV44pYtb7zUeIUiUk9auqWsavUl9K0n/bslzBfsRGkl
vb25hTvIh/B647u3/G23nlT2rmjBlFqO9uPfBvPmI043BvXrPolb4/F2tviY49smoyH7oNKuFkHX
11k1G2uO5pYDC+P1kF8s8KwvZpbNFTTjwM1NJ83zGnyO/qhB0lpBCotTC8hQuD+5FDHGORjV7Yyh
9MIcA1tBnP44TiG09Dme9V6eHOsiwq4jkbQ+cKp1hHCA+4r44LKjNDKc3xueBjHvFiLCvASFUCcv
7qpFTcz+oX0PMAR4alsZcF0PYWeiL6RC2ZSShe2Dnk657LhZcFb+vaq34TiPxco7RZFFUWgNRlmD
loFLFwiz4BpQKjg+9UHbuiH7/BZ0tXVvYzNbY8qQ9APb28oWkFw800I9N4kDv21CNbbyKy2pwk5p
0lg+Pi8s2k2n/BdQh54kFyNzqcTMd4DWFQrgy82nnHoMlSPAVAbjHQ8MO+ZtOL0cMEL3F1DIiSYs
jgL3A5Tlk7jp1JU+A9oA2Oh0GeZ7PVMXAvqNScCsZuHFE8OKnRPISorVabvPzxLmjNPoeXjz2PtD
fLxz0UFXAGKgpSpciNxL9MoqN17wbvMOwCCZfDsu23HGjBrSA/Vd+mDo/4ndLE2F33XqM0fondrL
RyxGMkGJXxks8WA+3jzdvdS0OBTqvysQPgdObtZHzQg3g+5hVU8CZGHENFGOqCMuNaQERyvEe0MC
P1+fg5MyV1HXfpL4z88d/IMM4bCG1uh36bWGuR1nXZ4O/+0hQs1OvyjQNUCSrpWlJ2AJVXn3FF4E
v5ruioHLuGxmrtUTLDAwij1K1WFBRohvzLbitnYYfuipujmK+w1Tw49s1mud3ULsJSIdWw25jtxR
tHpLisoG4+WLh5G3fCvCxV72tYBRw0hJsiiFCI4u+RyjDj6QqKKr3YgrfLVSwdFTV23VB7li+K/d
djOoLVPqfXQHNlI/EJbYM2buKoYMoAb/Q8XLsV2aBFQTjje09oBlwxK9mPz42ks6mQAuOhw/q/BB
iBtdTuh5xrPtZ06cap2nYLz1MOa3iEavBf1fCuOjV7WGrMJ2BADGwghuoLRsPCDlub+QXLn05kk3
GJ+jNfcUdeXEyTNAy1ZV1zR8R+4l2DcBI72sS/wyWf4L/a9lkUAHJ9wOKGTfjtwkODDrM9wUQW+N
0Xq74q6EhI7vl5Tf9Os1EFl2iAarNE56TKCT+MswYMq4FzAnoNfucYEDHDw+dtoIPBURP57lU1Cb
WeqEaKvKCPfIyx94f+jrZ9UFU8+XcsHYodx3ot1tVXfFlNQEXDnvn1HmATsU9avgL7e+2AaEaA2f
EYuSauBUXcd6BQgzFqgQce2HyfQK6pe5f531v6aV6xjvpLogscQslx7Cu+Lz3JsCxMxND4yX6kbM
361DfrJlyfpvJGdFjIXJJh+edVlgwPaALtyu1ojWiu5eoR97AIBUN9zJESPJ0bTi7B3f2gmhnVRf
5eD4kHAjp2O8+yfkDHfZ8R3twrk5W01qp0axcxFmG9/axVISnGNEBPE/rwa0VfYFr/NAV/pSVnVJ
YFikREDOMVrOcvB3qYUcr7U/5epUhYrK6+NZ6vnSxHexX77KsrCNsf93EQuwCLFWHSgjFKxfxHcq
yxJ2CGTyepeAYBqvj07TrEiUsUH2EhUOZN1dgN2oPi6MiVrQ6ztf8cMu3GNZufvflZ/OgnAXKC77
35kI1Rs3FN8YIyNROIS4nnc0RhaAa0A6DttIGHUcILx5HG3P2yeNVTxPBQi8oaZkbtzoB//smVlZ
IVKdcffjXnzS2kU03NeGEkvnO2hWEnTiIBxNHssmESGeRfyQWge+BYoUNPgFLeHwnZ0CL8ufsRFR
PP4K/flcPBS6e0+KN1mK4khg/f8qPBZMKKFn12ctibm0zivwobA8RLXut58wCE67YfMosEGNDiN3
dVjCI3v82yotGjmqNGAp+dmqfOl2F35qTrK/b8z1VaImHwaRfUtBvHnra8nsvFOWcK8f6a8r6keG
GQh/gYK7SHI79FykGyxK4czjQJZMgLmI3595jGIjzbg9G6aS5jFqvTBLRLzoMgnwYMyWYYmBOy/c
gxFl84ZlfrTdlGtggSVniJMoVrIVGoJU9lYpJyJgIFRfE+/lUNYHb6WTaSi+73thxUdIkmbLiVSn
YlBrWo3OS/Api9EoCf14DkmVeJqjl2CRHeozQiAC9QDGi8FXGdYiluYHXH9rnc/PwruiEKe7lNcv
3zdlOxcSImvvSWo1jxRgQSBezeIdE9A9BemYxZ0p8UiLNuEqYCINmp2nynimaA4Ov72caR1DNvuJ
UTVQtwdU2ugWgWCySWzv29usE6goY5xxPPG0AtbjwEeASfSD8HY25yRxdu+/N6kY2CmMnovOHqPw
6iaqPyqZVWrz5LfK2XmCOUZXyQZsMwC9uECwC2O1x3UoX6HWjlTWi9lPaff9qEJtoRnFpQzLslrU
oufYebaVOwozAfSyr2kIS3x+Cq0yeGP4h7JgOofJT1nwRCIVK1R8G16uFGgys4Lx1RenYn2clfLR
BU00qqq6vUtdHuZAQXQWMrkQnlsnwq7t7lLURwAHjvdBLYtfpda7PP6ptXrQnCyxWsKcrqj1xdso
TypxGe384+KWsazSald7I9y2Q8UwXc9eKw1ayddRSthrt8yYmm3IiGYD3Iz4H+ZDdsugHkYZAKYu
dIk5P9kqRX4YFL86yMu7fkZ/KgZE7LwlePBrirwRL6miqLlwvNkuHDl4EnM6vDNkdPEqMc2/RQs1
8m0RMpopxlmfwNXPjtLxQGCo/kXi7GAbHxi2ygNB1riiff7vh3/UZfksDYF9xOxZHHRgHWB3+3+H
GPV2pWRH/lC9vKHBXfQzxY1uQpIJX+q4m/Rpjp1DjGJ3NJo6lvJr5t6hI1b0qECpONrXVAtfFvHR
pvsnwzA+eFuaRkg/20vrXv1mTqISZFKhSAMc+iS2BypqqhXSnPLdYPnTGU1zoEtEHk07rNAuV0ns
da47h37EMjFl6VQZxgZT6JmH7letAdO57VSAV+Q6PfPoJR95YGKitq+bOQKNKm2UaxGn5C8JG7HN
t8aQQ5Ts5ktzI5RrSkcvZlN05CFyD4gTL6ytapPEW2Jz+lM2S30CQVk1VZYrYK4cocI20HWNl5zr
y3ssE6fSVH7yj2N+wBuJ1qOwJ6rihaj7HgcNfwkgI0wTkmACwMOyTjrWk1/lYHv66T8TfrQGI74Y
j5Jcj406e7w5amTCXS/HhguRzuYdKfh2e2VXrlXi8OQC5DbSyj6YjjvFufW7Kfy905fgdqvcYcf+
7zdZA36sZxV9wc4cQC8mMNjgXq+31tPCPNBZoxAok8ZiBw3p/lk87NaFZbu5IfOCw/QZUO9CMOeY
dKOd2hOpmusKsNwB06Gwz78rKDxMxXFUC16YFskrtkZ39huercdSMDzVsGwexT8VzEA4iQqtEDhq
5e0wvleDpIMq3eCNE3hGbMmeENFZBCDdRFnVNCdF8xqmTHii1WK0Jp+iaX5vZ4Ls0mIGxwDUQXni
ihOsUeDB8bR+JrxcgoVPtPXtEgjG4rV7Vz+dABQFXolFXAeSR5hMM2OwR0dl88PF1VeLDYZ7CqG6
0KnXlfL4xyb9+fy9tQc+awqG8pAP1kk3Hl5gAZfPiQ26TUhSN9LKC/+iDNEh3DAUxwyR5c4fPO+6
Nj8LUnCtJNQeUf5FNMkfI+jOSEZkkzMLEasVOZ9fxOs39hXKuAvEmKiKdY4B+VKikfTRvNX4t54B
S+o5TJq0V2Uya5K6ufswXemh8oHHJIx+bJY5OHaghAeRopmITBkQz8j5Zn9XPhPBssmHH+D7fGRg
WtGRQZLetWwmSGFUqUwjCPwkM3cr5ojyCDa3OcTWW9MRxU+1q2t9THajiwKWkAeduOQ4uHLWN7bf
Qb2OZcPAbBCN6a0WxeoO22ddTLJjd2kLUJiEak8KxV5hVDZgKptRQhtgaXiXixttsub3W4m7TLKE
X2An8WcghJX+iBZGG6Zymk/9YwCaqtAQ0wj7EdP/Z1IuLAnZOM7oxMueeNUWkLfjMLDiwG8GaItU
eY/pn3jajH03fVc3gWIHhnGlOQVho8oWrxh8ovDrreqjrliQMVq7l2NYwyzlZBBByqdcvOsxGCNG
nPI7URksEJs+RawGDe4P600jAAKg7suDdYtDbl5bNbGjCSrpgvmIZ8XLI0PWCXoG7W9vGunBdN7b
6QFFhjsJQfFrE7A7ERMP59PdM8NgOIJYpJTwMayigO9GsZW4jQmx3rd2f8dxRkcWED72v/0uKZEV
8sII5TFBErq7UaesXLrhBXQBaUX+1kLoZXe8/5rI6wTnmbNpIdW6P1weM831NSzpVcb5FzC1KbYS
/ViusnmO0MnXlf26Gzi1o7azYgRR763wA88kgPiEbjzHQF84E08V2G6RqnBvkUYJDxeEvS0OKfkt
t51Oi33y1Otbp06DRwwzJqw7WTbXB/pBXmhwgA3XgM5kmLbA0h7vy5xu+rIUaR1+yqCJfJ+1bQQC
Btcj09hocsp1nwKtEzFAgS4R5ATxfua/LUtJhE+LGUhAzNlu3q5oxBK3ZBFcvASfaU4yaM5EvqoM
TLOoxDZhKNBtV5hX5KNbdv7RMNzFitOvNVVBuMrwOb0nyj9BDPZLKkq3qc+k5aqpbNcCKZxp92pS
+B+Zhbn6xgWZ3FTCOSjlHKpg3+d0sTYmmGhSBwcLZgOVJDm9hHIheuzuGCo8h6zMvguuKW7e3egl
yku5IoNyHfnwch45PWSdG988q/3Z3LZx6fvdy7x9dsCvg2VKXDhKup2zoFiPxY7YP+jF5kyYXj2N
3DU1dhhjvyQ9BjxKtKOqx0Z96gHUb5wSeM55QQ4986dBOZLjoTcSUYQ3DKMOrHTUSkzNcJ5HtcZC
k0sOo3RoBTkLYr0p09AHvN6Soc1SUe+RS85HpIadDKRZ88wiAejVAzEcofb63QVuERikxAVbNlRz
lW7N0nY06udPQSA3T2YbVtdrJk5v4jc2nkW3gov665C61wJKfxphZupYtbW8zR6Sal+Dj+DAbxfW
zv5IUUQvOAE6m+9Di5gK8YeVhNotLNYGuCzLknTQjtnk8Uf+/2E62rShUMIzGZPG5Q5dOmkwZ8AI
us7XxGZPRe78g2yfxC/4wixWGS6GYQGXj8fk4ndZZfTYBG6Wd0cmK+k87wrUgQA2Ya8yLTzyt5Ka
w0FQDQwLwIr9ccX1xjxQYqGUQdQF5f6oi9AJVKtyHeg8TVs5vfY756prDQdQSD55oYjvrLaL4zoC
bVIGQ16w/aBk53kIK2bG6oHS0vvH1tNrtA5qFO6RrqbqpdQRYL5Qe6xERIC3uoEkk5A/F1lGKrHE
Eyo4ZJT6XntIBf0Gky6Pv/LSNk8RH05CmhOgpeEs1wKnQUUItitcgn3F+t7JRPH9QIpvfseD8gwN
QZ7UwrSPph17y8z/29vA/59r3OcpFaTPyJBFa/VP56xC0LCWOOSLc0bPotoiWT38LTLv7nDjmrai
R1KGkYZQomU0KzdU3OUJzHkqjJe5gQE8/mRzEubrJORsoavdWRtvJRwaUfyQZIig3qc73Rl1Qdix
HtWAfhS7spGCm6q4e7WowPaNOGZ0W4D/5IjDqRcBPnvAYvGC4q8OtlQw17JHX3/NCGwlEbD5Gk7G
JL/AcU2OzrNSYyWrZqcbUNsZvzbrEPbSNTaH0xuouIBnunz1rNgTWgsy0DrMLhroUO5aiB+yFKB7
eA8jo+y+iL4sgSJpMDjsMgbIG/ofar9oM7Pt6decj9CNTFIZSZ/yHHsKnNime5kpzBboFZwq2em3
FsoyCXiPrXFWD9eezVTBQ2ZjZrl2rRXMShUVdOaNN2017qE8Sdbylpk8bU4b0J7+euV0mJOZ1/M2
Vze78inuqR6ho0qqNQ8vKHD4h8D0LuOESc2BQQlgM5Euf+NAZoRmpiJ8bScK2NX/MfcKnZhLX0sz
K2yECD48OC5dPiIA0SJnWMk+ZOztG7EDD91RsoxJlanRkvub0hMPmtmVrSCQPOys+yZGh3O1A80f
HjmhDn6nm9B2t4x8NSLc0WQGHXnwf99SF6cR6MeRPuG9pyRNTXKgOe4ftJK81Q7IonU6IunlYH/q
yN6zunQgviW9xuqR+zJzCjaU7y7uFthwWC597yVyY0d1hdtPKFdsPhTymPbK6Pf5Ss1rd/ylV5uG
tJBPr5b7jL36NYRQI/vdgvEFjtYl++0UVGvISsTy1DztdzdSmTscwPAUKL9MF8HDMTKr0QFGENu/
yIaEPPGus5yvs9kuKZ8zztPuohb75IxW91nCec8v/Ui3yMRVpRK66c0wntqFSOAB6/jRum1zeqGM
zt/XkjM6zMgdYy7Om75upIYtMIK/m68Rn4BDIrhjQg5QO8UlDpn/SeWHsNL2JqSSDFocgECktUtu
mI+KIHPNN2Pv6UnZaYz0IjW3+14zhY5r8ofSiQn1V1tlsr5TTEVwoAYes72w6bR3coBLfHqKqqps
XxMb0fnxZd78P/sWnSML1MXZggMMvqBJdJOhT92z5tJqWCRgP/IknkrDLoUVzic8Lk7DImO4wnm3
nqc4meAQQ76vWzGAcb8UhEgl8bClORCVrxP6RfonvhmLfEKiyGGOq+MBwgapm0N0BieyiMHrMRG/
nKq38X3lFtxXywEGZSFNZ4RO5HCLAZNGC7WWTzPGwmZPunhQlw6bynTiA+UrgRroO9+R/Xbhum3q
xJxa6GWMKB1BoY6wB4Nd441j8iuSX3S5DDt+VXYBHb9tHBVVtvbzsWh0TCWI/q4lflXmsLoCLeQM
hzLnE8BnIZ7T/ibRNvKpcI0QSRhzk7ZmTaUu+WmMstw193ZimRyJgdrJZnN7GHHUk3PE8kGImto5
3MywWnMibIenbnvlZfUZvQwCjz6VXNUoPyk87yJ0gqkANhK9bPXLfyULo5em2yL3hVTl65pHewn+
f9dQRA7teLzgK92fo+T6QNvsYG1EpTN6Ku5QL67Fe7BmcRdnRlmTKU10tgjiuvJgj5Y0iIEnVZRF
gNnFlIL8j4Fi8p/P5idvjjG+718Sk09OWOv57pcfD+APDQmqoe67jvhKPCrQODv9JBT5JEsr/6rU
6ywYvilxwa/m7J+fPoJcIfaB5GYsbupZbYq3bADZU8ksTB5EJgkwzKnmcCflxOgUQhz+taexuzcD
eTVP9KaT73U3gLacmpoGMOx0aVT2mY3DDYuNvhRz/ejMFYVrSD7DMikEtfVVd7eSpBufNqGN2GKF
GDZvSu3lsP4pfQYnP+jhzVniCqI8RSVHDNkJ5Q+6QLFI2RtRJ8wdkgmg7Sh9i2efW/OMo/QtpKpU
/mA4gOps+kiZv23EdLUlE1gDXuKQIb9+MwiBvu4jQBXFJBv50iqenb/C5xX4eWO50rP49S3YKvft
JlQJN2a/UCRSsaFegHg5GcW4/5dQyVKQd4wwXB5iJDTjgEXbxIsZBHuk/EutVa7bbcMoihduA7eG
REU79pM7DSAMWhGZaCXeiEzIGTPzOBfo4wcmfU5f8CDZ6MfUTQcqYdkOiOAqtmU902JOX8aaJAg9
JvLi+qBTDKNK1u4nrG6R5J0rLVznPrAGpiuCEGVPX/QWZmZQLPYWAwctMh3WuSJJGy74slaulQ6E
/9KVHift2fDtvXy8Cy4Pfgx7b8oJMoko50d1jpL1oldzXoeTEFNz8hUyN00ygWAWuIpwo/QrsPs1
7AjyxZfGyGlFaEKkRsD43LpHLk4XxRvQvhB1lTtIiQIMcpZVCpwzLKqJoGAMZuWoJHN45bnhuxgH
6Cyn+vmd++SMXbo+2f9wv34waO6hC9T6SqzIA5l0sGfMsNgfQMvS+fC75NoWocGN/QHOHW2nPKLU
o+T3+a+pCQVSH8Pv6PDXzjZ/mGe3VbPVmmlL/qWUEjIyx/4BlLawPSEJqlm5ZykFNxcR+CWqdVsI
sKbmueScbcF+4wWwqwq/+ZSKQnPH9cWptWGBuUKAKEkkYmyEY/G53wWagoTmFAjQyT2VC4SZALJt
j2DJjEQip6Ji62o3anr0nxEWypduJof7OnIUNhwbXVL3b7aiJg6QUiEZSaJuebgEdgNuN3E8M1rB
m7MUfJ9V+uwTOISmgaYlEBnAFlTTsEQF3UykpK8KwEqUxPZ362Lz/r7YULUZCIoBf7QdDlHd27uN
lOiKtlEwmWFvA0lVDOoJbbx6zlz3SEE7XzDD6hpFaVkYkAuBjwX1OufACEcdcgNMvaeJFZYqXZQ4
Qrzhq8G8lxdtXV/zTQsOHzFSDG9cVHUeBdLIVoFkNNBw0ew2u92QLKhlwq4QBjglJsV5B0s4Yz1R
/GYMkXIITiU7oDS1oZ0VhsTT7E6h0g95wSZtKiF2QdT2fat8FVGCm4i8k5mhTGOCZFpqYr8+XDGP
LvHRh9uxeDYSOYPoa+zAslYYuAEDA9ZIPK6RY9B+sm24TMsSYDLnKG9uiaw3Vnhmn+LzmidntSIX
tXum23Lxpqz1pNUwarpel3v63id1eg8Ko81XO5uaUInqRakCpC60zdMBPFbRwf2Qr3hcNLP6holU
uJt+YD8VUpxyU6dtvMcgMPsXZl+B3WcAseT6XblDsglr1VN9yf/NhiMIfQce8V+OmHEC84Mfla7v
8C+JMK9gjXYfoggrCSK6GHw7TxDcxAxnnOLdUArMRqO+Nxh4FUFJRw5XaPxaqCpMBKv6QD+PUWtG
E0db3jQLZB7IKzJTkUmj7n4bIy+/oiRiexU2jgxb4Ra4NJXBEosHmWd8SYiUBlZM/Ac5X0IvPIqM
B9cXZfaajW0FW0yYs+wMZ1dlsu4ZGpv+nKNUJdeAc80K8+82YYIsldeY9tKwm7jt1/OZMVEDE6JH
sgbpQ63oOjRWFhtOroqH143ghVveBGdWg8tdBUFTvluvi5sKHaPFU1wSLQp8vL4n7C8RSFU3b7pz
3OJzDr3No25t5sf2B32PaNJ+bBjJu83NOoSCMQwdf5u8q9NDfQVMXonhxvdgCzlejzA4gEwZ1YHZ
jU7OYkzPvSlHhVchXFxCwu15dHTFwk1Jr4sRoh5pbJKyhy9eb+PmCuQTrmIbmKZEzCLqr8RkHcye
u16cuuh59u8C/CqYJhz5Ptw0AwJ/5WFzh2cBLnW5hH2arnEtMr+1hANRQeCVZM1RR1y/qoeQr2wk
Bkcs4dedrxrirPEdV5/XTVgtkpYAugi9ic2CtMbavMV2a5PwVWqIc81txdKEl5suYcBQrvoUnNyG
AwN8CxIqBBaV2WGW4JLATXsw8xxla0ilKiCp/03TO+KCb1kOKBe6jVwnr57WXI207wp64b8oE3YE
DQ+69QqMrHYEE1DvTaAf9psBpRTNjQvDKFdfa2jV+svaj3tNQh9V/ZfsawD7qx2TgY+UHB37pB4y
eCxyjh62J64zPYJOsMipwjFPbIu8it1DpYtqt/lR5vQ3gVKSm3/Hib4kvuaJ3T4nF0zwywacpZlB
+yWbsQfHjVOI1eT6x10meWdXeZ0fT6PcDPI2+m6JnmgchP58aUB2p65DiGL9QvGBPPUt4mdHWLUW
pIr8LlZ+a3xliA6CsEm6Vzw5xOEhCYaUF+VxS3tyUzN+iL7QYGLkSETaC7YxOWFnBBNhng18GyJ0
Sv4Xaui6/Xv/7WKAosHd+Wdp/KcIqnXZLk+B2XVEE8RmqQ44gm/bnuEPVt8A6dl5nMOEFqVOt/HH
IqAvJ+p2nPeafd0DtnF8DmQaewR0TPhwa7iE0TPxfm7+jsGlMAkQ960b4n9dNqgQHY0OItRj3Fbw
nyGbGCZrfjtHY7xAH26EHvICRYVnpUhkwTdr6N5cu2AY3NHjSUZuOEOXybRxo5EXT6aXwAZOP4u1
5JYBWOKB5fK9Keio9REKvbBDZdrhIYtZhsGItzKNO2SSVqf7Z3JRtAIFU3noQ/tufpYiquqjPrH9
NT/KGLttzzpQJua/hDnHDUt1/tYrN1Uf91lFC+7RFmw3+3oy0UqBM42a/hRjRz7lOsk1LMfzU3w0
biw1+eHfHWaCPRBtan+BZZ3DXWlk4ZhP2ZoeHAiivmJ2KXyrpsPh0awmpnnAhsMBsFzwAXf1nHRh
sI7BNz//55Mii3NKohcOs3tfZMmg6JM0H9nTlrEVBS97CZXmBC6NH7IHsh6BvZLf/nuzkvQBM96D
Ul8ej7dIzjhaEi/C/uemWgLmlxsd/n18Z3shkZeJKjYTcLPLbTAzwbDDnrnsJmZtN+v4JuQokZpx
gXwn/ILBF/N33sWQ3CJyxixPLLjNY0PFR3Z4xCRv1yX5Scxfe5a09mNz0VFRTvwu9I3qsgQmYpqx
crrFhP3ihLntmBd41AhAZiilrvrjgcDgOC350nnR+HoI7wqAvY8ietEITLpfOejxqXLNpl9641mg
mFPnQUWw+1fyLj5q5pc86GhAV4hh/tNXq1Dqn6NIBhVD1dnK9UwVfrHCSw3heuOmqgtkJ6nRtsQz
dQZOoPT17oc5E2mBSVxKkWUG3g2o5wnLK4eEOLD00MVJoMtE/b79Q3qb5+aPUY+/J7EwI2dpefzE
eozcVSH3ChtGTBncwhf9pJBoJCUJZbwHIfrgQgMIg1FJbqPhcwpXCVW7WandmQHqAXKSh4Lm7neC
a3MvYRE8dtawvxyJH3KjX2NxycDjtZ9GZtOSWUEXA65OElS1GEa5AgNnrwVbkaCRz+HK74SGFLkl
vkuM2W3Kz6BSdixUm21vy8v/7E0ZX57SOpuaVkQOx9vshF/tv/mNj9sCpEvC1feU/Vfh7EPY4reC
wGuZFbYuwVNo9EOE3ek2HSJB8+1Jd3308hdOcOkvp8PN3lqnC7NhlvEmvGsvsrU8tfWrZMkqAa4E
zKWQX9tRH/sHInYwcAdRYOpENEbrv9oGgmRylGbScfvkY5A8mjw0uoBaaqVvFRCqSiO6/RV2AviK
szjHYnDXUbjlrfzw3WaGYMpRcA0I6jX4pIZp8lS/j6JZ1WRN4rgbv7woseenWBb8HmE+vhF3NVV2
lwioWM63MWTwlltLVij+uZpXBACKjuJRMeTvwkZeGGHffNs0+q1KjsWqcwNMgcHwYp4twYUR/cLB
arLWvzpRaXnLGb2xsAmdjiIDKcpe8/offYdano35pRn8VTqd1QwAuQS4OR3D651VxFRUo1a0Zg5k
hXHIRkl8xp2yyeITC5TbTt2YleUyrHznBGW58gT4mWf3OzKWYSQqadIRgVPwJTFTMwpImyUkqJmB
78ykIHvoHXnUqDJqU3/hZOPMPZuumiXZJUhPl+7UJQbWtgm746Efde4AQih5OXbdGd9687CmcL1b
cbG7M46w3GlxahJZ/wehMQQe0akEG1Npp7f6EhP/M61JH2F+rOebWmNWLkIiFXwHKluSzPcz4cyf
NGvsX0z6wLw5wPjf/z9wJJft6mBZBrys54i29vnzT4GqeEt7yWGzXMuIFErPkb6jtwo0uopG6XSX
gYNvVNmNW79G52+mqIOoAZVmBeFaxFax9Gr+8pXq/IlH1lGJ+pfgepKch21P+cXnoRVQEQfvnQ6f
UsJ8CwhC9GAhntXL5z/sPIaOfGF9p6/7Q/vRh/ReHY6CQHDpahr0CvGRGlnvrpYiyx22Llq7AHdc
SO5tOwnhytn8YDsyjiHbvKDI7EZ66gavrsS8HQ7PtUEFbBXQy/6IjKM1dJsmPksJ1px8nLbsw+y4
e2kAqe9JGQGOi/GRnjAU3wggD/apjo3YLCPYxosnVsIJ8RN3lt/TAiejSASQ9VnCc9AZ0IOYuQkY
+xoG6VIKfn/n5ucL2UtZLRBST+TtdN1xqWTLkro1/hdcv9GuLu7/2qMfDJsjRqwTABoMbdBOM4mj
BDCIVlUpU1P0r1tZ1Jo0rJE7vJBgUvDqxlVFT99WfGrrGVoWezweWHrA4T1x1fyYrtMWHhlc+wcK
Icpj2YZqPQxdkiMmBEIhQ3YjOCzTa/j4+OZoCLshjTa3JbGGgG55JY5CGwAQ7c1DIM4faOf7xuys
dv9xkniIzsFm19eIvVhLCPQPZcGmed/Zhwz5bkBTqSQq2Jvxd5MuyJE52wZMiodkWg/B6MQltkLe
FrJ4RPiKF+7EBTADG4rOnEWoCPkllc4fX7x4GkryPNzEOiOdVf4VmyEgRzTUGUo+flS5vyxAPvhD
zitTG18jvVMXkVzUg1Xzbf+lhP6Jp46MWHFW7Wg7GKgweL5ihY3zQMHQKrFheQSFoTMajcDyokCv
CyjqZY2JyvqhYkHcCzsw1EhZrYCqA2HVKIrJ7tnzq4UKIXzoRSkxyrch268ubHeRIelJTAeoa/wJ
eaBRoL5/4CRMbn9jhjTlewlLGI5zQNJXJN5V47LiZJNL4wHY3yhn2U+n7RmWwgkzGHUdkFK5YJlt
Sd36YfMKlkxnYu7BIToMKXSdIS4YoKOFxN/vWug5yTwaliDF99Glk93VTXzJ7Jn+htFxt0LwNpb6
/ZBVPc+fp2VbVVmWPUShT262shJfQdqsR94SZ5xdbF1of4kkcwDRACR0CZRGe+DVcyE2VKPk9ikO
B7P0A1fmbJ9XYm+S4cxD8sfHGDTXqHevHnHKzDnbpV3v679ZE3Z9UkZ5PrOhZJPoQx8FHRG/wKC+
in6gF9n4GKpSiPMHPmExiysQo5hLHSlKl48X22HdQfHLlG8hAXHpBb48kSY+gpFxZH5H8SKjBh/d
vN4C88IG4MWFxjG79AV8TKUc0hjU+ns8goM7uSt/2ZgsIoy/eWxFSLsNvg0aWa00r8Ik6lzGrUsx
BPs5z7pmVWBB0r8oufnxKLhVZULPzpvJYEDVs6Kgjzl9xpbU3e3prHjQPcd42DBXlqcACpyiOlVO
56XTjV3N76PRD5AJRkJFBhx2te3Q+AErI5jrmJx4j3WFGTtUtDDJIAjZs0hjUTh/Z6UJDouge57D
wUorEIOuumHmgczzrE78dC9DPh+2hkFoQjDGU1b1gdLADb7VdB9691pjEJUkmT5P9wbj/ej94M8p
t7ZTLd98g/vEK07G+VKNHu3z7ySnAMWZpMzLfBz84Je6+BzoaERzzSS935SIcuMw5LjdHk7STS4s
xdKW1Qxa3Oo0WfhPAyNo81+45YlAym8P4sfmc5OhC97hGJES2WIaCbwGLYv2YH+VqqmAUa3e9ffJ
HzoEs1vvyM1Z9oFgeK8RdgCh8hiG/SsoCcvJIDtLPN71mZDvE7OZvkuNVDoaXxDY2PWTJs2quL/C
hs+7P4ihRRGlsl6SGgLRA7S6/HJ3eZTZ6zhJcFq3MTWsq6/6TOpPGuKESMfGzq0seY6TBc/XiBS/
bYwTIh8RLpFq1OEYK0W6GeKjODnFGdvpPuIUw2C9i5pWQOkA/HjQgLsF5Kd5+cxRaLjTH3XOR2eK
1NiknsJwyAj4rvvXCGpz1GQoQp0B1mZb3xlZA8vn9kNwtHH3UbuwVq0lO/i7ZCHJ9ecEZUxSNZnA
KbB5GtQNu6ckCbvN0gFITAk6fq1Zsq0jI7+bR4uEnQBm9yM2MUQFNkJr8DepsSkNcgoG8BiHvINW
51mPBakDDvNjLcJuRedimE8COoeVqbdvuMYanYbdXIYAlr75h83ZFr9UN+Gub/xiWkzp90d+NO6V
SxoQNEmGI/LiZDAA00vhG0iDJqd/aKvMe8h86jqa+JsGaKOxtzqk0J8qE/ktW3CYUiqzZa/U0msb
8fJLw90J5JniAcbFyRTMGyBngJ2HqDo9H4PTLRoT8BayiCBL9S/8koIU8POmdUYpp7O4QNASJkep
dltLLPDYPGE/6dpK7Sw9w6e7G23ML5wSyJ5ZUDRfaodoAnPZlvjOPADr+Z5EvnU0TmBo0gFFWyN4
Zu3QjR0MkpIqRMtyY7mmiR6rBsPjkakoQkzetfX4pYMc065jfXRJ8muwxtTrxMzr9mYnsQg2RGQd
lxGIz7z/f1s7ckqLlMIqhlqzMKvjbiVj8765JCdg/8C/lE+uPCsQbhNGTtSs9lVXfzc514f0sD0c
CrcgkPO7xW6JtwoIAKajMiJp0stc6Y73lcfBJRMZLHhW/Fi/+0Eg6jkPFDkpJIQmhSDDvq+AlURa
LIsJla7amRttOdgBWGZacZ9rMuFWPHjNT/4OP+Bropt7L08YP2l+dYL7BMQkx3XiI/pzLNBqNTJa
VE7iGZsF8TTOwGEu68s3JKjc8YWmf5sknghSJBcQ+8ZUEh9AAGIffm7+47Uwfwu22fWbcP1THhyD
1zA9P6wDKbacA9ONxjlR/xM9CoWWqXZA6y/6SIkPyYRFObQjXCMXv6pkhLea7Ft0isUeJWhpW2Et
6HWKX0lVGUbqs9GCIOmoau2yb7lJsgProogWjMeNCZtseJhG2ZSuve/bnyyD4OcyX+5TA+swhR4V
itDpO4cFGgnljCLyLNPhcRiUhHr/D1DLxovN4NlwSMpsyp4THcOhkZYz/A/MgEAXz6Ee09YWzJRl
46pbX6WMASq+sqS/Vo6MG+hnm1gO4u1b4bey4W60p3pdSkSQqkSbNJz691kgSBP/Ir6t8a9kGAOq
w0Svb4XXMH3sxVgMeNaS3zfbj799fGGaeoUitIOWravKRjI4SGIIRukpBYgzuTMRPgxBmsV7hy2T
uW616v54yY3cnX983G4Ipo3UcoFOF9gBqLUH7NWwW2g8FFPmQpD1rJuqBDQGMmHFUP0QVSP/75N6
bLHohV1SCXRoGb3bn8xF5QumlaXSRk2whulvrLFIdli5HtetqSxZBICSn/8oHH8DYRDv8MxFEVSw
sj/KCQY+hkfQtTmxs41eY6KRK4Vwf/OPEjFlG0zX6FlkDSqaSZVjSZBm2qNOKMJj3QTa02CQ4rWB
1y4M8QueMmL0gwd/6hGpvYQ8RRaV2UP3gwQs75c3ooGAHIXIVCLednocHxmRzXYT9d6GzgVt/Kd4
L+yPh7TjPRbrrdw3e90b+l1yoCYCd1vivXmkSHwM2d2DnBpw/fJnkF2YSQykOvgi+RlS1y528hrg
xlBzl0J7VVc/U3OXrRmocbja5K7DBOps7bqkDcev4gWAGGbn0A9vIHwmff6kuIRrKBx9Wp4ehQnE
Q3esB4xnlYCV9MTcHyf7kr9/E/DSeCGI87kIla8cCW4nVTVtdL+6UFyjWF/UCzO7zMs4RvrOPnhs
9jgy6nvOs+ERcBH38aP98XgUxNMmwXc5YBDN8H3xw1IuJHcSTXqD7HM3K51iKKXwYskN4nBij7LP
UV05Po0w1D7FIqoJVDUXkStyvKB8Qi8Lw8wFWO2mah/f8EjSu7HZj55cU/WE+XlEC0HQALhmGtmb
l56hetyiS0dyL6IUyt7SiCzU0qqk9OEK8KtS3uYubmTynzwbpr69nBna66no3mPiS2KBoa1IdSo/
1/E2zVOWDlb+ePHkG9U5wp1oiy/35ZczT/+jRjhWXnLmTGzrSbPTEqInxA3pN1t3jWyYJJI/M6U9
+IcpzQU5vY+GQczo/WIQGJC5b9rCwKFAGSPyM7d5ikaqIj88o8GnOqlYJzndK9Zadzp5bJhRO1ei
4es7sFC3GaViwAjQVQcD4Z/Pw9U5jf7Go8KbFAF025MFH1O4a1k0LGD5giPV1n1McM8XVp+cy66f
2uppXbF3sntcQlh1gZZSPDAH0e+g8ako+vhd3ApoSVk6QMR1fNbSD8lWaUrPmTERYg9IYw4Qjo9+
zyB8I794CUQZodHzkTa5K/UscclxwKP7EK2FSok01UQbGSgUhds8ijGsurYTZbc108yjFm8Q+C85
VBLPN9o5YJnKEW9vfqbC03kARn/VmukrhPpQ3cNbJqELIowZeC9Jm4RROQeV8IhAFgr41yBolEcq
rozbzsN0NGc74H8KdAV31/IVYR4U4vsChrMz+vgw0xPSpsSvKt7QD5dEOPX2dSWjzGToVQFx3f9z
wfYp2VNuqKcr6pmBMYDQEmW0U1NHE94yObRfKVu53bI4MBOA0lyubmCq4hwnGeULWn0jrNifk1qN
00UkTq0+9HMRfcoP4cjXCWvoNvDBvs/cxSShqgt8czT1ZcvwRwLEkwqdvBgekiNmOOiJ6CtuW+AA
JK+52LOlGdggjmsTDFVYdDXT+y/MCn1X9jVnKXF1xHol8x9JSzQ2jzCcXIhyYc9z/H3zTWVkzGqn
oplca+pj85ndMqcRpBpxWlt+jIs6is37TSMX91/WojNb7gQqiLMiRHbDZ+15xTLmecyMJMtkhkRo
N1bP8GtoS/2rRQUeHlhfjMsrfQAv5RjU9ybMdaagR8YV6GbP1fMlQ6smminE1O30ZSYhmB/6OoUO
etHMKEHiDYQQgN7FnTQBElzv+i+sWyeASvfKHawrJ0KKRdj/M8ugHupY9ilSBeMvjdwnH/KQVrgq
9FWM/BPk+Xhbnb4p5pPZVaHpHbQ4G6HYcAnaF1ChmOng+b30hGLjNcQtwWpMBlX+8aJOt+W9d1wN
5nH/M/NHt8EIU7XWYXYJUPh5YFObFU0re4+Ab845mdh4ZkREtwNi592TEQU0jJ4jCuoxs8AxyF0X
anzb9UskUEWAvrpB+phu2KU4lBmEgKmgZiEtcAzjUHIZjD9e1C+sE/vLn5Rz3LcjMLHgtm+Vun+B
H0Le9Rs9cXji8hIZM3ZMizU8jfuzBUCXexBs+a6IKrHxLyzBzJq99FlJJpUdZPdMHZqCA7EB0bWr
oa3F10hQwwxZ9PGVs0EWiRHMwUSHP/DkeBZqkpUOuG6e/qiDg+1V0oNYas0pgUgD6ixVaHYa2N+k
KxOSb2a/SQrQLCZlJJq7wAIxoMiE4i6RgUYM9pnHuLL6UoP6EkWvh/uQf1Ael85PdiQuYMZLuIJj
RW9AKpmgT2bavCS2iGed3prgo57as5WONImtS0vTAdB3ep8DQahBoGwVUHijNBH49Qnta+DXuxZT
Fwdc7WEZVbkNfKh8B153djfwbBI15W/16gqF+zbZ9wefkLHGAzTytvg1PA7FGrbNzLPKLV32NDSB
phj2083AttzLC7LIhmwIl/VB6DRD0AUSXu7vYct4GVdqT+gaNtyi281/rpLv5NJpANwg1NUNJDhz
8CDHRVwbUcElFSQsDRBzDbZKfoDy5STG8YYKHOKzhP4AgbUC+t7AnjUIS+pQ+L7yrRnZ75mu7Omy
9r6Yc0z8/w6y7PjcJBi6qo/ErzdJ937XmSZ5aLo15r0T49tzis8QeKkd/X7Tg5B5/k1IkZxtK2CZ
0eIzqUFCV0K3O+v4v+20Mzq1PtvG2xxoE7ZPGG0EQQshG+QC8gcZlF5iRw1OjuAuBkVMjBD3y6wT
UwnZy5xJkeujdeYrqLPoB2mLz8X4CiHdhK6gH30ItSDxdyUdPfCkLnCmwyvb4y63mHBEeqCYNZrW
sUnT4hVJat3Kcw84EPhfyFRs4SNQNVZUQpLz1/SVd9uv6sc4FqyAShqh1YgAolm9nvnK+pTFSVmS
pXzAoX75viaeSD+fh8eGZ092eS9bYKzV9PuaKfg2F/YAGr/C54s9kUaU1P7PTnKld6LdBszR7pvm
ctrZBQCqD2Jcq5v8AWRwhBLHyarqiHm14FD+mGFwsPqbjU409uUzDKHf0YiEW5mnzDOt63H/APxP
gd3bJ9DSu7FYuK57kwXrhnV99OVvqrr6UjJiTj1JVrMYCZerEwIcYHZCe/mWLhhRXw6GEwHyuV2q
MZulN1KIrjf959AKOnVqImoIu+fbgwAkA44gFrb4RNijVfanFPqVPdDL/s0wz/vrBv0rwbGV39DE
LQUv4j9tv+MDLsfG9R1oiK5y+nOGw98z1HWWTa4kbOU6OMreIuRYFzoyFNFoYupbSolB2Tj5sGEm
NXmHTt737cFFYrwnht3r/4P0sd2lvILICwlTVouTJPBlMcoYHH7j9aq+yrh3Tf7Bm7vfTDl17QFT
7/zwOFExBB2GYP82YKEcjuPo2W1h6uRJCFWkA2Vh+ZlHZ8lP+5ZkunsAB/+iU43lnqKWt2wi3eu6
rDtR+YpS4M9XuVFV1P3tXVlo2BNUekR8B9tmH5SVjk3ZphVAcQYHRyBSxmOmq/A3dtZE4pIOXAGF
G+E/F3mk4e6ZfYNehi9SEXblzvnc+0bGqeNk+v/PkOUEziDp3btl+xYnRRov8Y/qgQh9CmG76g/m
Oe5zDsRCXiU7otMtrLhorsOkdC2RYpb9wR+9hYZvE399UxxoPxtMoDiYo/3edZ6Zeqoxg1blKYns
8l8vnxdtpBB9eHyTK5NKL5ruLxjr0/iXvh+g0izgVYh3UzWMX/dd5HTL/rWIfdTjGJAqkaGQ2grN
2UGfGBJ4bFnOBf7fEB51ClrDE7zvMAthwVb68EbHyRswdwMsifRhSYwKuOcWiGRbBS590Na0Hzb5
R0dq7dwK6fyeQeUrLCi+f8OSF007p6zSdCj+qXfGgqthJXc1FeNcHpa6A0Fp8pttRqXNNvxK9gSA
ymHPRHJqmtUlVqkR2OvpMDwhPTj+C/tAvAjtdCRDSGa+2ycaq2fj4qZQhPLFTDDPBqWBo2Elopnt
jLuj5iSC9mL0EQ67k7IrsnwQnKY75d0GdREY8BqisJ28uvjIZr4OUrb/7vYKJjDdiQROOmto/IGx
LC6jc+itCsmmrqPPQgQXUFzi+VDkLezQTkCyTGw1eSkyfT/pbG3FpP9KhI1gfEMUZTydKp0RLmOZ
l9VDFMytxXJOJHG7AqrkfxKh9u073JyeZsTOlh5f3P54zipddjmV1UA51MU4otfvz3wY4Abv2jzu
DnljZUHZUPKBHLbwUyT/3EnVwuwGy2aiTqR8ndyy8KoCmpmhszUiqfmUpZtSERnxE67XTXUOPBoI
FLrS1A8HdJuEY9MoO44E+Wk4+vCRCmZd75zWzLb6jSEIPeMTDx9jQ3m4St5zbmim84NEIJU4U2j7
mUl29f/i26Eg1Ldl0vpwSBMBLtHr5gOF2QQ9YHC/lwqrfhEo7EpcEECatiWykgxpGS0PBh06LTga
HpGB/C8XsLkDEU7CCCSx85baUDszWwMuh2WQiULlIBoLPWpbk9SqjQg2pMIQ/39mlUYXEvFdfSk/
xajiuhIwvaX5YhEdg/U8B7C6OzNSo9VvmXDEqGs08pss6PzKV8EXHDO2YMXj7zd+hRH9vNyBOFP+
fOamKx3bUjdHdNA4YCa6D1QqPnrzx6F7mO0qpr7e0IvTGTV5SDCqjhE4V9oKD8zrvGnUYpOJXMUn
WV6XSdKSJhHS+6nIW+kpsSQRNht4mMSWD/Mkn0g2GHINmNNa8DEIyfYY+KkbKrKKQNMHp5DdLHMu
J6esLNrL++NJu85pOHCUwGJxW4E8vktyqobe/IsMEQGsrLPJhXnkLbw41tPSXo/NGx76XqLq+Gtx
IZ2yxUrfgrtJCwrd0dO9/ikwIgM+zLZYYBWS439W5VHBdCkLe3s7TuWlZiP0eomFskNwjW8RZWEM
Bs8EUQkqdzk2Yu8AV5KOi9UkeRsbiXzY1kf8HKZd/MY8S8prUsO7z4DV0j6YN1D2pmFwo/VsCyh+
3evkMfCDxH89G/N4pAdCpuo5hc44lZHcH28WvWH71tiz3qmIsAcC7RGYC1QBMF4GLOTbfxwgVmXc
7PdV0BfYkYH/ncqDlfyI+KLQUXBX+ySbu2aV+J3g/RmVXYmJvxWoQsOGU9wWLt6iO9pCg71FAS1D
Ctt3o2vYD9gPVA6V8ag+2m/tBm8QwQwMDqXecV5haZPg1eVWnu1wFTlKmH6mYY68Ce70A55AgOmA
zJIYOaZ4qTcX8kLLibogi5239XuhGGBE4fOqMjA+5E/3MwF0vzvA1Oy3C3Ay9H/1iMJ6KLfKkgUi
vhx2T/+gg22dcky6P/jIuyVC3MYfhAsANARodxDxCrzoxp1Uhnxo/4xfTUT2AXaKdwmrEnBcF3+A
4jhiSuiKB6UPzU7rdOP3my93IbTlvBw5ZeDgmhfOxadNHO+M5m9MXT5d8MGxduPDNHYPk4MpOtAv
LvDn3RGPMyOSus9Xhzvl4lfBUc6kpN3v8oxoHs8OKv8uj+aNtKuUMyFgo3ctKxEswH4UhA9RdnK3
tE93PNJDZdgGRDPf1pc2yt5HYuj9IC4gSUOI+zhMQhPcv3BpTWJ8pDvE4hBfM5gR/0zKNKfg2dhL
3kcUM4xlWHvF0NmNwjcyPT6bhC+P7FcbPUsrlhrGwxF0rvm+V6wvr8ZNM0hdTabfxPm4b0q2Qukd
/Wqmkx33ZAVITh4Peq5fHXz1iIqJmledzlCx74znReSNM1tf9nPscU4EohIWePpO0XcjzH3uBEV7
8r5tvBdKfLoYsWPFDMHDFHNc09BiQtyiwPG+WlgQiAfW45opnO396AZj1UhHPNxCIWEmsgZqw22D
disfZZae4dtzIg6rl4g8tf3V+mQgP14KiB72tXRvPiWEqrYQ0BKMsl5MZNQu3q3JC+Bgh43r5w4h
jXER0KmgCDS/JcAoIqY9Oa4AHrCi8DM0jS+pS+5D1y1yzhYZ/GIxqhwRgYUufElbbLWsNCnCEuEL
QfObIUCN95tlfNhWLIqpn68srR3Z9JfGORZtD/jfUGd99fuadzFITSaozBeXEF9G18YZ0g0DxRxS
aQQK1Ag5iDEbCd4LXOyiqOGVCbVg7CtPcQLYddtaLvXRwiFRxe68hgoISFjJHdu8zvDmqVLiKs3F
XQWFyIwmM5K1N45YQVjrxrOaaErlN4/ca5Z3cvpxiAQ6tUBNuKcDzOnYNuO0GcXeQvHKvrftlYuy
2Q6XIcEdnbFly+l/3VJ69VQPTfs6Fwv7oNatwNSrD6JGmXL/CMAwXcjY8d9WSjIP+hn3yMeifIzi
76qqdtZ+CDmqgkJ+4XNb3noNIl0P6yYmWXGh/RMcaDQxRkKky3FM1pBLSXcGlPPAaXcZGXRh9aO2
yne8mX/JK0SwQr8jtxMQuwxeAjLxLjZtB7R6/FDbHW4e3wi/8tfunE9cAyBvFLLyPD0Kv6fr2kwq
Vx2Fak73tiGhqdBWaAa45e5N3aa+gJg406HxhUlJxOmPaVs06Bo5bVUlTtL0h4i0uDYBciYVp+Tj
pkAaNOqnkU8Vdq7rErjBmfLcx+r4kFeEYKktssvY3rEg5/qOKoRWEnFCO0y4PtOwKlSXrO2WzzvD
5cspMHQUPTXZWYbDNTYIvjHA1bLanhI4bk3DtNjAmuHGN0PLc9CgI0Hqlol3S2IwRq7ACSC1PLOg
IDT+8sSPJu/Qx/GUHCwnh77wii98+Jv7wNI2JIncfQB8RnBZM80twckRh2ZHBxHxcHcbr4t1rYBn
yiaZxtJ6TZVphQ71sOtox7eRXK1gs/r+OPDHyhDSWCVYMcbsYRO1G8Su+TosXbnlp7pEoDFLizu1
vTCXtFoK6auB8+OWXmTPfXSYPOaODL6S8d6dG8P8+mK9CTZPr3a+OolkDGmvAYGBYnMufuzxuQWk
vkeJjR3lYNhM3sfks3pttLjaOGC7uaIcVGJ3WbC5BIKn2dTGzFp8o8Yu/TSINtKsCrsONwIp4exx
9dVTUO9iyGqGEjV/vA8uMDKxgF9gDTvkDD4n5fJv7817xFQdn97YWoZRTwUyzvYG1GXeWd0cpyTJ
i7rV+sywnw3kr6iWTUcyPxKjIfl9bwx5Ngfb/sK9SbcytFEWGe7BgIyYQVV5ej8Z0c/VaokkICjN
MUhKmSe0QoWQ7Ubh9QNB8oxl0OT5cIPKZiUMtqG+z/vjv5bIa43c+QprP1NwpTx9c3Ert02nHVTu
Hf1jxS8it7Oa6+JOkmw079KRRU5CgYj+IgHE9x0kzuClPmOx2kU17Pvg1N6q7bJlTBk0g/QVq2VT
XFtm4zqky6NV3f7aRtGk4cdmEdxRNp3eSJ5FwAgnHAhqRl3fpu/5F1WYmccq9I/u7ViCpuWIocpa
RBk/K+iyM4vRjZZBkq+9mcCLaWQ5zafngH61iFjyCLM+IkZxjmoMmAPzBOVXwnXjZoo+9WIO77QF
QC2k1Cl5sKJow5UUbH3NSkMIbj3znIZkLVLlQAYg/98H0pQbJ4vdxsuYwnKYh9kWGfZ1jmxM83VL
ZvoqWr1paab8gNXK1L75D7uu0ZhqbTQRhEc4PCmGKy4emndK4inIlDdD54mxfhvYdOjX0KI4kJ8z
UX3dH7FtIY79t1j7WKxuPt5cModdMPByFosvlzmgoaD79UXXY79q0I8eUa5g06Iggu3M6vR4o2gk
uItWh1G/9uuSAvLWxJdR3B5ATfY7veVa2U5VTi7kKPM3pLl5Dj4D+ud+tou1XCoMxdTQji6hOOWy
O/ZUirLp4ihLCN6ufVRe3/M5WyDJh/yzGK7k3EYeMZUwfZ0COai0Fe+PCFAd7xO5hDcA1YDXhDHp
iX3qOsBbhpGccSxJjbuGlHzgfi9Kw8pIcFBfMX9LsoNTy7rPVwgYB7bXKpkAW9mN4tdjmnK04NGY
RGSvML1L8EZ0YYUkMQ2NkEIMgfmDw4CTLE0lzh+kaHmDWar9VDcvTwnYBhv5zzcJIjLlcr63+KBT
x2BMhwz9g5LzhmKNQV3gQaYcO5gfybIU4vLvYWj6L3Ug1zpChHRLa0UZCFJvCaTs58Od3AP6ieh9
S7fEiav0rmjde1NaiEbAzIHkgi9A01uZSsASIm0m8acbI9SfmkSM8pwus+FPKMhQENn6OQGh0jnB
oeNsUP4igRtuPM8GfY4HvNdj/stdPCjGn3uq9aMR7Fk3Uwd5dbwNzgoK/mpKs0KmS+mqToFccAcu
ALWCWEdBX6kRVwVtCSsPg+JbWer+DVhB6w5z8+sjXkI3d57XdZMheVb9XKpExO2MOVXnaoeMWPtz
7X2F4QFZET2HF+rrzTSPu3BE9GfOH3a7EIU3f/HeLRYaJy5cPlranciZbWDazldwxGOdCm1ZNWGY
MvWpCeZWHH5/P1ink8H7hmwcdHM8adybFtQw1q6TQHqbc7M7PG6U9dgEn64r/FhrMD66XZbfvJg9
7TurE15vbZ+R9E88TDelIebWMtIUuI7xroZc5fzl2rTSR6dVzm0wNnFYrq756Dm2AkABlsv3QQNY
3izirZ+sBtY5fEGeYVpxZaWcUFpD+BQU2qppLcGb3kHRgQCj1Gqw+diQdu3Qf8BL0EXBRuAzO8nV
+HeDYPmZ4VlO/aa7tN7nuDCPa+hZQTtKffAWnjBTiZTRAfmN8lXcpRKc16AY3HISdz7S8Qae7Gxh
2NcEOLWXazj8ncBEBb5Qhd1X45ZfAYtpDzJ4c4Es2ovj1XCAwvofeG5yVNHNw8ekaCm1aZydcfxc
Wit9ARHZvyuNr3lDsTlaMPKpp4K0NqxTfGEH1PW2PRYrSuWY2XA5SdKsqXeHofVhq4lOPz8T67ON
91LB9hJO9xgyT9DWDQfgQT6nx+GVnoth48TuGcl7r0lDybs2+iT+kmZ2ZJrbHD6HgY2G/POZPWUE
axLpTc+i5I9IJu+9oWcR4rjOuV13uj7f9BnluYJnbugTsw+16t7/gUPJPLT7RL+XbFP5tF1TMLXl
dbO3x93pQZv1OvZ0FV/DOubsK/KwJFCXgxwnOwYJ9BA7dOTPTnbpSM0Z9DEIy4vZ7q8/N8G7LoH7
fpOOC9bU9AQ9RdPlJTS6vyF+Xj9k44l6IHqH+g9NVnqRlcsSS1CDg73+49tP2KYCn0m5XTR3Ig6v
nNslsRJFURYtVpxzHpnI80mIeZpWLfCtMh5U7QE80UKJK/E9uRpaBo5WXk1xEt1OpaTFnPiV0YVW
KvbhBojtAPp8BPt2ZPaF82ljrh+9+wCS8q+v6Jzcw13CdHBh9en0iGAzPUV8DEGZOyuATCavimYu
5z+nimjQIwGZSmPKldOpc+77zmV70hbQigFr+Tn38+bqcaeyb2JzOSsCX66aM2UTDU1Rzdw50VUu
nBC0tURuMbpRvhQZSIbN+dfZ+hdNR9FG6rAlcyyoJgHRb89VYu9SrNHd/te+fpEoDkcQxX1Axr4O
Y1j/a0Q94ojC2l6R0HeUQ1W65SWTcFo2hHLTf8L6LaSOeuxyUgZ5cyRbaOIueCXikrkO7lUuspjE
emJzit7GtXpRXVZ0rEcaxZ9I/6qYSB8iwBpS8HfcGB/TY+93/c6mmElvIsGxeb04JO8xdBH8YHxT
765tYIlAE7dDrkKBdv/Yr+7aZcIcWuUAtBQA2rR6nRhXosPSiEQ6gbozV8je6WfYZPAIWPp6M2Rr
qfHHaruNpwy0DBvgM7ZZD3h+98LQS16HuN9if10guw06mYwtsoen2pYYqnMpuqPobegyv6InUyjd
jTmnXI+emIMSzBUVqBuXfpYlJOpMVKh2YZaCQa/LI/BUQZGjozDopXTEu2SNqjMs1ooa9K0ge/zT
zzUvxfAEKd3L4CuTfjf9HQEuvEY6Xj8wTK7ab+E9LLxoFsf+/Q91q2m4B+8rNijf9xu0KCm7VeC0
7kKobO2vhgK/9FBngJvemlC6RaprMm12Cy5azFNKPYDCAy+TNge5EaxpU7o/mf++tX2sSAO1BIwp
GvuAd+57hzBYsXbrRPi2NY8QEnyzWv8aLL7LxSbWNpsJ9+MNedaiAWlf+IdqQ2HZEMf7660I1jHW
ctsq/QvyaBWGGdOaNsZW4M+OZe/+D7FuNJDfDRBag/cm87dG268p6SJbl8MzWqtNAnq/6lHeyTKR
nTCo7xR+7SkMJukV0p/+prYIf3vBeq3ArGSWqQGXenrT0qDYcNcvFzU+Jy/2j+5VMJG1aTIOmm6y
1wqczpKzTUVpnUN2dizzpVkaYCjTq+xM7tpBMwIV+FqOaImSF5HalfDEWUAw65Rhheush/6+Ddqp
UW+byHuY6OcjBgzLbXsIgo7aamuR3OLh+BieKZ9g+TXv4ug/RN0uvFxFCG6Cb8x1sfJLhHpe2U61
wyQwwKhud2oA18KMl4lapDeJNEEzdUkLhr6lct0lxzhX/S2Sofc6pqGNQ+xtB5HvgFXQQXSKoCx5
xcXPYNLJcvfgWu+0pl5lRQMsGn9XvVVcd/baxX80ECWihj93lw9wRiiwk44gZd0++yjQyEr/SOhY
ExZ9CqqVW00y6uYXJP2nCklPEPiW7hvPvwtn170XrvyYrmzcdylT8te8ZTqHNdd3Tc1nU2ucS5w3
DyNpwLZtg5iiNDqmV8xAnDNUrl+fahUuTYsVeBuNliSTHQwjeebfFdWTJdKybWQ589czmRFF5Joy
8gy96tJb81/zk396gXmag0tkw4UtEe+reOTT95PB+olqP8crmFjzlF5ZWG9iC6XZm76g7nGB8xuc
G3oHlM0UizRqZZLJvtOkS4ho/mGUwmS41+FNctWoSy1r01l+B69np6LkCDZM2iSc0T/BHDcUs6zl
Qc7E7qofHcqVRu6lcrq5PMmnn7+z9I3YFGlg2bxjicUY3AmHjU6tcenkqj/AtD8MxkiObDgi7R0g
dNM85McF1+5+kW13WOSJQqVqovycB2qgEDKAgDr5ZcbVr0Qlon27AJvlLX8oFow1eHlkpqRZf5Qe
9RE9RzpmkrgZXU6cOYnsDwfgfdZLka9/akPILITBPQkhvDiN9Tm0iChzDrnpx++I2j7gA5F3vM2X
OXoPTabva/RlWR8k5nAijYzYgu49PVA3eTryBSid9HIsqc69xxaJYCedNeCFNuPnC1ZRHv4w9lkC
ynAfCKwZB9V4UMPWEOWdBap/TFfVM1twmtYpf8PbFfl6VIZ4cYrN8j4+Xxj8e9CQT6u+ZpgeW9me
hE252FdecQcvVc4WiQM7Z35BooMWl8HynuAh2KKpF9MvyyFgTy9FXhAK84aM5B7TsjtllOnnPmBh
pln3PjDpvnFmaA8j/4jXVGhWSXoZWdn2QJskpeNJpXm/ZTVOru/njzvpRl6D81vkq0/DK181ylvK
wICBdpTHriZ6ItVqEYLQlKsfVn/ode0dMgaTBWq7bFsrT+yF8BtIQPKAd3IX4/7Bnd6O2hGO4xKQ
7B4dHJermek4KZodxE2EuSBtVX3d+FMsyVrogVmOb+Z5qL7pPJ4zO33BcaaczNlyjXOKKqB4XtHs
JTAQAR/CYkgjiErv+n2CxqYjQkABZ55nRc7tO/nOKV+mXvrniV3UzUQqVqEnjshN0Y3rvkrmvxrb
Mc10UGXjXsDbqODHdb7Kq/1DgpYYYgTgtca1NLI3LqEH3h90TDxLicUNRHtc/8MSCWUjbe7NCK66
7eVL8akpZ0ThQIOsO+dVADqeUBStGVzEYC8YeF7XQs4QmC6UwsXT3JWZrji1oji+4hQpoH3kzz5k
n++TNpdFGo3mu3+h3oyFyGIDA3wNbncUpCoyeo7Vtu+gXoLCBF81QfsqvNoazIT4eDVB53ol9pHa
9cFpVnoqgZppfTuEboQigNwoXqUVybGoyvnhd5Xe6vCOSN9/hnWveIN6co6mOVMIPipMzbUVIyea
rm9nnHoykSqwnVZhcMKqJbgXQ+oX4eR/NJOiSLhbWl+vzm56P9AQ90rzkRJcn9PuhsScNZ6hJ+A3
2anQUZigRGVM4Ec6qjV8whwJ3nMFcpbYweQ/W6etUF6sSeJXzPOWF0AhOxULNfegYXCSAExfycXs
e+JDFvwFsonH5cIWcaao1sz/eIld3zhUGeQV2/UfJE1kJJrmibLxiHhRJ8R2XErXKMHTeHKfFxXb
tsw6X2KvWZog8RypWINuYHzEjZ9JwMnN435TYtJfjNtricfaL3D8owWRGhHC50mXYOqBR9QPcoEK
K5f2Sj//Vb0lPYIRyL0ak7asWDljppLMg+3SSDPx1wUkvd6KvQDBaRbZt0YPdN7tZ101ETbPAHT9
pJx9TL/M7+HWfV3l+8r/GBE/5rg6zFk0P1JchoQ0RJE2VPoxlVT4wIc508iT1zt1/upeq0O2b5d4
vFqZQhrweZXsseDu99wG93XWTFfg7tawexz7BCyNfmCYLGJ+m24US46yAwpRHjZ0EZaIV7L/ATGz
kMPC3AVJRpi0Q4XSowDSm6F9gb4scconCjwPtRGnuMAjTRi2rhTuLPbzkCYIxoeCzrxtzufVU5iq
3WICB6eOEMyQjHPBxDlSy3LNycD7+l2UgWer64CH4vrhSqy62CoLy7NX0aGlSI/aDk5hrgDCHcQk
Zr6al4BLLs5dRH4DoJ6IrEDekZcKw+aSjaCkIqHcn9ppuUhLLmu0gnmtejFA51utNU4X9xW15mA8
FUl8Xb//uJmQhHoeIeMA/rdryHLeHF/CQij7t0sIPQiJ+zzBopvKYLAewar+T9ItjskY9mhje7/9
NkXWgyziSXFZfzCZ9pHSw+e3lfMkoV+CTqJSyR20Z5DcJuiX2TyElG9H6QoxudPY2Xqtx1sJg/KH
LXcYJGGIWkeh1UMfD5rBdCp7Eww21EhSTY6tHKFzk8vrSqUgQs6e6WakcLPB65goSTl3hUR304dO
W/97LaRJF+5F0wKY7VLZ3neBX1tEYsS6cdQOJSPC4eb5r0y1paIGzyZatXe3VohA/oZ9XD4C2Lz2
EAJExr1Wawz+LRLt6xI1OtVd1nPZfuwX6l8na2rPil+xw/08ho+nv3eFWoJHTe+a2BNM55GDf1zo
Fz/EQmMWMh/iTs0ZBe/hNVqLslgKerHzpNRdajih6ScQbWPgXbwjUoy/3jET8q7shiBIAhE7D4dQ
2VZAnmhATiRahf5iitWpsofQqOPS8anUdzQhl/Zavmchdq5tVAct59PF4BYc8l7iwd0KKvBpO3ux
Tabec1PIKL/Z2XoFi047I+BayyoqWrbalycobJfnbqbsvUGcQ12wkUirmtQUk2sete0nXTQvXCPO
BvhiSXl44Zaau42iGCWWnCjNMZctQICJK0ygyBwHhYlB4VKeqsf8x3rXYww6x/VAIq/9jY2sBWk4
oilNdweEXJgwfajRfG6lkhnIb5XvInhEWVOesrJD2ya5tiH7XdLO1SEL5pCcWj+ggiRgX6wnaiwq
iDFoDNOl/bgDeRc39cY/CQC8p6FVT8Wa1p24g9crsNYx1DaIzPRob7M+irzNYRG8hwTG/GCkWqR5
Cf6LgYY1oeniZ4lGhZb8VjhsgNh81GLeVSiG1LWtlQy2TVLqFO3h5ZXW059zXudlO+VKSutV4oC+
pi4/KR8TFqqn69ssZjLo6NzScR7HL9lDDvlXWFmi9P2eN+avNcA2HwecaT0nrBqSNXlC/vJ8ummR
glRFxQivaWc9IOKlRmhwZtpXxSN7WoOKpvOJsIBqBKBuLrnhLfmRRRwNhTI9kZO9Ep46yo9awy4A
88XbFD2bsVZGqQU/UCw0v2Om165qsFsxlXjfwXVwqWBPSMiJtSuZE6lCuXgXlFF6YTmRf5/baLD0
uDkXE4SF+tglR9AFsg/Gisz1rLz7xpumFkFQ1o5zZfZcHEdwVGOgYv35vaXtro2h4RoWYZ0Msz7M
cj1wVVw5tx1DyOzXlmn2SfaEN1qssRYXeFONkND5ekJ8teVQHZzvqIk+8tQGo2JfRsGWQULGw62w
UACZiaIEQPyTid1DkSWy7cE6llecsfpeM3sidKtkuiFNr+jMo9bv+QBl9YKrXlIMSQjRaLHremny
+uxHmaTv4Gi9ydlMkwBgHQ7c52DvJK7b6peB5R69H0fhhtD1zqm0olHN0k0DR7qJwug+M67OnaiA
vzG/Kkzsgrz9sw9yfNgFkVbWIfVH4MrhyhPmRvDxAu0nd96vBW+MydtxpVLqfUetFyHkh1og3gQ7
s8lUR4VHC8iFazk7F4Evsl8AKRpX3BvHI+9oH6QNabQUeahnaqyqwHjW4eHY0ROZZV4DDHw/YkHM
UxZGoY7ziDbMbUEgrN/i868ljBy00y8AGmUZ3OSS3l5VFswrYcfHS99hCqTylrcVto2k8whgf6Jp
TPUNkNJqCu9Vzg+V3bdLC/BAaibxpgB20ES33pHr2FbJeh4BgV6+eH8SCh9ECUQ4F6thGB6xKkpy
I+LHqHFXs+5UmQkHXw85sst78hmIM/U4LHpIJD03RDGhs57oGmtKPQ93qVmNuz4j0vCPu3XQuS0F
gC/Q23c7c11Ve9RIBTyUkaBVLu2Zx1uL6jodxX8Plv9ooJ5CUpCoJXwc+pJY8+6Iasd0umDN6i8H
wc1iW+ud+o+6i1G4+zmq/3DC7O/wseLm4iEdl8FrMiStEPe4bcpcwcX7byf70gFa0U+qNXcnXjbd
3JfxBgLnOZH0a3wgCGfWN25Csy4fsEIfkC97QgkYfNXDdhDQYOlyddaX0V9vSLsr/NxIDqj28J8D
E7XglX8eR3fsrY/lykGDPG0C5BxarzFS7ysq/2CUZujRc+AkQh3I34gak4pOo63UfO9v8E3Ydvwi
Ut0e2SJoqRCW2LmnOwD0QSlFG9GwpncYDCg44c7gAqUG2bwKBG5Uno43utzxUM2rwCJkldXUin5c
jd4YktZbCWocVjkYjYE9n7agUbgnea9p7+W4J5uEakAZfQGFXOw8wOicFauPp8LOht2f+dF8wHqp
VO41mGMjRO2Da/cveolmQPgZZbMW1X2xBsTjqtnDWue903LtLjQRIseiR4frG9IBXDgtulj4M3qy
IrktjxXpaCSzHWfUaU9FTmHjPsKsgx0hJkgKSchnpiUxg4EdtP6IRakkFCP6QxPOOddxqFYAlWnh
sajtjAm/CTs+tbw2G4Iqk0qkdAGIYw4xNn+ioP9fnK3H0W9t4d+x6S3BNwmWk5fwUEOcEjH/UpTz
MF5Q3UyfM7YOoZphyK37xnf2ByIGyTN9WSmtU0uYr5LiXLx/SQ6MKa9pQcl60CDNwDzQk/6x2wcW
ilpyhRfwLe6Au3x3XJEByfdYFUv9OWlPqBSdl4tV4J//59XxebraNgp6ugBNAA4AouCzE8T86i7G
4BMRX393Al4qcyrJL92FHNAWKTAfx7SK/MTt66JssJnKdT1h1JLSpQUE+9+WPNC5IhCb2rCUvj87
MlsQqx8IG+q+yVjXpFGlmTrvKaJMBM1j/tZ3EuaGc1Fy59snwyUCXfjC9TO0erzuWopiDQQy2+UY
BvHehtE9tx2+e9TvrFxyiK3d36CZoIHxNcaADC8yswwTNTuNvh1M+hnqP52Fg4re3WunqO1YsSPF
kA4RKA7PDpiVn5qOv1yl7sq3jct33QFZgkWDSQIAG65y1tjFEJu3Qj6/gUOPqmZiEgNiagMaDSgJ
GPKoE0A3FRQBS98VM9AwD/UW9ARoyYO1145YGHhdh37g3MoNkT4r8WQEz4GUImyQFcD2Gyu5JRCj
OLNn5iLbs4g6oqyOjSjKyYx1g64kusXmG5ELmJVjUy9UfneyN/iGXlp3bVu3AI3o86y6yIAGvsYJ
fjFHEnww1utsxy39JDgltLIyusH9Xu+YLvtQviJ6wO8u/EEfwkAjZ0VpC4hYasoBzPYj9z/lsXfD
kknYAcFGOmBYvF9EAx2ESlJQwvb/V0CtTQoho3adoRdEtdVMfze4W1jl3+ulR8ypmP0xT77b8lVW
s/stLn1BM/Q648BLUO+V6BHhlxQyTUTx/lonPboptk9DAr4VDv53ifA0s/8FPOmX9JZaYze7cOSA
FhIGfL/bLmN0fTvSv++h+bRaTpigUtS5FojVuelpH1fIiw36aDDnJkE8tp79rfGZOBir7Z/jtaxF
uaCHSVDamA1dgiSysgdaU2NEE2y4B537X37gAdkDagEMAV2IgjjSLM/Yc9JwlQC4XtRZj6EYKcP0
OrAjEZE3yoXxVIYbMWFFj+xfcSAdyk1CmNgJ26uvCL8PlnP6pQJ9jLjjn84+r3LEslaqZ6MxQJT6
GUGYKKKDynxlU6TDADa6Am97fTqDG6qyYSWCJUMb9vMcJ2g4nJNFK8BqJdipPCa50lrnq2dlIQ4w
73AT1Ja39/fO8XwJyUV1rcYpM9BzIZDSz+wRv0DXJrrnyZw7F4xVKaVVnmXE4Rm8jBpNo5967QN+
CHWLy2SVrNu1kCyRbMD7a2KFxwBA2QZdk0SBkWngbBKe+Y+TYC4CwF4zGvdMT+bbWPsELKyWGiWj
U2h0ZItQj2CNjXNmyyYWvHrllR0kK4nM2rAP2l9U/Jd5norXb2BRrYg7EfrSxYhmMd3Vn0VnIkCg
IXHm9WofE/0rti27T1zdlKTBHTvlALpTtM4NEs3wWQHXLIAMiDHORDSfBRVoBHnTQGX7WJu88/AV
s9q9LSGQIa1ClUxYI3qqK1tzckUfcNOJCvbRQjOAw0VAAqdik9klAt9ZYu93Jja4A3aSgsoJvRBs
f1dn2siVbJMKWCBvhmw9EmlTUhDNSlCRRumEMqb6qloU+aXDwphTEDrZlrYGqMcfodL2xV30ZX1Z
oQzdHyLpQlbu87j3eW9W5T5SK2EC69WJNr/vTt88s/QDoEwKjkZzoULrSKGAjnAb6H86Y2YajFgW
O7/Zu9ny85i9OzeTFlz4bkRmKCoeJp0j5+3In/pe6vNDAFT/BG0VF+YfoPi2uLSyjDzug/sRGuE7
s5iG4E6seJoNzbee0dXnmfSvVITMlif8KnuyL6fWz75+5T25VL0IiXSM4bEkwB0wBsPadJeAoF81
3DNqwMhTnQrkPVIdNDLLTb3g2ijNdMwdqOyHv7NlqV1bVRpmT/LiLDihJQ9n90CZ1+NPgQWIB7fj
VXakSpzpg6wpnrk6ahfvwrAu/lKbUIi7NlOc36CABMoBqv+HfHnWEI2li5o6UBgjjxzhR51jIPLS
EOhqKQiuQYnXBZf5s8bv+6I9VFgyvaSm9c3rdStTSpCw+jDXwE4n6iTOUt/CcOUJzJNTYorLVFDv
zMPoOcdPvut6FhpY4WbU2SdFNEFzvOKA/9AWM27s3O9/5xq6cKv1zTDcRSkDZ3FiC6XglA6HDYRt
74N1SBm2a4lBqimc4HSSWeelM2H0ngZNFLR8WgWduljXlq62XYW7wiRIjfRW23ZDUZysGSN+V9rE
jXbFtTB6O6HS2pxsk4FZX/ATemb/bm3zgi9PvEXL9fSV3FcLtU5wcZXTSR/NYg5kCRcufRj1RgWQ
rw2ktWjvSO/eSOQwc3cByemgjyYVl9HSMIjx4nZXQd+ntc2Rf8KlyfSErTxxYBlIqQZU1tviadIQ
dYvlkxaKfnmj6Yj5Tpj9u1SYRs5RWoX3t2KBbJRtqX862xrW3N/UWmWk3hlQ13GIdAVn9e0OiURl
usSInWtUA9m2WmOusj50C/pbjJW9yTafGmgej47Uecj8Uxa+mYmK/Sx2yD4AH9q/04/65kwuffQT
1/joiM8zUPK+JoQtp3GdN4Ednt6VvHXsEky47lICOp1ro6xgPhfMW9I6gDq7LMqjWNt+UPdzih05
rkgv2gW0milIk2kGh1HGpHFLI5GPXFXhI628sYO2v0w6+6xnkYsHc15xaE5Bp/1ydiQA06CTwWyE
dKOct1/pMXOnV2AtvHQJMIg9AqPPmefTYlRCRPOSv/NGkZm2/XX8kV3butjdySUVro4YeLennsnG
yEpq0w18sSEpbRN1aq3fqX/xDrl/4ZCwrYxDlqnaZrHSX1+vjq5ivsO5WpbDv9HnsrRTkHFYFivv
WO8XrPuaDgRalom6jWC9waztxxm2Anz/cBeJRyT5M7vpAOw2VcPQB777RxoVp+/IpYhwnEAtef7p
FSmieKo645xekKxgo7hEGoXJepP4tI0XvU0KwvWCyGm17qvCnjj79goUPR/BTvPzu7wjjaXcMfYG
VTvSL33+pQx1iJGQJcDn9wjqEPUv5e/ayJvsRpAaaKE5UA0+fFWWwbZgpQPap6DfLjt28AxKROoj
a76FF/KvLTGuVk0tRnOueL72kmjAkHNcORB/3sP4NVBFmTko7ClH4/CaJBemoWqhe8usSuysYEHg
oR7D3IJ7hFj0O7a+MZcuQyYQcqfaA6PdfO0kPe9m8ZnKsz5zp2VDLX5k4gzWsOzMTyPyzCySwUZs
zc+lGTFJAw70S0XpQuvSoTrnRTr3paqSiXd+uDCWuA1YKne8xZweFDeUA34x+esk78c3TpuMiPDn
3mvyX2zdHmh5+SbOuEHEt+9CYsbg0g1jJNSb7t227XtcRE3kTyo4qAD/4uiZ2kZc20CtQU+t42wn
SUjEtsmqZeECirSbO+sHzHIsxN/qUcFh9vSrqTAVemyyD6QPhH+7buGX1O4pOOTdYZBjryyI+vpY
yJGdT+9QYj/A719991fCmC8HZL/XZ0URWvfjkHv7SAVv25GN2P1qRxpKiIgN+A7FJTOtZB2xA5Y6
Eit01oTyzAqa/OolsR36lWCLilQnQ+ZU6apOXcdhdQjqXcd2+msODygQAPNie95nGMXqCUF34tM+
2R9UV4iqzyLZm3d3Odt1kcoxkvWsaXhDEjvl4yL3LktV2GhTgb8awnwV5pRp8JgzT3i3MSDEd+yP
aGhOQAD9lJ4mVDr5aDns9YVFNIJfpn8z/YPCS7IrQvxadq+08cT9/FDk91WH2NVbgkmOuziRLET5
GfgQzWZICghRzCtleXbsw5I8edTI6TVf/3HwY+E10DSAWO+93JlTxMCzT1Nbw1kbtWwMZ30ktWnL
XfblV+TnS+yYMUYFIKSN9kXYoz0fquX6uOzJxGMILfTSYfF1EBBlJgEjzKvnzW8cJwUSv+WHkjZy
PSmcqRkJ9xnZ7THMf8Edw+ywuCiQSjv491hdq6lKJSW3e91SgeaPoYF7hFHyMQ7z+TNKjBPWugx1
OD65PL0ekHr/tNzTWdkj28dJ7tFabfJtDMXllIEwBDuqo0aPaeYhJWWONz2K2a4VBW8nIxcuxrPT
yT2RBsZigob0uauFH3rCfS+JTWt56BPVuMlf/TPdl4B51yLEtW/DR4n8zEL8ciiSn96OzrnAydcV
U465lTxYIZvFQnagjb8gJmSfUoTFXLWRVZxG+TsOBEKHqO+NkWLvxI/oAIPDwSvPR30ACYyMuT57
4DEkrv4ZGXXn3YdviiUK70K3bGkTsxZ1YeJ5G4JrxehicLOVy/x8s3ujOuYgc0mClYAPiVnjnmOy
ZIxyPSWTzdO6IR8qr2ovBjRh7iDR2XUAQe7yJnCDGYvKT9QELpSx95GEwdiWoVtgXQ2l58gq2tJl
r5jr+opvzslUv8JFSxq7E3BZCAEmYCWlb1c66z6NWy+DJlDSxuFbUXMif9RDJoOYHoJzZddtEBWL
FYrYmUe+W3Ko3l0GWpf0OLbQhpwtodgUXbyRI47gtPts1+MW1/u8eY0WSIY5O+iN1su+7vkSb9Hf
h1i1r6yBsaXuol67W9MeVPViVYqTPCJfcpYhUTi8GiB26wJNuLKQJndeMoElQ/Ij9NrvYn77lE/4
/6Vio7yy+TX5VChTQUo0+l9uYzoo8LqcJu7q3k1b1BwRIE9GqhbCqhC1/RmW7Dl8hkhyeq0ddys3
IiMC85YD/Qu1SI3EQqO6krwUuw2+AxzfISeHmrXjC01hhSqCMQ8azlHGoJKgKfVcieYSYWo2ZwSi
Gx5fBGvdOXJxeDSEGPOSlTvVyOsEaADTxPfVnBXmNhR6oHGXLxHg+u/s6MUPEEsC9FwJx8/IDUCs
0nIIEHa1YVA29X9icSfSdDY4JAOqsiGOsnkktOg4V2TY0IAI5OVJ8H8AL0pLIKV/spZkODuR9qyv
Fqno4y03UyupPfBu6+c5PchIrGd1HAm+R8iGY0PMVzhx+RlBSnuwHZFw40QLz5BkIje0wvyrGLI/
r5caTF22WKMXkTB/d/AqXm8e8qSZyuGdwCiTSrklL2Nt8v3lxDPruf7oXhssXxHLX3lbPnL7EvqI
et9IM4blBId4uupgb5HG0TZ5VqT5RmrvOsuKg4MdM+ZTr9+Wa9BVlJRNojcfWfRbo2IAvh9n4Z6h
eJ2yWfty42EBTCljvYnhFnqzWKO0yXOkWQoWEBrlc1JXpwHkjNtPTfdH9PJSWGzczUkiYIUMKs4J
ITAhIPGtb1Gi8gerdWi0iIfKxEKaUsq9OcN7loPsvaV1q9bzuj9V3JVRiO2bNELmUqn1XuWB05u7
D+ChV4FrHDrtUVRj72hKqjmtM9Nru/+RG1oUPNaHOkbACTYu92b+/OSgniP35IlQNNutQjjrltBy
YtR3A13Oj+D8zNUTZMZkQRZyDaTDi6V+FzgvamxcVzjKVMwrS/AJ70W17LveFY7pTaCWOd5Li9i3
MALooD7l6u8jGa6xAOiKLr1L4FrMpfMUJ3akLk4wGHT2jG1jsA7nXFYvF/pcgQhxfrxN7Gpb4h01
fBm5dyTXyYNQ9/o6Q/VNHLJLC1zyVwhd2seMT7OLAtqfFTmExb5tWhfUcn4oQl6yebsPECHie5YY
NvjkhZDNkcNTj675wAX4CEl1W2c1fPUeTAujUtfRvQu7LnUs1jRvPKA5T14Df2iWPT4aOCmAX+Jf
cctODmwARVIVz9CTuJ3aECQDRwEaDH+/fl7pNf25mdaauA4/+n8cjSf82LuYAj+8PCSQS5ym3TYA
5XE8Tz2cfnVA0Y5Kz9ONKNuIeQwj3wIEqf6Fs8dsIhvcn8J8JNJXI2YeTA9bK+kS9E08vk/73L3K
J9gET1u3FJNyZ4coAFVJkQkSepuuGShLXw/LSSWAWOqYSp99x1dI92mJmkp1/lqRBBlpwUcBrlWq
SrjspF31Jp5C34qcu2TTMumwixA0oO9o/0547mJGcBLGyk5caZhsRy9NibjJaU2/sMK1/SZ5dt+m
DSYdW6n66Cev0woWBFDnbkqY26gto4BCMpOP+dVdJ9tGFG3MGi2w749t45RUq/Ck6bY5ND9f7LWE
SQchGjhroNhD5BXqM6AajiOLJa8WhvzAAicsoMl72IirnGk3EFvSJaM+fH+PB24cGUH/XBeoO0S3
Vq28XpIf+msdi4QkNK075fEOAOhnADGXcWNPPz+nHBvslqDLymwiWt0UyvxfUV6lZ5yQx1GOSM5T
zNCnK0QGAwT9DSAiz3rI4rkkZkuLLtCBC5ec7M5djO9w0NsSYiQyB78APvRcSv424BfLSMLAf7+m
zuJ48wnfBHxJaAM3pnNhK+NrOqV7MUow6GwpYdrCs43ReIWCIYs3H+wgqF4sqEWMeGUmex/Y9dsL
EuKJV4sn6xGaCLVbp83UvVhCIqGjmDX5PFNYF1/G2gJpkagDwgVEf81xf05+xTICQg7wGw8/sLKC
9w7AO1S8Y4cc+4HQBDcILal18T0qmCWdKpfXSA7aSUTjCC/fl8SKuRpvcWE+YpBx36pG6N6751Zr
UVKXBqsW3J625TXp+GAZ0ox7cO7KDDVIBAz0WRmVfBuyOvhUIwo5rShLtyyqhcyKeZ04zUklzmR3
XfDr6m3SpibCcIskAemdKqm7wZtbGF1FbyXhF6F+XdNOlu0e0v1TmKIUuUpuiiLh8SCJp7EV9wI2
cCyxvBHekkauh5jyHWTkHMghSaIhSQgmK9IHAhKjEaetCiILwO7lA657xC2ytkVLIQxtNwG+XFdX
N6IAli/9DkMFkYcq66y/zA2NiC73rKsUr9Lyge8oJirhv0VpjdO7sBjVhVwxprR3YLxSAcND4fla
v+Med8zQ87P9+dz7t5ei/pyXNc+FYDywBK9/N+wlIh868iGx6oR4l3k75Xl0nFKV/gxTlPWuFQ1i
1QUWFnp/FNSI0+9h9QFBDcFbTKrN7GpIqdqndiby6by1SHHvI29VMqWLFA19QoS94FGtv7kESilW
e3osqBrOmEUkg+y/ym2mafbY8YszUSTZPyHOIyL02xOW3daB2yMkFxhTx5NS2uDO+kAzfm4HSjcl
rTbYrmNUxQ64rCUZOG6fiOf5qF8YrdQLIPFMt57DmoSgnoOpkcAgn/VP49LZCWFnGt/AuChoc1to
OOb/hF55rIJKGGTmLZY92kpFj/uZPuLfZZ5USf+iRf2iTP07NX1Xz0O/ZrDVNGStKi0BXfQMNjy4
FoBoGe4YDbgT17K5YEcfD3KhfzB6LKoGpSBNZYihDg1Z2W71yifdVEZ89cczIww/RzVsZ8DEN0jD
MfV/8RIbYykVm5EhvLgaC39suBfitsWT7RuW0F6145/FGb6rR3ViDUMy/FncmWqHim5Z2B21lNTy
iNU5HTWstsKWkh2IVkry0peroxXyr1Qtrw2hMmM4aioVHuSo/KTq6VM89Fjg4UYqH0N2y4tCSCB3
qUUE42CRPWRMASw28ODWTp+h9suN7C8PwjqsdPmP7Pz0qlZxoBmgPMG5dN+/i1YExKMm4YEFahBk
27OTNy6KJf5FJTGE2opNseMze2nw4BMqP9TwJcD0wAMP1HsMrGuv19VrEEqKWJ62Um/debXbHwPN
Hu21vWDPqsEY/BpS/hrOXb52eDWTeQtBZM/B4V75VXGJWRREoKpF81cActKS/oKncjiHsf12UgwK
aDFAPXcHbtynEYYUOyTYZxbVDg7c3S98rtHt0SF/GH3rR2w89I78NS0P65u8FObb61INZtXinKYR
+mC9VHv03Cv28zDSjShodszQTaXnx8M9/bvOiNTo2+3Cis9toXNMX12V5gAwQ+LeWZU+CRM7hzR0
n/6L+vuKsRwb+e98T6SsTMsUzVnauMrvLmxTCpsbvNkFiCTl1fcDIDkgcETLqIMOniWA11QyMoqe
1LNgWtmI0AV2TEk2SpvQ+k4cbE8B6iCjXg/hTSbWyKBtnQkqFevrcL7cMAa6O23+tZhEIN0SCTtC
btjKSJbCFw5a+ggX75YarWnyxZIYxQIYpdJPyj4pFGwSWBkwuCHYAQBEgiKKHUTVqk1gVrMEK/8v
jZvOEwE4pH0dPxRdXFW5fvmr5juK+du0Ydpl23dkj7WpcWjNUQncmKDVQvVSQDFQ6MpBfTavCKvn
YR2nZXIFbpEEB+BO/yJml/uYK11v8bsSOP7d5P2E+8eXsz25qDesRg/1XMyRxFO6TTLUWisBo28t
KQR1Fd6UDfZDtVi27OTka9D2UAldiaTOj8eW4dnT5yq4O+A8C7m++dFyReNrbOA/NrjqXAf0OUku
bId7sw9DYMKejRpUVb19ZxsLBw+zwigT2PsfgSMqg8ndPWJNy6zojtcjRuJPVLCkRgPRL/5Rsm9l
yw/ldCOjYhvGkgTp0wWVgezsBvgVJMWZl2dRx10AW8LbePcB8cBYWKG6jWTgi4zKk6itI36zKqCA
HQhZKBnZXxQM3ZZlJv1fLOAEkZ//ni/1AXWZlJXBV7SopshOnxMxdKH5NxmuXSpYo7PoSIrMCw0t
TLYu7S+/H8IIZpOh4mlPXqVhY+oPhpryKNmTJbb1Y0PhCIZ6Fp4Jb7XMe5jKPrGE3hmjju69GXAZ
oi2ouShFN6L2AKQZXu/iBYO5aV0+H+YywrPT/JAL4E967PztUggbXdQe+5AslrgDzBmo7yRy3Sbn
cuzIX608gGDECC2QNgSyV84OGAyLtYRME+HI1eSWF4seK61a9gS/2sC/BGop09OgxL6r1RmD0EQP
M/pvih66qFyP+f7fVwDqMTjAuv0GbJOlPwdtxcLfAtPpk8XWact41tzeQLvHNyn0Tgfg6NWVcogA
9OYmsm95jEtZIpytVg/ExMInym6mUDZgDa1Xs+gLAKCRbE/Q0p5FVZTmZVTfcNmxGVxH++bGxID0
NeCqbLj4Ut/o411VYqMrBpm1tNie3YqY1w3gOQT+qLitR1Rl42CclcwfZt/ULxQFZzO9c9D9lwKO
iyvL+LWW+6EG/H/mCyicVKQGFw6UfaF+5wSI+ZrvB9QMPsgR71+hd/d3P7PwLItZkhzvMri6C4gn
CZrLRwvQQn6ko2gTbA5v1gfIUIIzm//NMjDPWqD5x9XLEsF6c6CO7BTS3MAq8wJUR5KJG+EL+VN5
jbhVBORgavGPBGyRHgDZz7/QEUIOe676QuVPb9+ZxQvDBmXlVw9cm0h19nzo4prnncylX6keczn3
ptJTk/02zncHkvu16Bwp3fR44K3m8ybfenvn7U3MP12jzgStMc6LdJ4mPQlN4P4kbuYie2w5iOKI
4NXef9Mvq8GZu0ifStjPrXDS+LRnBqiwp31KBGWAiLl/YWNOConKvOsf3RvEZyMcWl3hhM3C+wJc
94VPc6TMbLd7AsCf/p1Q/E+AW1a4/Ot5/qEWHDyam+HYJzecMcEVnRJohSfYIOsWrfzT7k84CbnH
nWtHvBuKflc+WgLTTzSIPaoi7IVM1O8F98F5gW1gYz0gLlrPuT1YFRkxPDscCP2YBDZWYfImDc6u
aJzHgsPyyf+vwy+PJl4WhcOSed67/Qg0Aq3MlK6MrKzaJSSOi7t7FlYaP2zmq/Iq/8cKmGateUJr
HNxGCB/UcGEymSFE7GIZlsJ0m015kqAQh2b7oRH0NZenFErVDbOkB+3tytzZqZkDs6Vbgr6i1xnc
o0pMuM21sWnhTVekgiXcXj0g1tl77NDifLUZkEPYarK7X79jj14JNm3T5RBr3fU3ZisHn6YEkGHg
pdlCg+d+kEf0Iwf75lCms1RpofRroPkxl2mvBjKr+TWt03N0AhyXxsYRUIiDnd5LSRVBBtdey/U4
6/u0IaZtV2m2xEYNfIb9SZKUR6v079VvahyZs7Ll7v5VXzNAwuyKYr3eYSB/UAT7pS+tlKz8uPwY
V8OAwGWJbzv0B3V5/6FvMSjGZw1pDEzCxw6Qrr10Ja6xmz0W1N1FiEZNGkXD0IBXECccwTmANMN9
VDqZZSmX1rlli5oMkt1qr1rN0hL3uyLhbbGjfMRAZm/SYnOMBQ8PGFl4CKSxs7gBsxYL3oAOrCyQ
LSp1dbd7wS5twvaCaojvryJLIAVSFX1WcOUYM+Je/oNv09+gC77fKGPXz//dpwMmTox56XD4CHzh
WPLVay+WmdwZa37ogJo8NEbCmU8S1FUbSS00I5P1ks47kIIZgaZjUqV9cZG8Nxo9Pq5PrKhrD876
haza2YuZqWUgXzp/+CncT2gBqhtFsWhhaga8MhA4nAx1RZnUk7k/VpwnIOy3UFEQtd77HcbAzbIJ
3uDMVEtgUy0nHaYOF+kiQUBuyDGuFwE+4ubd8zAKKr+u4ZAWnzXhnaYTRSuUW6ZbdiURt0NF+xku
QYFj/mkzRP2K/73NYRCcWgAacxABQhArqP1yR5NAEHi5ETZdIw5fqDgx3hxBMLwYqckkI9bOkbej
RfXSctiVgGHJSTZp5vcgOIDWnsm3MG9uAgdtze3YjBTHmEx82vbFPcKm0JdVH183mrWKnl+2rWgf
0aD5RKf9s1nNoDnwN5jEyhwJ3QmzUGtBbw04lJe0BQ76p2qCml3Zipu4YRq0pvDioiCqFRuDs2iw
VSFcWD1wWvhMRar0sK98QT28LE1m0A9SltOogAIwCJF2oHWE0CnklXffeCJw14m+evCgqHvi8mT0
qzMca/AUzcT5PZLl0iDy6WkSVJ5C21XWGOEDqVnq3ftSs0xImWYtDEwyojv5d6IpRjRCo4s79cs6
hrn8xY+2L6wg/0UawW5AxmIDiE2X8AGz6U+9k1j30gY9snRqZnFrGy0JZhMPUS4wD9k1CgjkRsGF
OmtChWYQgf47IpFlDxWh4g+LBHpPOkuI3/hh8M69HACVj4EaZkkgIrZdQe6vDd7tNDY+yKNHqPe6
zETVWcAxC/2V4wW9OF8wxtHgzBDC6ABr0sIjekGuG2P+4JqFMiTz3kJ4kmvVMyaazSc5mo7U6zhT
H1fji44DIpHRcUsNJ8rhKtlSFG/2wT7HrEsxVHB8g9iglwy5d5UriN8kY2B9XsViGKyrObDIw2j9
UuIwZPPO35sxwJtgTWcR4miMmCi2CLfH1V7u93FD8GH/Jp8BZ76drosseRXd3isHaFD8W4nvtYP6
5LBC2/ktS3BQU7FhHJNelB1D25ZffFr/idrdT/JnkacDcWOImCl0i9CRAYEAA43DS862mk+ujwml
DOhe7EQ5EyTNNYjU/UbBjJo5PZmkOau3SE0YG4h8YqXYSo13vPneIIRdn2t0GKZOkpCdRf5OyQ0A
QCsyagwGjIY1HKQcDSLSWJN3jFpZLD49PP3XmGurolrZ1ajR4E0PC+xY/nPqrf0VBqQL7xOJL1Qb
BdMiJ2QUkGHhQvhTz684S4IrEmdVFiAmWaYi4BFhGuKQ91+pv+DJwcFvWDzzlflkvsjNb2abHU73
xgtLj4lAaSkGeQSaQK7ceA5eX64wGEyPK4lQ4D6k8UCHFkNmWuy/e6ko1RJlbLymqzxIr/lRepjj
vln1R7RxHIedRIuub3YE4gGASWXqdAlmWRngX8D+ipWnsq90z3kHb7hawC/hI4vWHa76Xtxp5ti8
bs3blOnEtfY576YdOZSSok7d1V2CPrRlQUvim1gxA72apKRuNgo1Q12loJcZdfnM6rpqeWh4OA8d
VZZUO++lngY6O7g2wQ0ZbbPw/f6Ru5nr46i174ygujwSLKo/oUhLB+/7SwrC7s7Z6rTrA3pRp97z
RZhyYvfkOf8QE5lZ4wsZuJ8/Q960Qgr3MsU1XeEPO0lfn8rJ/1BPljtpZxhRNkgGxWxWZ30x1ZRe
1Msgy9bUfCAxwIi2HERzK2iKWHUzmzJtJIWIUXaxHlhQzQ39ID9wkjuaU2Ps8MWewsyf+Zy0H3qJ
4YwHWCEw8c+lbw+ceMEifx9C46GXkFhz1Q8BXPOx2Fx5gX9q4GYtAC+SNNie3RWJL4d0Cq2gQ/lX
KLKJR0785/Hxa2iV0SY02Rxz8/lyW/rcEDA51i+mr3a4nKS81bJJ/1iTKrW+vzeeLd9TFyFE74rE
gTwUtu3NyoWb/vzeFD+Dg1Y/6uE/Vl+nuCJ0h0/0OCNhFVKDRXlMR0XSsbLt7VrPBTjoy9Vs40RX
sk5s5PKQi3yLvUZqw67mNooIAGVdb8B7Bs1OMa7bf/CzTnHZ5cn5+coQMWiWAcmIp4fybr8n5pBe
mfPMaG16xE/AmbKKneXByHc8xWASwcgoUaUe6czmDfJ0saERWeqeE5N0lSbTsEdveF46j6SFiQtJ
29cR/T19C+ffLPZq22iYr9CU9GvkRAd/BwYRPWp/4nAC7pkZMY7R01E8f/24spoy6Y+XRBUzY5al
jcQt6B4aQxcMaddLUsB4cOhPjq6DkVn9nN3dyt90mkNtGOtbZgC7ca74Y2pAf4UGmVttHj5HtPL0
ey/VwaumihByICUG4clDjX62PUlvuCxVZQPSAh3KRkfJfxSUIuKi3MNHT78GZeQzYKOntRt5j+HU
bR7gaqpZv47MPaEd0r8DKbFp29ECxVKXBpcVALaG3eZQ+STYOlSf52sMTfVFXhKWAHy8NzK1J7Pe
6dE4vOfmMwhDt5UI/SMXGeeAJF3tlzd44DzJMCmnNZcYJGGcGDCurCD1WXnHlWWpvRJaS72lSbUU
7RV+FIokXQnTbP2t7W2DLU6yUYyVqV6xj2he+LpMwc4Pv2UonpFburXQWeEQJ5xJEvIzjMr61OP8
pppRc8yeJTmcSJTBz1Cg876Z4+knCHYPzUKDZXCkoQ0ebxqSrZEZ9wjUmLw4gIbLiI8U/OM129YH
a+IV0W4REXEz2dLF28OWcd/0HZS/2S5asEkz4+H37OHVQzTxkyOAW6wRCV8SddKqPBRsoMAEMYhO
P6z9v0VGWXPp9y0ebfdmEM88dsMO8u9TcQWzEuGVPc1KvPE3oB1WuJQ8qSUcgFcJDM6/UO0DBAJH
JlHnMBwTyPnPwH7wadhCGSfa1GXGHHZJu+2Jz3EqOoTUFzzIpZNssYlNf2LZEJRWO2mNLev/VP+M
SQ646U8nSdlNbzHC6Sed/ERLNjcDKiPir8IK05rFivcnQV4L84auesWkntu80j1UKCXhWOOHKLh0
ou0m5mxOXdvfYP/qhrHl4cA79ZJeAPVhxslavhLEJ+sPwB8M0Xb//xizXZDH+xlO1EVXuIWIbW/m
xM7nJ/h6+E7YEYKIf0/2+LE8f+xvDuithZg6kTznIu2IGy9nqySkpe6H633Vj45R2sbV+/2AuC0X
p4QQH3elgGaYKKL3Fr4H2CXphUsCydKpQ2W5xGihSBCTqhtFMnHn4zqu+yneipAWLmyZ5rMoCLMl
wH+d+WiIvDpVkN1Y+k1c7Jy651D94qq1cAPPLeTfzFR66mKXY8QoOGW4uGrt3+/Fk1Jxhpg1ODPC
2ipWZY4jg+Vbv389zNf/xofokS5LiSDbZdtEA86qcehS49pQ+HyI1kmvBbd6OQu2NRLR+NgTOzwr
G41hSU5NcMApYZzFrgHLdtzzwErxvpNO4Rc6Ap4nTN0fId/kXogO2RKiXZF8RWmjdjk/ys6/M8MQ
Dk+n23rb9pRtBki6VK23ZpNXNB2OY+5LWmjcROY7zm05zztKvOKAJ/nQ89DQYug0GVEA37qeHpzK
HSGZRJopifiIOBWnTRvhT7rCdKPdSCvoR0B+T6syAnhGMH7q0O96mKpFZ8XV0zYfYhx59A2Jl+w9
GnGRfGced2U528ETr49gYwCZ/XfXaGYXZASm9ASZLuQ9zfYXpmwT5uzhTgiXKg866ZduDjKwuZKL
uqujMekOw1wefGXF389hYImAQL/uR2a96wA1EWOKpyPA0JqGaNaERx7yZe9ynhtXeEp5XpDLzpUC
CJfC1rhMhDWAWFR0HQ5bbyKSB57q+WUBAUWXffDJ9rcWhLWTs4yt3LfBEvA9yNWODTGfyqaukFdV
eSIeeBPCxLYbLp03lmK0seEaQnPxDWVb9SgDcjh4bOKg3BpwlsAPXAa2FC2+PpgXHexI5pNeq3Nr
GoqUdEtP+crTGotbihbpLl5fOl9H7160Feoguu/v/3DaqTfM0FJmi8tsI5xR7mPHqvddgYhQt8C7
aWNp4DmSmAiasdgvUxyJgAjc/fPwGN1V7gT+wO1ouDPU8eFEwedpVLfaoEPbLrgcrPs77qLvX+Bx
NTVd+wdgC9bYaUhM8TGZcA6x/0SRqkneM4SWYGlNFSRr8rmKBEi62+PgFIBjIACvCvZopVN/r01r
4eF+njeea4p7SoaIwDhhiYl3vgFcfKffHFJ/zxfOfbkwH+T2tI3GQxWKheGpvqy+XLK+otzBSHSf
doHgYTpvP7VOKCQ/g/aMlYnaew1hQ/vs4NB2htO4P1qHWJaPE1Jnxr+H10MpcQzi+JRsykt0M43o
odTfpvc8ylmxnTc8cS0bLD8HGkClQxS5wEZe16+ev3a/op1Cfd3xi8Vcg+2/gGrTpZZWzYLm4l7U
NOK9QKlPhwCjT3RYqPoETGEzGlk6zbSbmDNhTxciHmIq5E3oQ7CsVQhWLG69f+CHrLzyGLjWRF7g
oMwZwjFC+f+ldJxpppM/NrljyoMDpL5iUvCiqyCEZY+uFFRE5BRUhNllYxNshqqGPHmoi0rocfmL
kOh6NXD9LYC7jIl0S9NdTz/zyyzShmPWS9FJDrDmA8tGkMDHINO9KANKdIeSElVCetCMwCgs+5uB
34JlcvzKTC9CgE+xRODPpJnTN5bEvAZrWGqJuHawC4uZJBUgZpNQdyy3kmfI6NXZsCZF0vbpmReO
PXv8rV7hgYIzCy7ct6mrMUuQL8pQx4C8W7Oazo+X5yGSobVaQdR4Kk68l2HRM/vyJdMRfryOzlJJ
cBpgeTJiYVyFPC8rQwZXKAAwk7iyuXDOJzD99RLGRXNQqb9hfxB745ABCTfGi73luGPxkGvp8KSM
ig2AfRhnfQW1b1Nc38VBYMMVCDoClKatSfOrb+Lxq58uqgA9AZhf7e6wi+B5R2UC0tk/DH372waG
cvxQWh/LN8EWcdcy6zJJ01TLp4PZtWBzi5VOLK1w3Eay1TXhjauCK4Y043LajHcVTJ5NC+BlA71n
v3tozdKX6ArYFZjn7I9jdYmxRgnvP0HXOLevu/W7QzHfY3Xkq2j7C4bxcSGHR6bZ1AMAUGX6RKJZ
9VjvKB6MSvkhihK3Gbi8Orwo+CNKy4p2IbDGj8LgHL51mBmr3sj3pdYglMcjNul5/jUOm5D2zQCf
qtuc7WSa4CXpb7ijukox5VC7jgFQ8w64dFHRPXhNgC8IC5w6I/LknNLh0yRACdhhVefnhEImVzTa
KBrigbBnQKLy6HiNDO+74EJ8kfRNIl86yeOaPP43Jx9XUJggbP3Dj45W+yq8bM1atE9XWckck+J1
pKh0JjTm1X22TTgoCEpsFe9MuX9a1nCoRKdCPk7K+ayTDrt9m/nxYMHxIpJZGI5gMLEaXPkUsBdQ
x4ee7iW2woC8KLCzjTccelntzmXVSjkrb3sbaN3VRk/RXYNa+d6ufybiF+iV4WYZCyMtN21dgk0Q
eRU5NoggRfi0aLuE9GYQe8VZLRB+xSpif2/EsbqJvJLjsHElAsu1/gp6sgwur847NAXoduqH1KDH
VPuPCHUw49B4rlGDUEBVgnbSqAJWN+9T5vBmKPN5pHfETupxDQz14AdXM4R86eNFNBx4zrL3C+2g
mqQQ103EP5/KmnJiqWSD5ZUQGtCvVEP4eieS+oWmxWCAI1tySNiVp/bD0pW3Au7Hwgm1/niByUUf
Ik0eDUTJGchLNfY4uZYwOB8eWctnQHrGQQFuI/JwTbevD7sxVbthCb0jfhCvRuPKiF6zQ/Ur4elQ
U26dvNCi3bG2ogq0SSBrxFLZGmug7h/IyHiAfIX+HOsmULSOZAg25akul2cikv55niv0tyyl2DyV
jSXsIsSn8gLaMDac8eO5f4Dl6K5x6JAojedpSrJsDGABA4hb6Fs9LDpLfVi2edehKO8Nww2JcH23
j4m9dLYzca5dooyJT4zAL6xAtAwR4bfNeSlBVXDYnMxkRBqVxvS+0inaos2kI+0eFlvLENoj/jTb
IY0i4ZKKwSQafRbQYCbjbLeG87d51yJGec6R7ws6DMJW1+A71Vuy9hOV23Q29orYGr4MzUrjHeBU
0cNNowCmVAXBEmqei7bud5OYkfLZzbowiT9gFBeyS3xY2A6G1Kjbt5f0jl3W87ERmqqK02E0MAzE
iRSo2LbA0nmtbVra/EVkFM5et3K9LqHZzMGdeteGENL0yLXKmVuLGmHwAsksJ4TerRInduQsgTRO
spLpW2YXISxaTS7VJzE91i5XU/fyCvd7OXsDce2bKj0B/+TotVsirfjcn1zpv83ywQhvLqkXLuHl
vQ7ido0kD+Xw8nkEBQW6+PEyPUke2TRwsvDxkOTVkxYsK3/2nJLtdrq1nYPq0NfKFHP6i9lor2qR
l22Z99r+HkqP929xu4pltP0Bs3wGMGb/3E0yEzHuHOrbjQl8As5vu21FQ73GjT/fnMVKP3v5VtP5
TWeTDzzKQSv5qz08P7P5VolTExnERq4J/6BiltpOIGFvjqAYdzpCDKdWsfitj5JqbOPO1ODq29FG
VjRL0GsBW/oQ+MNJO18sZhgcxE7XfjtvN3OvFkXWYc1O4Ed4MwPlqjeotHHFDrZjjhWSOLo7xGoy
XEe86EFQ476lqLdwPzR805XKiBi38Nozvp6Qvo2WQXUFF4dDY+Og2XI9+DZYsRfQEg7ZxCu1O1Fz
lrZRq1GAtrlEfETywTKkO/pCZT+HRBEccUXXU6x/bSQehd/P1smK8R2bCkAwlG2CEte/CcuKRg0n
f9EroMsjS6On4Di52WuRYEJMeydV5+LvTonOgxo8BTbnWUN71JtHmR/hp1kVSt1bztycwjcfL5Em
77Gxp1jm+OuFjirr/b454ckq4I5WeuV7NQuDhoHBJcxt7gPz30vuH7fOKvNPBs56NKQFPaapmp/f
V4+BXPNFZ9fSuMggfaiYiHwfVDdlDWJBnrIoCO+CMXaA2/whUTtrSDUqLZrdaEkJptvw8Mv2U7oZ
KHmdm3jk0UyUYKxhYX7O9UyJL0nS9P9PW5MjF65uVtp4+zIojD+U2swT5xPG7UPGPC9YuMwd5mGt
5wyjPKz9vtouuAisx3QCBGE1ItjpAMAiVa4+JI48l1MQFGjhJhMSXae8FekiAM8OIlLByhwEnoX7
WOk5pS/pxUh1TGQB+/wF+N5cKKgeP4WX3FslmcvPrrB//TWROAlQXR/Lmaj82U/U6U2cUuyapiaN
QcimEYsSOtqI6uTKsIhPhRc9GHr/XJ5JQ5QM7Ubv3jZyo74cdfi03iMic/WAC6Q3HBvDfUYbINTR
bAQ8QOTbODnReKM++w/dFVv/Tcj3G1EZ7C0M+ka41fisBt2J3QFvb5c1TV7Cjef2LuVxbCyPPeD2
wAp7ExZu86u43WOY1H5Hd1Do+TKKvVxxPHTZYsSZQqc32fCU1twTc57AeHnkM2nnTdYzFHa0KfEh
w24nhwf35xkp4xe86M02pH+1/76y7qZoVlU/OUN/fz6P9NfECHSZ6LILdjW9grMB1SzXkKy8ZFxw
iB4jCqgGYKvUMI+i7I3deQH/SfhA+OwqHO6aBe4pOu2IghAcN6/x/cxFSSD2KvONI3ySWZSqRR+Z
lH6pL6IOI+TMCiJthOdTQsjGvK6r4r2kXs3zjC99Kni0UhKoSa+x57Ss6kB07EbkO/XP08u7ssDQ
ml8UksuooFzB6UiKIp6U7Rp0iPVkgbE884Bih4nhbhzWviwiJ+9Y15cWmt4zP7uPASELFJlciOWD
4cl/hzO5K46JoM1hCC0PDbDj7BhWtORwDZcFs0+pY87rS2sPO7nogSLAh60IGU042OcSmp3G8WoN
65GloLeHEOvzqpUBtqPyeiXbZkG03jt2fGBpM3PudUsfnx/QwWVp6k0FMFNJJSs66QKrCX5zE7x7
nzFkCWiRl87Cy91BZOzwpERth0XuBGayjG5S65IJehiJeopG6OgxzreQTF8/IbDCb8O6BxmLzsDR
swh6njbnVONzERmlGaVNDZ7KAcGek2hLqK0el/rZYJeAQO25gvurk1UtfTyvFq5+2d42jgOnlMxV
whXj12/l2+AR4nF9JOHtcwfqH07ltFWZhg2oZ4PPLyLZ26sU9++yQECzdR1xaJUAn8Sk9wnVdoPc
S63RKKpIBrDTCG5vQu5ywJniD3z6kGjHpLI14L4OFV8kUVf7fYQBfuAFT3kLsrscw/H4uUX2jiEU
Q95JYZmIcTTm/K324CiGWvDKbW+u+DWKTeXeUFqjdNT5+xLAjHrIHFJigIKaiBG+hgFPBOwjRQrT
IxTklzqOT4ALx6oc5pM8e1tNKtQmIZUzU6NIPMmOxBjS8q540mvmFJSK2l/qbWFkdB8s5u68paHT
KPRM2t2qFiJrK2YU9QEkr1VZrChXxCo0Mqe+CT6w6A6d/64w0sakP2jVJ4OMOujQ+uVD7LtgboRF
iV82yOJsxRxBG6E43wlzNKIBWKAfRMpx9VIv7ceUy/aFFwXYGo0mhb/iR71IvRy+ddbAUte8BIwE
pf86wV0mHkYBSnwwrz1nex+Htr3CK6/0V5t4OJkqNCa0AE+16UKMM4t24qq6RSrfATViwUHSR/9W
R13eHPbRDAOwvrBJgzT5K64uiyV+42gLwD7XlD7vw8LrQSaMuAmg0LkAkaM/7UPDTLG2fbkqVG6z
Pv8+cVQUbviX5jtqsU3pvR1swisSh9w2ZDRUrfuL3Sy4MiKvH5BfIbmMh/vGJAQqeghZeL5/NnMf
CdxJcU2d66vctuJsF6ttVu9V3D6fM9jtLV7cx4wF4O5r5vORnXXudchZux6dshrCbCsOeh8qOQIL
b3w1+6xpTWW+0YcgAmnPvFlwvxaKNJ0AkQsX9CkQWlqQXGSeKqHOpz4ePmsRN+N3GIb6TopIh1Kw
+uJ3Gungql/EryYSHXG64Q6Kms3mlImyxdVI3qyWC6XZEFp1Y7swjmpyNMCz+oJ/808Wdjtdoqf0
awmWXR/cK3E4hcnG1ydE9eldJirUVRi27hMSbQMu+ergY72wzV6dFBe+Of6Lgd807Nk6byGi1326
fszNrwINY0o7vfI7FC6frFzh1RQeeMREXC2IZ4UDacakRi4Wj5ehue6F7UQFnMz5+jMxyxpvEdLN
4asx+EMqa7cwFFAfcFyhX6ye6qgmcQl9W6TYI1BqETQ1UJCH9kXhYX89WKouHqd+Bc9tlNUPynZZ
Ye7LuxZUtcdS/urcFNHqKmZd2VYp595MoyfXYyXCaXFuLeyXXu5PFge4cU8Lo93c0IL1GJPSjQVt
9V1hj38zKU6ciqieDsOo3NtJ46W9nAmLYlNe66XgxT9V6MYAHuFQdafzOp/BDV2zBTzVJ8a72PcP
v+ncRtcX/jO9ufPDxSrsmp4xc2gyWhjL0ClucmAnf4swEs9aukF1rYrDZc8ZixXyG2U6lVGWuPYZ
3uqe//v+jqx84OSDlVwLuJvPAWj3pq44x7a5sZBbcJmZEuL9iEZ3EKVtz//K7RxaKN2GyTy61i1f
3SBKQKUrvC78njp7kGAD0JwsGkX8C1l5sYbzEQ4ZWeh3Ivoa7PZD6gpkQFspqG97vdtQaP57rp+L
62tfrCED8KwYrM7MaYVNDSZpDSRJbbMpUsEA5FLOjY9Du7tGHXllpiuETOengCBANn3em+q7nPPa
cuSC5HqDNrakAhWMOeuCXGX/HypBUZklzIyv/MzD2vUXv5GDD/2yrkV4Tst2GB3aIUjnpClSjSeR
HB2smbM7HxGuC+JN1QXPpwas2eU029Tb1vwCcczgA9fiE+YXMX7VqkgVu1TmBot+m4kTMT5N705M
cmuBcntpS1wtJIIF/pqffRnPUObEf7znSdsAAv9mkYoAncqvm0MyxI8fdUHjCG9Jb5fPkvL4mXNS
rgoVC+itG+nTYIkh0YnRCNNU9MTPrzA5zibYScSyNnT4X2zY1La/hpnHRjtvTUPT/HVXnNamaz/1
yjiNEh4d5IKS14QJ4DESOycRsVxPDM4FIgE8R6O6ChOiUqvhHyqmpqbB5L+3L6Ly59I6/SgOB63l
mtdEwvqBIGoxdJArgrhVlVv26mxNs3QrqDrWhfj14MC0Z68MuisCAig0HRodMarutARLxmQU8K/n
xIDiOiZpFGSr6BDijuDEygGSkTwknPEFpRZraVKGvvGwIZDpQzrS17cfnx2I2k0r/cayzHhe5V1p
EKK1ZUVaO5AjmvrnylH5PXgGajUi5v9+Mw+GMENISmt9v/Mxc4XfVaEytYz5np4EEnnPECWup+7N
lSdZWuI7UM2ZB7QoK6naRFGGurGEmKQVixTkwuuuV7O4Yg8JBT0WouQl45K/LCFbPCaYI4EgCn5c
UiOu3Ul5Ik/XxLGmY/wv74sDUCKWt8nF8rFpTSBav87/GZgwjPuW7muQOLjr6PmH1j8Aya8h8nJM
gtYjVXtJCoVobJ1a1KWoyz8VaRE0Gj2KVMo9yNjMy7s0tYObbQ95KEXOQsccuz7QIZ5w0BOWhUf7
5UL7v2mXBBJQDAbpKChNxtQOqiYkIWl2/Bva03YFXgCcKbA1TCtpUpFU1rE8LHfADU7Fvpw5fNqT
5CX2dDS7mXD7Na+Z+oUlIIuZ27wl+tphjhjsgxKIdeMFqNy10R3ByvjeK0oXWtyEfz+pRIkH4rMa
JtSLnS3Iihugbuuo+w8Q9+M2NSwG/1uSdII5VLGmkDnUopN91uxND/ihidXXcqR2v/t0f7K1NZMo
TgRV04OY/ockc5rs4+1WN4WpMdhxk+yF/lUxHWjIBORd2b+Cm+xdgk1qjzjFbHNI921SpYVhIgcf
ntB5+NqGhf4oMwKB8pYNI+TE1+jko3owWldSLq7/hcQCFLZtEQlbdHACj809AJFj3gstqpz/lQw6
iJIHVd/NU6/Z8ph+cyvR3mCnVbtEB/SHeI5cdgvrW3/H3qTtvhxrWHfDIOlV2hyZtXhndIsL64n0
Eg99vKWdbKn4a0z+q6i6iVXZyFsiD5P7IGRlcA9ijHlPO0Q1I68nqmSvNjVb4GIA3biU8b7Eflix
qGzpWqtqOwHz4x31UK8jFzSyE219RgZhgqpt3skrh5rEqid3j0PeCY+UYBMKab1xqBjYt1qBgiMB
S3qrhJqd9OcZ2EunpaRhB83I5UYgFhi5Ud7zQ5YVKR9lFwZ5TKv2f6pZ5v20uysmiYtSgJy9h3fm
Ccu0ApLwN+xRWDElCTlkbgbuGzsftohiBQxEyLcsTGC9eRNO94AJP7+QpBICsJ/SzntUyUSbE9XA
8Go7CorJ93fmCikQDWIC3UCbNUrNZOb0E1WzV/CZkHm1rEw+fdB24mDmxTSJsp5Y/4sAmT5GGRUr
Kx82v6WgEKRsfoEX9Q2y2KFwGRSvJc2avCMWKxEYdHtykysjuRMIItnNrH8rVdRFrRQJ+zGtL4x+
0e6UApQ2xSPbWohhcJE1/NtCQydmaRtjvK5++YD9ApKxV20dsR3Nw9foOf4/aOiJSzBQ5GRKO9+p
SJaaEoM6H2OvJ6JioSTqQftj/Y7WgV2E4PBgAtYRaKguXWnl/mvHHNJATKti+NzSgHnTTwGaZWmd
a/v1aT79g9Mbn0kF/LvB8t5vP6KP1nRCAO6bAmMYey+2bpwHGWk/65opoLlcgZZSLdR7Zot3jXOq
JJgFuzUHvdMjCZ0N8gezwoUMdOvlM/Tz7FqyV3Mw7yK57BQYGCxYebTvUGHhUUYT8HvV80YK+DGj
u0LY6i+401cCXXB0EupaQ3PznEOwgIITgl3tu5soBdr56L/rmc63cK18mzWMUVZNltWQ4LDHB8oo
Ghi4xqrOLOJ3emIiWsRNYjypwfs7vdA6FVFfxaV+9iOM8bJWQNHHQEy4k2wrdSMdUceEVM+l80T7
oiJQsRZPkn+Fx1zmfa+J8M6x79r6AE1zTC3X1yv52sXw7n0aYxJnaeJc8lG7AF0IoXjbwWiJLhdn
o0oyXLwsNKCuL/luQhc0x+9Fq1ca1GuaTnWt0i0Nn91SfTR0gLDV2y9Ssd+4JMQBDaZOos/Aakhu
20F034CK3vys+GYXFF75GlQYISD2BbYzOH1KMJYwlW+R8e57d4Z7nX95iuJ/Q6MThV56TI+3gZQg
Bl4YfkOxa9UjmZrV7h85HOo/LWAB1yepYbgQcniS3wXbShbcG2tNK4iKnpdtB9xYpV4IfnikgYrF
qqJLgye7/SIpnJL6eaExrmmAENe7z+G4jyhJ+InNsCNvbokcewEVEg9moq7YtPmn/w9nli2Q4CfB
6BB6q+HKhA24/3YEs8ilvUbTwnrOjGYIsjzcQW5SDNs+jdYpZeoXDs2XKlJ+Dafh/S6Abi6gMq1q
GAvR1Mkj6qU3zU4u2U4BSMDWsCs/8/e39GQT74gKcNq4CgWFejtMiArPC1NSn0YBVUZm9eu/yi4/
b67pknuKzJiYBHC6Gk1OPUH1iyefAx+iE5pLrZh/gj7HPdvSHNVGJcCp4mMv9lSxAcUa9yW9GX1h
TVjNvQRcwtakxxBcVzQ4Kx3ASWQmmkUYwMIAI74xcgqO5YPcdtmv0aMVJTY4P3mef2avdOCJQRxR
H2ETjXlgSnLrnprHX7xeKn9JzJ8gaMg8aU/3ZfGdQrqtzsCS9+dmprmlFf0vGydowJH/qe+0Qnf1
EGIXg9INxNZ0kR1COjcxC8lqGQK8g8fagHPolEOGvYtUs6779FZS6rqI0WEjq1/QobmvxCIMK1v3
sbng6mHKyf7HQ2ChVVWnOZ1UhWG+OgGkEqFYWRl434p3J1YyIKG675wylixUU2XaqWqxzLytEAc7
dCxpK7Se0oxQqTxwkfOq521+di0qydvB13dsuf+TJTDHFJpeA5KtQVmoCuQKBz/It1BJh14ZQ+Di
8UXEy8UpFSTl2xGQvVwsGJ2vqHYHyeqIVXUnbWJPVUPy6dkBw6zWleBhRbTada0LGLPJfNXtTNYJ
KhB2SvfadGtt3bf9dGPXXTDV6htULlKDZyZztLhiGiLkUq962dLf1aINFP8GLy9Qksj33cXKv0WC
zwBsA21NAY0ciAZ+8D9TlUDZn3xKcm08tfdg3V/CWFYSx7nONHFJaYOxCtVV4T3GMHp5yOjOoJaE
/f7ry/SPM6u8pSAUjAlsiQRHcONT3WoIOwO8DBw7d5MWvR7weO8DzJn1inmLG1rpQMNNm/RkbSPa
8bjMqwnYESBGuPQYQFgIJaNhARMNKaxxF3kW73DSkxWqaMmQrp18bYrTEcA8E0zLVL4Rz8jueOJM
cL1DlCpxc0XcLOhDaYRMlnxYwgt94s912QUX1XQRrKRW8JBAGXSnzyNWcE2fMTBPOn0GumK5dOSQ
X1cQvLtsKsSSqbB2zlc2HW99zNguUueH++5bEXzrtVfsmTgVZoHY+F4+yhXWG+5pyrggRCpavVI1
ldYmV6IkRtjt7FGoVuMLh22QBKoErmsM0HdtuEGE9EYkP/iiQ0qksLl2LaArQ85nHO809VtN3gR2
fgslVq4aTGjniG2raV4UApv4kjxnfa956SXOo9bLPUL5ni8BwEe1tXpZHQpK1I1Dyd3leg0M04sz
mj2tPjgw5HxOS6son14S6+yrZ6lUHXzPX2pe0V2gQdRI1aanWsoIMQFpssk0B1slZvBkAna3qbN3
C4z1LP/Dz0qn0TIDhLnFw8gI3ri1PSLmhkLkRU7ABQ3tByKaG8+XZi8E/N4sElS9WAzs359RzN0J
f8VdsMkh3dU+kKTrtEsg/1t0gsCNdG4OXCe/JpHwhcMAJ0GBqZlJeV1DS/8Ud93g4oJILYPy0bz5
hi+eGtY+n/ogpxDxsVi3OWou+S9DoFe6i2dY627bl6N7G+SI/0UvzpSoRajVLQkeRM94aAYVPqxg
pYpJjs7nummjAJ2Fqwc9GqvY0BTposxMR1zzzzhZ8kZtTfDcx4sOw83AKggEJRbto57q3b9wSvFq
AE/mrS55xGhVxO5AW1INgtaZSY3+KabcixPmIEWPJ+Tm+AZB9FGB4a2JHrwi/+KH0p1zZKw8uGT5
RBNgX7pLuppKMYrAaJ5K5I7gV+nRs1BjqqX73RObWlzBlYC32VIFpaWiB4JKU8Q02IUbnIcn4M79
MOU8cQcGge5AjIR07MbLoYuZR21I9ki7mEK1HXmC4dKU8PWOfo9wC4JOy7mzOT3ci1Ei/SwhHxvF
5/V5RA11c04oWuq0l8CQbVbAYNjFg5kxZwMRHyS2qKQ5Inbel7Si3erqZMZM2GdKBhE+bXsMX+xM
EOojsjccTAkNa4KDaQR3LrZoAriKp2CF8bIQFWNP7GP+73+H94crlLq+o8e+3SrrUcARdI67FF/k
M56Fz8K2TNDuWfoVH93t/G2C7PYrmRyYHauxrqUQHjXRwOCHBOUHA0f/JvINZuNPNcxCrhP8A8UB
2OrrsdJsn/HnelDSR6BfhGhpcDHJkWYFW3xouK9uLQnKOi1dwqNYCOZG9RZ3mn81jA6m2hLDW31V
GCsNRfuMGe0EaVqY8FExu+GYFr/EhJ3IqhyBBUr0cZpPtBqlNbFtQRb3QdkJEYMBAhF/E97MG+8X
6J3HyzucjpBMFg4xa99B+AlAbrb1o4jg2GVAo7snNp/NnkCuJtY18wL4Ky/vTQfuoO0Jzt9JqDzq
8QupPdJQHXZGzE28DzLfaeV7lGhyqZzav8AyK2g9iDXe4VR3rTP/zR5xLJwDcSpJSiSI47ktua4l
vVy/G0I02Gw6AJnuvj39u7PzAKOwyxVa0LfCRrymtJdsGGIWt1rqe+VYzqrLNq/fU8elq6Sxnri9
qJ/aWiXj98SoV7uQ1MnYCzghhVJBRcm8QWu+1iifFkeHRH1VUcv4nSHGlu8Dn5OwjDwkUxFybVid
bA8iRa3an8OPwyeqU2w2L6TJd7OG5AkMA5/qdN2q+oSIDstTWQfDe0YdWuMgbRqMxRsA2/cDq8QY
U3wGRA2pIk0uTsSL0yajIRgWDbxMjH877dkS/3B0HzlrsKXwApe0UgMwJoY2m+brgfDmZs7tvFOV
L2DEU1TZBZlePwKQl1Zw5VZr3NhuZdwItxp5gPqPePM+RsPVLsZFqW61taMiGpjnp5GglpmHJN9b
lzcXJaaaoE/hmP+I2MlM0PL13cNbMd2XW1TK0BDLOfzk6ZX9elHyWUvhh+4FyUhLGAcODO9YbWlD
JDYSRCtn9GagXA6ImQuqexOSWsYz2w+5gRpk3lmWDBAin8uK5e0pi7c8jXtIycFMe/TX77371lTS
bfYHUazLU0HfrjogUouXXsSUZJukOh9TB65EVBsNBH2wHkV4LWrVEGHDlcwl9xQ7uan8pWkhnugB
PCvj8JQ+ZX3hFX3bSazRB/QTY/zZsTxjLDcSfnSy6VRlxJySX80KEykefRkU91sp2uoOmMmnm5ah
VEMEBfELVQDk/x3AUsNueX2picM78g9JkLJ3IO/EIpkRfoiZcb6dy/d9mHQOvZP8EX2NP3Pwb8Ja
KOjCHZKrcCjIvN/5fkUg2R+qMtREWVKnhQYX++0d3bs0kp64eOF+D/3sIb0QST96kS5aaJccu5ZP
l+A/rejtwmoiKzZgOFIG7OT9lpCyGfKHFF4EcBTwk/Pg42a1IuVHKRCYpk2JpuGAGVOrTcdmd4FG
xL/EvlV+Q7DmEgeNc2C+QxpRCJW3J/pwQncDfiTOOAmFAvQWjsjBiE5bdLH2jXLMzRE+M1ejHrQd
/AiDmZOYwKRgcJe5e73lHsnRaLMd/ClDCcwb5/Ti0a5u+JDf10NTxZoffo4Q4ry3c9JXeuLCGjzB
VoD5+HC5/EEq8AR6wSUq/jMZHdfjscVBjwE7ZtXUVDJJtdvy8KK7Rpu+6VtUP514Dt5LkCN97NNl
qkxSmgbc9etCu5iRlqH7Jff9bbPqcQamw8AAZ5G2gLOORPy5IOpBbqevaGkIfOQKyQLyGCxCFBCM
9bY4FXUUwN+tCiLDJVb/7z8fLR+ihiZdXXJF77VAYWMa+diIoZxk2kuwCQ/ptv5RBbTKEAKqEX5R
Y6YunZDVcLCBZ+qZuGKAlhVDPFhBs6fnAUV/HLw7UhGun1t/WdxQM/muFGMg9xTUEL6x4h0SN+tT
NIXxCzbyWctijFdnW3y/OVHpaZz9/bT6YAmkYTzVh37bvwsSWi5y508SEVnUZ80IivyKNjaAaRfq
FyTkM3DxByXqTP8UVcsb0tlWdTNypCjOqxZCayaN8jTmW9BfHtC75qVXLjp5GuZ91h0KBnFZ0BtG
weJWy67RO+OTq0yC1UUmfoq4t0yQPoSp5POSdOZ283ECi0ffZUPAdv5D352RVwiFxboJAQes27+X
zQnvh9cHOemgXAPe5b3A2sveo99CPTDaGH61DpE/bXOjasRAH6VGRSvLeX4q5ano23Nt17N/dtxC
5Yk8/9xmut7mdry5Lc9CzoK2EKQaBgX4tS8uWAQgfIyeo6680ZjMIrzr/ducooVTmWz87k198CSh
1aWgGYveA70SWBIU9V6E9X1NBAfUprJCH+e33ii4WKeoIHZmvnZYf5vKoblfj9yLgOQEVcEJuR0a
NL50vyWYuiTyvTJ1vU3hMwuFtJkW3e6GTpZXxg8QzbrM0/MeqY3qFJ9OoU1wwiiDGyMKFCKLbA00
vg+/3m3hcXgpU7zIAUMW7LgcYkw3OBwNIqJZ0KSsQ6RNqizT6pZs3f4e7EC2dHjhFR7CpukDxd4C
C0V1nq5Zu8fXcM3ANheJlFYbvYOWJ1qtmCScdmzmNsXjObdmg9u4lUnybJcHRlog7nRSwckIkS7V
LhZkCv0qTm63bmdBaH+tdsrUK4sLqPXgQeWS/T13H7djq+OqZb5D/FGT6pI9W1idmyFvoFD+dXMD
l0/18lyugva2xFffviiifOFv1B6NSmwSjMFbjsN7yM2S0Y7IAT66UF4ZlTzU2y0b49rE1QYZC5mP
yCRI3TSVe7UXmAY9SzakW9CdRxGMDR2AXrhAo+4ECkAntJ4Kp9BQ38Om7AnPxzzfUvjXDNnjGdpq
bugFfuKMdKSHSNMoVS2dYRA9NNfFO2T4aFf0km1hSH7v+9dPQD4nYpwjMfWhxpnnp9EnMrtp+j5u
MiSQenCSiM35YqMl2g/Etd/vcVOA5XEG7imfWDOEm8A//KtOtFxCpoQUINs+7+8HBIG/8ejgP25K
HHgTo0VEXQAJ4zrcfpTb/p7L5snXjcicXNiIP8l9xPaVOwsVgE+sjPeQJgguwacN/c3D0ZBPPdjH
Z/lMxyAu220wy4op17/A6yCabYt/JeNzlX9YwxafHStUqLVYjbW4lRp8B/VMWe6xWQxAqWkpOGyK
DtyPVUUfsxcltbkGfYarpoFKluOw7qe37L25PWUtCLj/UYqY+7FFeZAzdWw+i7V22hXOGut475Ey
MgfCUuE/4CYIZW6QzGj4SrStIffjFG95d1u+XWzk8yEsMcFUV80qVVWJXmDBzm9RaNwiffKyEfu8
9OEa/Hb8QguZGHxbMnylRPqOFxOHLmaZu5epqy/rHmO1nwnohFjIVo6mXWN6NaGXHzaKGGz7MQZR
yhHZ3TjJWXpEojyLG3ozW1eSUAIBLfBDCVFEgzPXdSJHzf6gglqmBdE/F1tG4BhMrM1w8xEohqyi
BHUYKBJ2UDWJMXkwzslOWD06D1wIaAilOBIfuem2oSTKfnzagM+vAqFWIu7ND5VNNxJJxfgxh1n2
+x5f2JptGQCUakzzw4/8rPj743vBtVKTon1CR+yZ+P8MaZYc/NOWHs6rwRewEBPWjAQl66OD86FS
bvATigUVL3Xq4KB1GpznOKZGaQ5YSiA+Fckr98/xO0ITA9R8zvViI+bDIcZX5fD0eOb7c+tr3IOK
Wh+aiY3/wHDZixLqRGOUh02lzVFnWtStcIppVHeGb1EZJl1GomTUuxqyO2krAjN+6ZxZ1L5kzEXJ
Sftv/hovoAHOKUs3756PoslLZquMwBXa58ypPoJNHcMzMrlqsJgCVqJjhnH8rtUxVbPYetG4X2Cy
bJoHJQIOCj8YWPV/V2v5I9bN3Ztcj0a2mVvM7HtobKcNdCwfxsWwm5I5+cCGEGb+P/DaUwvWOo6f
WRwEgb0kvv5upG7ul38smIcwcIHfaw/CILpRsX3WGfvo3kjSg2Fv8P0Hx3qI/rnkcEpm95DdSe+w
nNTcLfockMDEFNhZDemdwE6Crp6Nnp/Q3zptwp6/6h2apAG4jM1OpJyGIn4dvbIAAHB6TFwZjLmq
JzzhGq4do21pH0GW7rybAIzgNYdOVCU5LfvPiRfPiMRlrnv9+NymcgW4roiA5UesoL3SAEE9f6Up
LBEg3f4VfdJl8a20lnAPRRHKRNNtuSWXIjsQg+ut61zdtVNXuoEuaCVDjeLnR4DrMMjKskSNQZVb
eo3LdnTyiU/5rodYewz+tW0XS4p7PrUfCMZXKE2OlMsqNA4CDrrEIRKI8Kul7JibScfzS5Bdvfq0
QqvjSexY1yEBPYfcCJcb910cKc6LybNNUt48H4JCVw1hvsrnb1CW8k5WPnh+zamO0odygYLRFO94
h6HfVLUCPwREyrG/rBGKU9JvwsTndnwj1XEsnTbo70VM65/wXgf8EIOULgo/2K/caSO2u92hfBbV
Pt6P7mBS/Nl2Y3XGKDskrz8Aen/aezv5jVB2HWViXOAqRxv5ahi/2Iy9fPIb3IEIwZXmo5xtio7m
0W/byhMztFew0/9MXz3agM7AWj26pZ1hdad+hryC9YJm8jGBaCVhoYlw1LlEKA+Q3Qc77d1JG7yV
DnEWbcE1XCr34Nh5VV0RweKvhR6TViC0s1Ip6JQ5N6TtyrP/Cd+BSOGac32YWhYE37P3qpEPqgor
L1zDQSbihuwCKt5QX9gEzvGGp8GZDHZncwwAFGuRPC46yb+yMtHq1Y8NDTy3GaVFK0EUItkOLcVL
jtryhLXPWYjbwDZH59d3RUXzobd8Q4wmpsUMxUZVKU11My6K781vnuoZYiflA5ZVLnNjpc9mGqSR
zx4ytrnRkCd5uZfQp2uDc0vC0d3QB3ti7qI1ckS6Bkv/MypFfbTQlgbI5mspxpuyOPh6g90IPwW+
GiqXNEq3Wl2fJxNfXwGWYKQrJ076VA0WwtvAxLawlQpbZIw72hmKPs1gLLs2OLeGtrHCuKYNyrFV
6cEET05pHdBVDV9RQVsfGGp8VAPBFRk+d/hj3TSxEOn/ufeUaVlE272GTUanZjQnHseeVv5cgKD3
w8+JXE0VnQcRlpsyXAg1EBzULLN1PQtcF7zEPF+dcE8ux20UvhlF/YLg5wHVrTjGD4y/Fr9cU9Gh
2vWol2hn4qsGZOSwk+t0k+stRq0p2kMYMudQUNRaGGT6ZzQqW4Jk58OzEZP/avhjhXmeyRmsxJ4Z
yJUw4WU9vI5Wb1+9WtS3zPS9nCccnLm1T1LVMKTnWVcV+S94kUzpFPXT+nIGEal07/bd0D2ORleL
u9xgyPWB8HZ6bAkGkzyAW1k4Td2iaq/MtPRa1Xqg/575iXz/IXlSZfo3Y3hOGbjgfzIF7X2G6U4K
sAJvmNjPP3wpOnWLqVOTHwt46/tuOGdinNxFEBDqlf17PgGrRAHtdx5mYTyLUV0WkA/gcbVpAxIi
HF24tSPy8FWJ3FkcKbNi6sdYW3gUVnv8oO9dqMc6QSNtYHNboNj0UKhNI0uvhkARYID1GRBO1Mx2
2QwdM5qVcI37hjnmQ0n9h87JcAVIb6B+8h5kjTOQs50X7tT2Y8HTdhIQ8BoDkIvvTHc4vcpsh35p
JCWnFOCgzNhZqDAG6IxAX9tKBXl76ckrCeIrmY96+/OirO3zqoGqkjYT91upjsHXsb/x3U4qpypw
pqR0S+O6FH3r/hvVbgkBqde9Rr458tblZ2f2sVOokEeytbgH+GugSw8Mco5VwdTwZfUlDzDVMv0H
nWqFV7LkLuptCqWvGSFvDSGsOHh+isoGKDI4Qb/oDgrV5oklYYdulrehpkVWfjRCrZKRYjnL5rTV
9Ke7MF9VogF2EpaodnqmXDTIud7HgVk6A4bQsxAVoRXWd4gdsH2LqVsaSPurO9NK86+XqoOK4OiG
yDSc9C6FuK2mRKWZzLhPxfWJqf7cqTKoI8+cr8wi4V1eOKjDnIzPSc5dE3JXiYqIvHlTT5/koI5e
ix3VIYALs7Vf9CRJeLoX/x/84/yZpbmhcWaM5zyU4zdmY+SRO+4XDi7gtBiFpYk90GZoQzio5J0z
qibjdC8F/efbjAH8FLERP3QdUP9z8DWGD6l0OOHXXWdfUJoxYb7R0lmNlSafm5hi9SFtrC1b26ZV
Nxr8rI4rIaJl12DD7BUJL1YOX4AxJJlW1Y33e3lo5PuZZQ6Kbvz4oZJzNTt1ErL8rOVVIKdpsoH2
S2gY7OFoA3GSauUQ46NfudlxyE0n+mGsEQnr3ArO3SYcuqK2qCqkBJv4QswSZpNUfN0DCPuUJU81
q7opvv1IG/1RYIJadul1yfuKRvV3jGOwVlD9ZZILfyCs8/Dhoydgs6BuOPaZWzk4BlD1g3pO8Hew
+PpfzNOnhK0CHojZNHtD6TtKljO9jdr+1BcN7J+JrUC2ZmRVLRiGQW/VUADlBwFxfpoljtbpgfBP
gP3ECa6AZJA29kRO7NfFV4ItrHfSjW+AIKzcThMsJiKiVjVbfC/padP3b36T16SupGgcBIQS2BDb
9Objmb/vMV6ZlKCOd5WSLzEM8ChJ/1TSgbk5qpza3dczNkXzs26mZUjCnBQVXKIiTg9dF4ZChgKR
9TeUZUocTumb1aZVfRCfYZdHYYrpFZSB/EoJOlQHKi84Lh4uSejLFfLtnVGQi126a6/9Jtc3hcMl
lBCqZ9c2WKMHTPfb0P94dIomfDsbxiJC8fd3JChW1ytSuYIy7UZ42PNdf4SiaKnA5agFA9H2igyu
4dRuXRgfmnDEankfvAw7YGmZFZnKOMIKJs0xdxxJrlkj6u/uwK1BUMLd4bIbSxZ06dabmma6w3wY
8sKcS733PViUs6qQDslAwTOPjD+aS9jrNwZmxoOkZ3hy2YQHGAsi8sCWJLJKU4bCr9Hk4i8kSER/
GZZ50SXUHTMpHtNqwf9CMCa4L8nvV0gMQIHytwaK3VGH2AmP6CYYtHw63lysdJYDndbJCoZiLwj1
9sY4FTGPI8M8atTsNy+Vy5hJIPaR3utihHqiP8cdsa1kuvvYeb2q7Cl5eVv14bqFWFkTV10tdw9Q
5b7qp2TSY5bUY2mPqOpOfpXuUW6tSZEx2Po3tR6MUVN7XO7Sm3Y1rKtOy7CSfrgtsU2j8QfzCzHw
iKYI7xZ9K+RzwFZjIFSRKpc1wKRRIjbW87HRuSg2tw6zV2JxkQyASC2srAjQ+4MUrihrmHkpqebP
YypJMTKXuPb1BaoiFmD9jTpTDW1LcezX6O1yFW2OZwsqRgqNN0TzbKrT0W8iWDIlPZCjBY1jqZ8R
1waeu87eDgEfsnj1GGbPEkq7YuPvisImZ4YC6CjGb/D7LM95DSKK5xHZ1L9a0UWFdibFlW2wEiMq
9lFiBVz3d2N9hu5iVjt8S1k07qzK5V8xKTUdWgRsDVPlmEM6g1Hjrr4yh4uPML26E+GPvpdYHux0
yoJGDmu1vLhSnChAgKwsJnZ9sV3KtNZYecnrSBI49kjzfnrG76ggVdiZ/QOEDBAUU+ZMSzFjiDqW
ry90XzoWjQb9v8plngwX3NpPtYew+xb6VCPO+ZA/zSyNP7CfYkhbFtcqrUZ5DmMPmd28ZfV9m02G
hazL2m6lUfiaKVn2NBjwN4qClxfXhaIxZCjyHXgY7gAb6pyQ9DCvXUOU6CdOTfnWscFr0JrDoqrj
Il+zv+Z1AMcNh+Rdrcb60Xmj/7826PBaghrVZ1MRcH4GbsUHny6wX8aK+YN6t+u9/+vI1oM6FDuj
Vz7u7AiEkY1GuT8V0PdAJdsixzhUFLQc8AtKs/CtIh6lNpaUVE2R/P2saCXumVvs6q2+qRf/x5eR
JL2G+EL4RRgi6gAi8Hs04IbaebSOSRmHV/jiy2HsM2i6oeVZ2rV5ZwxKHngwOKLe44IBPH7/SInc
QPJfydcZFrMq23xUAgEaP8eJcxkxsAH1xcD/BPc68xO4FSKNAhD2WE1Kq11c1sA26e5wJ2lvSr/c
5/TtHtLZZ0KySY1YlT7ZPkIM+wiDP07ezKxguG8GIlSyFeRvcMrn7OJvQvwRDpylgIRGpKyQuei9
8SgW4F2L2Z97F1UuB+4xXpzyj0Q+NmzSrW0xXU+f0HaB3fu7jfCqBTJjJ4oBtyhw/Ixn8e10D1b+
wRee37X/DFWk1IecXq9RIxmF+crcmMySdMBH//2ozJVWRyXB3MZbqldzYdByyr5n027GtY6N2Bt7
HkIYyaqWnZNi75RVD/sEFar+ACqW8HhkTKpRRnCU2tHss5k4lq9XBwXE9ENfNZkz8iX0e98o5am6
veVE+vo48rvgeA6jJFcbjASx4CHbWAA+lqPQJvprbvM+kdGecw42E3eeb/7BjSUwk3T1rWn7DRw1
hxmEJ5m2VWpW37kc/rBEsgMWwCRV/FzQangfZ+Hx+FViUozmLhkb9M7TQ84mHcU1eLuW1Ebhvnuy
vAppYzsIC/5dB/6vXV3jYuO2hPZwVlZzRH8MXsj9swN53RS3AB1PwuB0VMcDOqx3MULrfqv7wf26
G36XmgXcuk8yt2YC1NEN/5zsmi9UwxwTxc+GlwqUMhUxAglQvenn5h0LR2z4cieRnvKujvJ+zrig
ObhlF3uyBZyYh9O/5gAOiE1vmym6Up8kvKKx4Zm1NUy00t19zkHwyYmXGSgGFWPtA4woleXPmQBZ
G/D6ApjVT1VldXm7GN0edcucjsMLuAd9ukh0In5uc1Y3PLU6XfzidOrhskYAIzEAkQiqfrEDKps3
St+2lQotwu/i8SA9AsMCNzGTV/5xogg8zjCGo89yvTxR8iQzBmCt4rYjDjTr2LlvNyqcv6pn4pDC
IP28YMHhIPn5ZSVpbZV0bPIsYhTlw75KKikjejl7FJDUOSLDD6hwLSMPgqHTwZ5n4NS6bLYj5AI2
DTljEHnRiE8SAS89LxpXEDaEEdB7rjgsSL06t0lTK3vxMz/qcxko//c0hYp6r6SD+njm62lpLAvD
Wffvxi0aCHLmBph0KxleoH5NpXEj2vTdXnM3RB/7cVyJPVTfe4z4/862oOYP4wd2t+VzpsCjziCk
9++uygOvF3PAO+k6GLTin6y3nv1JNQSfoVl0o7Lvl4BYlU52+zPT50+nA5DFUuC3hy00w51mjkdd
oDDbxrutvOmtksLpsbMszjWj394sHLnSoDpmGDKyRlX3iBokJOS2ue7XEqyHEIWQnEjWcTmfUGxF
b293+xxiS4bwkQRvVdcSoIm8NW639ep9C3/FgogBQ7BT30Db/KTkCx90G5AfdQDutQUySeoXISDS
BSOe490LcuX8NWJ3RT43v6NTIWCE13kfepIyUM0YW+Mcldw0V2NpXZeYmOwmLtF/3GFlIhxyI+ha
vUajhT4F5PwXoezOlHyz8CRGazYLMHHaPceLtr8CGUYgWyx8A96s7qGNfgA5BvCDfnLcemMHe156
aH//AcNeMDVj8NmoH5xp4UA+dVhfZOSqMeRDkM6AJbfGeLFs+LoxR2Jnj3tF9SJ07ZMi8BpfYCrl
VM4shq/p1eXo/6EXelyTja8MAESKAcRmMCe25wCHA3285ajiTPtZlfpYgavIUhdIrd8SkjAbgFp+
dYKDPdbhgZmMTHudVtAWmEnewSsjYL9v1qXdqtrLMb8Nqaf+5uDPgtrni7guxL+Cfxf/+7qrrysc
jGTV8nIkBIYmfjAClFkijjIgTcyAvr65iAe3zq+csboZbv65E5lwWYiR9vOUseyVmykb51FABJoW
Jqt7xu6qMlvq3kL0iayhM1TYbwNrhZZUzOaE8LPiJX77xjDZ3LMMTt4/1g6gm4rvXRbmO6i3TXUf
OYaxUthTiVp1vfJTLj98cq2QKmtO0UoZpEyBCOg3okK/D8bMk/jqf318qwbK+wOdFBg/M9cnJNvk
hR1aoQ/2KXn9zr/jUahYf3Fz5hp4JLiZjWOkcHJiaQ/lHFFmp4/9wg/Eb8/JHErA2DCQGsOFo8zp
psQK3w0AE6S2fuKpH3ZZkcY6YSyH5gfGKrjX6kSagh8Xi4RcB0znb6tC8SMiCZyzqzLcGoxyMcZj
7KQOmUYhI3mNXsFMBLXhyiHx9cipGzVhHm+4L55nFNfjX4CqmbrMqPhIo0gP3xbNlog6rEHw5pRi
YJlDCNavVf25jbuTVYotUZV4TWMcoUXl1SjyzORXOAvJ72N0wgfWq4UTClKfTOJmlrlEaIOnLznV
49GQL45PdhcHMnUOgddEKt+OQhhGDhQZPZuV2kzJUNV8Q9zS+AqN0sMt2HYcI/XQqXqMpUkYxkij
0zwoAgiKN74k0UbsGhh1qG73NQdgxmxbB1da3oc8qE1cL2GWRDUcKd/aNAkgDLJxyWEtKGpr99Ku
jI61eW/fJfK27SU1LTBVKIR2LG4tWZkWsnFPN0ZjfXWQB/rhxZrXoLmCQG6XCCq6ikO9cSgC9Fel
jYocxBfZGD+wR3Rui/iSz+Rd80rMi+x9/K61OwZxlPjcyb001feUAwhed8MCTN0XpF06yrz3cIef
MaoEdI7jHv9xN32DBb2oBGpa9gRT86g4RjVh2/MHQvZ8Y/cG7Nymet7+CcDAsJFLPKbkcc3SNFnI
k6uGGehsIU4ruvVEmEV9F/9dzM6ewdeuXUl5hMpm+Hoi37o4c0TtDC8xPo2QtVxANZqE4sHCAJQM
mSTA57PcchuZgaBpSTqlJUajflh+sLAbwnXIHXY21U1322bRdCL7HlOuvz2XcwKPTpXMeVxS8uUW
k0cJQre2DrcFG35LVc7xIqZ8XPa5+3A+O0sWWk6xP2HKMo2g9dBATVKf5wlQIEGSTBnd2/T0HG3B
8D/L3Bwb4lbPcUIhdR7dd3jD4WJ5M2mDjfzPlb61PBkjM9cFcpRM/C13TVO/W/sw3npxwGuC6zgE
H6X0KpPPub1T1i6/Ky/xECmTEhkS6MH+ARXnI++ecmJLVy3aVrbQyun30Xp94Uc0QFcCSA+jC6Uc
wSdqAWZq+g5Nuyy+lxhHGszF2MTejqq4ZDHVGn1qkplWJUB6n8Glw4yyPf/DjA7uHzk1FbaCg1Fu
0KI7FfoF3E1Vldah/NSqgd8hCkoXlKKzXphEAK2Fk93kh9LsoVx2xT9/gelbk8B7GIGTxNpqLGTt
xHaQ9Vvv8EGdWresaa4nudt/J9LyiVcl1UjbzpD0Q8tkR302DaPq3fC0whiRg4cmYN5M4YE/pAmE
iot5mnnnjkMwwg4wwp267s/2HxlA2HZ24pnL2XNZRV3yAFqPyEewBWZm2leTAyPtnwhB2e+Wndw+
nh4VkTNO7VuzHPozESbEn5cyqp7mmysowXdh8A1nTls9IwiPnJmeTmNLMaH+acZA/qHzWK0J0ETo
7S2VJaYv8k1B1RcFIcFyC6ngWMIgAEPW/5XmshULR2JdsssqBPlv9j3J7tJI8RNjhumeQm4EG0fN
4F9P0FkeGY3PuI4uADjsw2Yj2uQ4fTXFSSsUpNsAhrAQZ5PJMMpA1SojAFeS9DOHwSTbgwIQVimz
hIc9L80RSpsX6G/AyPAwJGf8ewrldA5UQsUg11DrW2v8ZmA149Ic8QM+yd8nk/4ezNByykpW05wQ
Aqa2UKuselmCyRcr+VvkcR0cxwZWmX2KEAERkZ6zDHqizQv2eTOTVdrzO4yj/fmmy8ldt+Z2c9Cx
qf2cJvxLyKXHoIn26zcEe32TvbkCSv4PzYwT5wGDn91QvVSB61V/o4wNni1Xt/DKXYw4XxjVciK4
jG++OtvZnuTxyZRpRCnLN26OXzXccV/Xlbh02qhl7g0DPyCE6RvKNZLk6Wkz0mObZKXwyg29zKJ1
3CZc+XEZNrH4dq75JDH+cuMRE8rO7Lf11Z29usGqEh17d4U85AB9ysiGF0CBbkB5aIOs5pp5ndXa
SKfnu2xTFdy7E9Bkqp+4fJQSpIbgKM0gESovFXRV/PSuD+NWl+Uuwvzhfhhft64QNLmUqHK+FLg8
vRWht/DrejOVBpefEKuBcMxSkZoO4fgnpS7xb/9/rFTY9/p8iWgGmVoxSMF7sICOroVrIkO5Grnn
ti6xk5/fC2B/c9fYcx2rROg6SwoKboio84/eF2xAPiy7JAr9h0sDW7NuAcNA8PXSbkHFL0b0RsHr
ArFe6bDkrdtRofFFCzwT0QLVRsRfPkdZHbXXPbmYlWJ9qpSMs7igbqolfUDBji822E8WyeVIa4Zu
kLMQ9hhQK2AwuHnWNtt4Ym5Nf8PrNGBhgxFwfR0KD40fjQesvnfkfWPQw2IUjEvomA/5l9H5/sj0
BXV9LP42t9X6SZdN3f0ye6kXHo8dey7+CxW8KJH1Tz+hkX+/jzNDuV1iAlE3R2YY3zsEbxK4of/6
YfHwr3B2hvA6zyfRcRGdJHfyV1uLtUtpInudqCkW70a/uk0iX9oxD92I0q7M/Dufb6riYBxG5uv3
/GJ0b+NC75vXe56BwXyJ2sSHz7nsb5IdLiU1uXE54b5dnl+Mk6odIzzLsy/XcR/utnsif2StxDwp
5kuwnUbMELxSWoOU5N8qFb1MacEkbYM+bye/mId++epOlwCO+yErqcCHb2Uo5lEMvKWUNEx41Pw4
A8GM6YokKPWtobzKddThrVXTtHZ9cqgEzUqaReja9+7pKQ2FtNPs21G6AQ7xSoumMwd/ZRXAkYOx
X4HQKchrRkiSTYDlHsGcpArzpZV3FW+jjnumLX2Zu8t7Y/3B6FRTmXyExL+qIPieo4MxoGQ4T1Ez
J3o3DwpNlVVxJeXg3pYcqMjI5nJSy4gy9ajQp47XqIdzWf7YD1WrW56GM89BFCOO+N0+Nlgk6Q9O
LI17BP/02xOQKw1qIRvfDEb9X2js3Q8QXbZCyOHiy241TR9fhLNzkJ4cJGriTUMoW0gY6St7oMhO
K7rDQdQ1hkwV8xiZu4In09pFWBa7zsDjZ0thRNjznM4rC6uiz+IhSm6lMOjELqFEWUGSAD5huwp5
Jx8evcLMBhftlsheD/PmUyMpGWJfApBtzIIZI7zx6DykJwghLntLyrCU7B4yRB8Zk0KHXSzy3zCm
D5L2KeD8rto17l2psmDeshZ255bCMwh34DWWG1TK0AFUhavxtVi6dwf5CnhKk+cWpA8rfYdoTL+L
37a9A9xjWAEQKyEOWoSd97X8G4bgvJ0Z4/JzE6iqgoGYbDurtvwsy0kpKtYuym1HbtIA1BErkwyM
G0JmiVSgWVv3fqb/1GvXLLQVbJ9qlyOSojnNKhhXzN01teCIr2aP040O40gVHdYrHKgtyI/SSq8M
LqFdC0Yhkz+zqksVcUBs0P/tnnVExnPKUV9xxzrAMGHfA8pfSIPG7FLGTamPqk5hUN4Vbn1jTiqy
SJxEaooqf5SfBgb3WQlDMsIwchXt38S/canf/5Z8v3HJmkh1oLyaZ9jTEnNZrbt/zmtWi3s6shdH
Mn0fTaCoXFlEQC1aRpCFsfbpRfaaEtSAVBUt9HYClEm5NGzU0wOajb8PrbcNRJhsC+NyoERRpO+4
XfXWkF7eL0pgqvz93yNO4e/+5gJbZQAF664EwEhKDXBQ8qq0J8jOmY6IqD1gmGSqCT6yy6YC8Pvs
2oRY2MJ6ElSFG7qB+SZeQq0HKSxtmWzI/NWo48OE0vushKfpXz4IL2SXN7MGsLOuGkLPwcPnhw2e
hpU2/DkNtKCY2nWbCSRu3HsbFROSFOarhFL3LcP08d/oz5FiXgWVdLKykjFMcSHAIO6+lfEJ8vWx
h1BtA/wwDiJhMgKDuXne7TX/FzO/xyRTeKA3Ivgbr9rMkve18728ThJnt+wp0w07yUInI7N6Kq6i
jE1kRfqrQ/Mm0u2od4A+SZRFZ3lx/AHsjPqDPuYr8CGzYm4s8jBKnj/vyX2/SdSuYoOIboWLJW73
qrLQajfxnLMU6/ewrxBvUfjRr/HhWk+H+M8E5JcNmIrBJN3dz7HMrlFs8S8d+DWd58y9k5XGDc/1
HZB7Ll8+SYMufwDE64maa9cBSHyccLWijYwvKFUUaN6Ij9+6SikAIOvNpU2OIT4vbDBM7XfQ8NBB
zkIIT1jb4IjE5wWXTM/2uPokPqa+nqxRv7oH5xBJP62hyEgHb3JIvMlJBnSlA5SV+oDeLsPcrwTf
iFtim2FEqffwiRIcKTGWHua8pKsDkObNsi/B41xaqxKmmusQmx35TREzIypIql+70kHPsy6IbyTa
op7kUbikY15HEIzIv4YJn0NrUWoAKNsTkjFh7l6PpXYX/aLj+Z+VEKlFLan299vbnowzAqIunYbO
VIUiZLkBs3sFZDPCZjACZDZ4egOEgp47gvp7FheGiLzr5hdTiXlxYb77IdmY3jx1nXkmpGaLcqwb
FYz/rDpvIpiRzTIti/rvWqlvsBWjoKnBhipxBQet9746UcXYpn2/KtJNgCSo89OOFfuBUu2715fd
Je4d9zcbxEJLTq9tS1B+mcakUV3O7q5XoPN/Km4zQcuA5CW+8KOb4EV+9karpxRQO02Bog2GAsf9
Ir1m/5VySANvm/8g3tpZ9ltNMk99p7Ne6uaiotZzI+fp+qcGOlrj5zRA4RaOpsG1hcCZ1R5T8dvK
WXH4RK6ml5NT/VoIjx992wk+WC/E5yVLKahdz679qawx8THZIrW2lk6wSz7EexwXjMYTr0hAE5aJ
r4a/59dnr6JTYe+cHr30VmAYXQBlQ4XzSvj1R5QaXNEs1tfEiWc4HFojP/pYuU6BPXB3IwpM4z49
s66eoj1I61K8wvznQL2Vw15sIxoL+ItL7WOueswZpA+6541oAd/l7/7aVhL/2tCQZ/+UjvGYbnZm
a/3Db4aceIvBWNgWpFDBNs1i4f1yl96XR/r1j/apNVcwUH1Rb7znDY65k9Yw86rVlO6pK0UJzkPc
j8584NhsWfDqX/MfyeERFXevupVlwVSqWi/R0yqGUFlMp6wiSh32ofLk9hEncVHfqENzPzFKRS32
0a79j+e0O7lCKa/RV+9oW1n4VQQyOzty09H73yTcZhQnAQN0OMSeJl/meCRBiEh3HWQnK0/rMktm
73rQiyeRKt9YvDD0u8aWMvBUh5U1K8R9TzpgtOhW949/H8XJlEAz+kYrgR14pUnbqRE8DYq09yX9
6fIfTGtZv01muJKZfx1d5ygvhuZ5rSQxUBvnrAiCDLMMbCEmvdRarmaC6iqKzJnieIKL64xibi4e
XnqDFrwwfKHeOz/btRav9J7i6Rd2uROaiUpS0mbnbncE1yxDNrv5QIQKNaF/je0VG9Dt7UaML7px
Z+bgk4UjxErMSTOUVUdqgmNsz3LOzfFe1FkfrrLElJNz6QnXj3mrsv4LS+Cm+1Wrtgs1R5fknS+L
LrHS/fF3iDEBm8BBQ7M/SxSdMludIUaPEwm9epZ5UFHVAMEf6n2B7zfGpyZ37i6eGdKpr/o6G9PZ
haNBEX1kFvOlPPnsaTLz/e73pPQHdHNUiU58fDSSgZlLn+6REVIDkiapVZl8d+eTXAX/bVh+2s/L
3rQp6cHJWm61GW/RP36fplHRFgEIGQqJ2GAeRyjk0QhXlq8B99bQRIR7nkFdiCVjTg1+dCDyqpS6
yhseD6wpi0Pi6J7jWCrvATkNk9bkMbm+Qx9S/IE6ys/wd2XhFbqhJLO4CsLOKcbeRrBtqDbCwk5r
hSJhZcx9qQYrqSGLHAPMuCVR40KXH4pOIBz3oTgN+lUszIRL2yisXoPdiKT2TzSw5zOen5shA01D
uKPYZJHtr6eKstNoXAZI+w53MR/DJ4V5OjsM7wQcFvKmLBSAftEeYxzkQe0ptBpd9vUpjDz3WEDZ
XodLP3i0DqZKPFr0/ak/4lLsVTkinxNcm8gYVWijxslD0OssC90EbjaQbN1MPdm44HKEbJ1Hg8jm
DaU93NMCNDFvI4RVMMTAwPMU91IgiOUKL0n62gx7YeU2CGyQ6FjfBZ9Pjo3oB7GMi4nDLLlpKWzT
l/3IeFnJ+iKuyQhAanGSqCERkhMP/TCK/IbHO3gXkqoBwljPSwr6hwYaBBCyh4nbg/scxcaB1Uv8
Ih/BYE/ydyr4yjH8dzj9XFjyrncaGTnv6wpD/xowGBVIpQgJrm30QpQJbeyLK0K8pMxj06HohUPK
J3cR9uVdfeNo0ubP0t5VFsr+B1mvhaUpf4dIpawL/dP4/pG88VjcBwkWJBfutsgLyhiDLTCy6Kmk
Dop0uSvVYd5jaJjSpi/ZuPhVvjcaNa9cg5rA/nBk+Mn1X3B1Yf9ph2uUZwXUkdeaXeBIVNz+oYVf
P9ukxHV7dJ7qAryz1MsZGvsvm8MvRBQwpNhXU7+k+5NN6aDpeTXRkBdZ2IAMHvTKUC/OTYfJ7DNd
JdBzqE9VdaInuPSJ2+VMtLCokydsXBITv4QgMujgMpaDAAQH9qV/uw0DlfBxBk89XDTsDB2i7DBW
XgteeZ1zRQ/4VBqQfSSFJZiqdJkTFpRS5pma2NiS1tcatZiNDx5sBfBozOutegcS0XA/siBSkc/A
yE4Qg/T5xtEuwyQFlHeHb4YacJEAjcexr6RuQYR5VOikoGmUPu9pMRDFQ4hVxZGmBZ7Sq6WKtgqa
g+DFObmisGfYCiVwlgz0QEORjCRaWhwSS7RlpQHrGI/AtwKtJVLeP58BYnvRaQ88/DmIwBlPszS8
3zWtHVWtUNbIgVFCAzMSv86OdUuZmO0Arjqrrl3xugv/Vt9x1+NCiw1mJ+ZrIJCMriUZlpKvhKSo
1P+Hbhd8paZFnEpM7tbuT/+ry69IMQpv+EDKYf25x77SdATUapLhoL/sIGpxm7aew8uz9ydSSqtc
+Yo2hD5Dt/Bb3F9BrpEGMiU562r6oaCP+wBYoBW6OogNDmlEwf2KdQ5guWbLB/9KUbavJ7D7oD7d
UsOH3+QmBpdW15iivIDTMG8vVPfULFh7HVpar48Ud7cpH7xau+yo/A4L699FJm4nWSKhCqgN98eH
67VB2fwoo1rsDsL580tfXpbuQdKAolyvIYsoyDhGYWVBg6f14aK27J5g8wR560hRTIB6u+MHPnwp
8JJR5aLv2dCPtXO04BK4AhUPJCH7ucyByuncCM/ZAWuzg9bzMGXOSSuiN/Awpds3ip8lsH72w314
lGMQSu44qtQdeETSINTdSj/P/J/YO5a+rA3I/NrsEl9eGkgIre/Ui9vrgzPhBdtzGdunJXDc27P4
H+yYXZ2NQajS2Xe6xJ3KUApWoSj2ymk5ZQ/OHbxusBXiirtmVU2fhfrqRFhx+2amb3fFxo2+F24c
4LE2XMkTS6XT9ACVbJvFiGNz1ztoZG9S9+zAcQPuRIDJYioLMlnxKf4T5y5+awTqPIjDqNQS9Kjv
wjS8mngNaIGF/buCWl47+iSte7M62cUd5NlxT7/NqUOh07ULwo312VWRgEV0XO7i/FkjNwVxRNur
wgZ3GbUasfu7bnV0Zka3v58s1Dsfun0XpeJ2OQghp8Xhb0K7z0YtVp0Ht/pPadcyTn8TEPkEtIcT
hGvIjlmS/G0ANI8qUiFxduX1Wv/Jxg/7l+Iroxkes7dHa/tJYBlUCyyD/7jXGdxSgpPd9DmoZ4sv
p4RUev6HnkrmsoW+bU8aGtyofkAW93hVz2aUDyL+XYBQ5vofBhLgFelYtjR2AKkEWyBuvCd1Y3Jr
sE/9KdqjlT+PinrA+y5tRvRNAi8ndWgxJbfZX1xBW3MycqDcL+5sCANZiruUodqlnFJHF7GBK9Ot
itPIRELuaL404BZpDIlP1BELYF8USADmdqsaPXoaqRl7GEnPEpMK5AOrwlTEXslMK+PviC4PIo+S
rhXKQTKnbU1ORSlPPHvcAaIIqsNsfrgOMHDc0Wn5fe5bq19wAf+aWvYVa5S9EH7bjh5iT4i3cDqH
SWoppxRMKBmhwFSfHrBG743G+nxG+DCz64wphixE9hEwcvUcJqRLkvoFiM2E/2SZQnfHC5e8cgvx
R6QlrcKWtDPIviGrxvPsz/t8tM3tR8Y+GjHZghhgbryn2TlGC0cP0r1z8uSQ0sJjzDhS6S0+XxLo
Ae0IMvZMNr4XuN1aHQO/znsedr8NCENL0zY5juA6rgQtdIrxnSxS2Ev2xumA96Cf95gJnoT6qYKy
fN8ISggXEEdWGogyKQxNoULlNISqbc3Y0bQU5h8lQ4K3VsyirlAqdDt8o8i+SC7qJMg/LfTBMNLg
lT0a3AqbERBztZC3ZHv/Jerq1DSyHgV1/JUkuluUBifcS2+hwzAQ8+xtMypA7jA9eSQlqFD509l1
eanKi2mdJPaZqAnlz4pZaoUsqCS0em1e1TNrBb1WluA0fOMCFGLsO3qPsIsfNwseq4ahfNFiVMQE
ML9iXpE8KHZqCSpMWXbIBbLElcTqNKJCOz+D+jxq8GRuuUW9ReteNNeZZ/dzeTjM5f1eccY+evAE
dLImuBHRoFAfL2ojxszCKXvrN9pN5KG7w2hGmXbeoHdBs3nbRjGW11VAmCj/bIIlPFjRhYbCiK5N
3lzl5orhpsCqsMSI4Ee9Asnfp447FV+Lr1r6FN+gzTKPV5VJxtpKP5M6At+OGZb/BQLYVbypzSAQ
7BWO6nkgJUDQM1R2XD8aoBHZHIrZeszX8EmTLs3EJ6/1m5blNqXjIRSsrXo2f0VCJMi6Kj4a0t3J
/qRB2Oc51JOeOxo+RQr1Gpp9tqzk2A34Uj+fwWlA3OfvRqOTY0fBB+VQTmnbeHcJmK/uJsSsdks+
+aVIhg5LNGRfjSThIEFH5dzecoL2DYnrW6YPYqYkG+MbWPox9y/u98J5MaHvs6Tf0QhdPeecyg9p
WUbvZrGGjycRrcnr4/hd8nDnw7tblaIOr0zRzHdeFhoO9/w3ekZcVlp7mMwptXy/GJS1Sfluu1DT
R9gu8iHCNFSVl0TNBgCVewOTsBTfscI7OgT9VdHgRQixa0fL8npj3zF3dX7VROv9X9OP+xlM0P2h
6cfrLpqiCj8LJ69niv/xt0+tDqRLmmaHB5U+Pt2ybWTjOyCL11W4AeYA/Ft0W2cgdj8tlnPxfHqu
HZRwuAoPSgTy+J5+zoJqWK4z8quMocYiqsJ6PseYwB4BrEKEgpDq6ckLZ1ShFQxUXQOiriqEgG8u
mwZGP51XXrKHPYamCNBiludBjR4zP0cH8WLBLdeyTRcUWD0ywSTczTUu+mzO/Kg2KlzXh9YKJ+a1
bcALn5FgCG+X9YoBGeU5r4DK2bHA/ZDER/iGYt5vrbDk93+EX3dJ7mOBps+UJ9DRrOaQ2yxI8oiq
tV/8qlvx/M2qeqZR1cUiNg5uZmeLjiwZKYhfuDOm+CiyjIGT+oyydMPpHeM9I8c8Y0HokZbDwLK+
SQeYdEisQCTUrdg6n0o+4e1hAogSafjRyoMsQj1J9YDuRLm39mjiOkJ61C1BnP/mA6JH41KfrMDo
gbTwH14NNnbHZMj/5GYr9GJXSj7sHGYmEmoZvD/BXLgSTRdjf+d41COtnHrIzjkagkZ+eGuJfbH2
QFnBilUdioanoQxhFws1+z39Eemni1hUsYhEPrB2rXpj26cEvK75F+dDCTa4pa4+2pAeDLHMYud9
Y7s/lGN+2LeMWA89ilap54lvUYKCcBkWo0INZMWol2j7NDbrapL25yr9iM0ordz4MquvzIawjdPa
vr84ip9k4PGHw3fK7wyQtAvnadrGPsroAjAZH2TfjI8y3UosS2BftveTJDOtS7PMtQr65gVOdBdq
uP5yseatAa57d0AP8FgcYFYY+yztzHSujqH0CR+kFPaP0dyuFweamLpp8DXul6kTWYLanLsxnXAI
SqEhJQDhuVgJdTYPSk7d3iPkTkzxOyQLKj555lFxGIZw9WgwlyzVeen1Y7RTlJ6HXv5S4RVsXuYZ
XCkpKvacDTcf9E36lFp1bX5F1wurn5CpxoO28b8/uIyw0U/YiMVtJnWMziGLVo4WpnnS+IiUrnQk
PQNqA1QF2+vJrE0uei9Vxk7VNaefq1ZFf5VtXLfJiosQN0h3BDLmBhixCAuvyQ+09U/R6jQas+So
VzWyW6UTlUCtqo3pBBsK2vh1VLNpZpZlbIJsBIYgjWkzlEOeHE5xSLO/mIIpL4xgLKH8Iec9Z1mJ
wXnkCqlrda4wWfQazwTg0Usezu5hZuVEZiWUILclxFbuU7eOfmH86bRpyxrUZSPcGdf849Qrn2OE
gvuRqrXovYJ/ZFAJJh+HcaVDNVYgNrKvz1b1HFZr0LSJsijsireLddsM0KMb1R7Hsb1cUEyDXq7s
gWtyLLqze8ojTwbcU+tK3QzsQvmoYtLeHpwrUUyOY6bRu0EiF3vmYF9foRy6OfeS1TCY5FfGisA6
hvn9mzgtv2YM+tJUJmCH3rqRhoS7sldSYBYc/SuifuKQjev7xpv7bzKz3xvs/RwLJBKiL+3InO/M
ZTK4dkx+NwBV0fK2tJx/43+kGfKeEBVvD6R0wv35vjQbiITBM6bI1ASNC0aZf+EzjTOffJHrh0zX
BIVHr3nRz/MmfMBD8zrjmH7D10EC7/rJEQ/boCo8tbEvwIiAIkrX7jezgN8tkTvfpPgfF62iwwEO
dD/zDpgdvycwgndkIpoS82mrQCn+yulrnRF9LPiFZJozNf7RRdE7g/XvHb0Ik8qo4Me1FNHwGtSb
BVp2NU3KRT80W+lmnCWzn1xenT/8lyzCL+mkvijBFWIsVsH2/UESZglGABpQ4/GdC9rhu8gGFGIp
kvks7q+xlQqiLorOZKIDeGiLbGJqP1hBuMSy4rKkDyMON4JFP2vJBLyWdOxw1CKXhCNbtfe0SkWB
e0Jrjx01o1sRHzJF1KZGO/B6gXUIVW2rItokNcgHgYCgQb5KWkUnqm3Th9iMGLpJckyF5iV7aQjX
hPW8CPQdFwFsUQefw38p2NLnwybM+j2FdYs4RvVTvM8XZmuuAk32xNvnldDqampbrWUOtweUU60x
2IYJSaVtGzFLk6vPsD100PLQU64ziObc6+Vdq3R++BF8Z+SZWK+Aes1x9Lv/Tm3OWKpskqbTGsr2
vznGecrR+7xnC+cxrptA7GrMmCapW3iqEjXW/035ZfA2a9rJY1qLhWsUxyFzjfvvZkOD7kryyftV
5LyaOCoc+TvO9ggNYvnWGksqj8MARX+YNmtK09B0q4aPSGxeO8rnLX//itJ4CW7ZRs2Xycw2NlG3
2LFEwuVISfCtLrgLR+CmyO1REGF99XD1ZvYVAIKS3VMUf55hOamFKTTyxVSogwp/HT6nENKfXJ9W
h08TYmZIPD+CSYRVZYA7xVkrBsE9epi8Ny5jpwRAzX74sKNHkMWRMw3+Xxmu6Nf9BFjUvvuwLiTV
opK6OxDIxfMuogrVEGk8dYxTvWHlUzZryu77TvL+FDgXtLlT3KIeillZzTZ1mhYBfA6/pKG941px
CnPPFhlL/1833IPmsXVHY43LX643UNbZKQ4Eb8DiCIoAwhgCn4f+Xb4IxnwFpgoRGSnf/b2XeoTW
M6Wn2zLAgz6X0xgA9GMD+KPaJppkUAJroOjaKb+32IGH1kaCTx7JjojYCMlVj01WE1auva5QGgvz
bEGNgDHc5c7lESHECV5suOyanUwuVKaMPymunsN/4xatXD2msZmElnUl5aWQ25tPoWx5VO74iipd
dHaG3r47WvdMO7wXXUrfwttAA0N1pTq1uoBHWCNQaSie2AKcDz9BP/6ePm8PLLDAPcSswIS24pNs
HA4bHv1utlAr+aHmipO1hEjfWgrUKtGgs9G/SwLq9w/pzET+EN7+7QdEXCzSGIHuAm7kLbiWkJza
qXXUPJuZUTjMNlOzMALQ2pKR4/jLmfrVwx1TD5DxIS5E5SKtk9nTL/HYhx9giDZkJQYmoyJg/HaY
6EOfxX9hL6sj1Iiie3xP567viuwLGUR8X2bdHuL8zc3O1z6A0ufkpr+cIkgpF94id7hbq5r72MGb
Mz+efCDPBpe/fUcysUzZvefmtIahBTjjczAx9RH9dPrQMGzqtmozsT0vvObEWr03yQ8eW6o2hM9w
Cziy7zJZ37hi2kt/NCQZaGSnuie2IRLN53+7f6AuiyQODacGUkrq/YP/JWAhjUOElJ6ScL4z5SAe
8T5VPCfzm9hF/8Yzliyrv3fMnemmEPGKNSIOUdba8EX7WHfk77nMN09cSt48s/Nb9tslY8iEMIVo
+H470Dh66jsiyL/EI6l2og9eoGMPwjWfANbGO5Li3aQj0bGARCFNX2m7BQk6xeO25Qp0IIvhDosa
aTSfnSGTh478epfsUzztDC5zrctInRgHjJd/VHzkYgeu8G+eV4ye5JfrtvXf0/o6mdu7tFATfreK
8D1bA1aIIZN9TK/W6dWIi5Vqx3u5EIT4SgFSNbmNWL1kF4TKjpHW8IQ57y1G6ZxfvC/EavbFI7ZY
y96SE0zVPALNVyfZXNFbVinyvbTOzUiMt1FVr+K3K9hKRIRdOulX5wOu/rHTgmuQMn1I332Rmw9p
wK+XJFADbcX09Qu9+V/unrfqG+R9cghQkfn38+qmTjC4UElTrYm/n+6JLW6lRrpxDavhybs+2Y/7
0wzH5mJgSl+0zkQ97Uz7ZTH3syEqp9strtNzy1sRbxa4k5BNlkP8oLsXPWl/SOVStFf37tvIHiBy
NcvZkRULvzZlRNE80vF6tdcRu/0OBeBBMpzby3r3OKwtV31hqOJskwoaHKH1oHr5k9TuWoukOx+n
otYpjZQxgy25BDXr/gFqxAxmTwtFstw/nUp9fo3sIuScINbSR8lBBMnhOIGu0AeY/7AAl0Ifrt+v
MgL4S334FLbmnnDAUbvWtfzHPMDEsaUJ97iWdL7V8G3cgpRNsOnGKZ0fVsaVilWQ7e9Ukh7q3w4E
0m9iduLuT86BJPxs5QLioMrNjU5og9jyao1TAiStRxwBOZUHkz0puY3Nf7mH1EPKak7aNgs+no2X
D1zGsMDHflpwkrB/o9+hE5FDu5hCXcJV0f0dKZAFX5jVI+S6GX3PC0Mh/NbeXpJL8y1K4TzzrA1M
onVP8i7G20dVAr/xXaBE4f5e2mXqvNqEm9vHqNykPs0fLnIU8zNQ9z14tYwElOBV6Rxti9xm8BFK
rhKee1AJEhJ0PntulKEU2YZ93jciIwxg6eTFBKOPWe0WgVuNgO1uIXyOh7SmuTDkkApoY40bNZnh
P2xPELajZO3+akso0QYdjveS2c7/yAPcjla/WoP7U0xGdik0htPxOLGp9OVdZxUbdYWz1kP2OHqR
logHL08LEETR9kNb8cdqtdfA/Gp5QMfpsoTHWGRPJbAgzvL1Os+tNdXLp7tjEwB9Clj1X+XfZh40
IBNI0cybHKqg6/SGrMGtC0KwNRR2B+7qIiniNXLiXdZAl8NG9CjND4L1KYB0KEmqMitsTany/WRV
6dnoJiUuJ/mMJXD/vDZcro8LMp1zyD1O3Y2R1jxFmJaZXQecjgagBZoGG4Ds3LBbTy3HG5OB2TO3
hn7sSGM/XFB9X8qxAehs12+Mz4Q9Ekv4pedUDiQedqX05XMzSQmTrVoL3GmoSwGfVKzzmmP4WIvX
r2Uftz4ZCE1y47d/iaCXgmqkKmWuzg8GRurMUarjafXT6OVr1YZTv5JGPBsAnuqQn9B0CPyaDgZB
uh+RTkgfjBSRFJ429qT+0dyNhJkIt9H2v+1ALjTnjtxNDpnRnsHTMvwrq0WKwR+j+66c/2n2AUpU
zao5qt9CQUAR/QlmwBv1JIX+HVHOGCC7pC5tfATWQR+XQvoMJd/mqQpi6imb18S+BVOHGiThIzct
u7l9Bf02Q8N5M1/RwidSs8nJo7m1SZspOZgjgEzbI2BWwnvR3VMxw8WXSj9gY/eJow+dKU9Wg0v/
4Lo+Ah8N9z1OuSmyxj9q/YzljX1jd60vAKK7zDf2OAEpOKIzFnoR9/6rFHV5terHyvoLd8qY3qWW
Y+pO/k4nvqfFOP0HilzcsSTV+HXmxS+5dMsh7tGJhzsmYLHV00kXC1J0bA/XJpunzhVaIH8RjzFd
rhuJJaWDvx12QZnisv/ukKsmHI1Piyvs4nDRI4M7Lz4K/jO8vMsqi9vrUh0o31FutjoN1ifH7ePS
dxpOTHg1ImL0rFGUpFLE9j0rRYpl8h0OmdmkRfpXqxvaoSIoXVUcGlHQKAOfBVP+KrAzylgPgbT4
pmzASFLwbi5y1BwGvcdecNjEymVgSAZ+VX07Xi/1GOyTOEd1z9bJQy8b559uYVTkYTcY1UkfE/4Q
dKLKjGwY+bxHx1bqs1HZSiXQLeNcOMb28IIYivTs+YffeHDZsBxnHMegDcZpU2X4Qsv+/PGs3GMQ
59wBY0k/+lZKs9V6LVxJ0/68WykpuPiaALDWla4G7tnGhj5vegz5O5TwnlxoVfdBRXwFkhU0dmM6
Byf/5RLwMbLMuCGuP0Ge5ilMRTk2BChbPv9Phkyi/lvgzZGJDVqrpS923SlZDMxpUBXUwz+FWGjc
KzvZBtH+VCnnJmfOeLaZAlc/mddn710j8OKD9/PgSaoVL0jfiR9O9GZlijrOWRIM4O5UOB2aPj0V
wkUHfBhVj4WVc+tHnsxqmwwOgTFLSfuFOCh7TusMhkn1gLST9Mf9jHJH3iNfqg6RVZa7wB+auM7o
QGPOewqNX7XzFW4LhlYXH0BwZk6nZsAqY5gDN3DWKTxxfyghUN4Ta3TtXK44WWFhFuoi9YbGP1Em
0YwvkVvdhI6ivqy/ac0E7541SGKj3KaR1zq/BN/MTawITA2dsak3eVsMWZrQhdTK8Hlme1IGJ9J3
aMt9GDxhxSGgNjs05/xOobdswib9Xl6qWbO9CtnYqgWromAtAO7bIBDeXrbXbHQyBThF5fy/tK+P
aMpGtmGEUe6jBDYJimK4cDumfv2tejgqOVPCDGBbHvT3ro+D+jzCNPWGWarTksGLi8Va3LfqEXXz
ak4p6n20s87+sum5nsAHngmrFBIFr7HWJiVROvt4pESCVkUPeiIIV8BT/A8xsbMtlSX3kO7TjzG8
1DrexKhtx0f9afJquESHDOVtZSRpoIHzrh4MqbI+5rTRXNhCPO/ZHNDDl9ePGS2h3NlCv06+h+dH
02mfP/v2PI1nPedijP33zpn7eKK5ZeBBu9TweNePOzZKZFZuag3h12+NXPmCm0vkjkN18xWFjw1S
d17tvKEXCmInuGyCB2qzDFnyJ5uTdwGKVO0YfB4M4JADCmcV8CyKe/pDtsRvt/DeLxXwy1D6HEDL
BYew2rETQy8fH0XuaAh+5CoSIeOBFMKDyHU/xsZWJmKFS/N3D7BIR5uZngsQySSKH2rWrac2Boe+
+2RW5RSfVeQl9Kufw5Wzs6xjTHzqurYg7adbHmS5NLsFc9kd1QzEwZkkFDjTplXKZPOmDkPpuFyK
P1g2nK5KxgqI6ba40CVb5i2XF6ImNP99p2Xv1txF4a5Cg2fQroNSjl2Y3NOgN9bQq2hSbt17bvBs
ctADqtq0qc2RIaZV9aiW3NAbkaNyp/7TyENuhbwdZO8abRI5PKsy3lNh6xXwk8yFVDA4TxOtVMCu
utbkl18FU2bu4bITMESUa6Vqne0/RN09F5lTHWvQDGem+pxzg56L/QRXAzAcXmopb8u06rxKf27X
vMMF7Rj3NjoJQaWwig8lUOl+5Imrsyyr60fwRfyH05VfyDB72MlxQ/DsZFY2Nv8AHD3YUIQXCp0/
VCuU8RWKjS9/i9Z834JttMhoto1uOLnIZ+BdW91KEXpNDjVIhKKUFm3hl8Q49v6XxJnl+Np1zpzv
F1HLnhZXamZTqzIjn/n6Hl7P8MbNcsPKS8LHuU0bQsHavsYl5LH22SRfWFr+XydK+SyPoIsb+FBY
Y6SGIi4csnyastap90SUFQz7EtL8ulfg+jgLSY5YZkp5zoJCXGXLHITQODLAWznRj5bny/JSN45T
twPVg6FeYVxlRdvu+p7Cf4p7oAlYsVR/wysIfYJxMFemCkV/F5AoJgc6xlZ28FFx1HIlmkgYCVei
CoPaYu6GSzm/2FKJKt85bdC8GAUCamYU9CjeLvNYTRt0SJS8+i6nwsFSPgTGZmLJ7UAZrRoA5Ckh
UgLhjs1tJrbIb1/mZ7IXGr/dLzP3itZvk5538up4N7t2NZ6CX3DdYcXfZe8I/m/cjDdmjLgIYVkT
4n0HBaamFxOZBicIlzJh6+Dr0EpBt0jMMIvXOkjIzXJb7am1O1emI5GB174b84swm/HjcunCergk
2d1D+1pQ+lS5qnath+xxvwBCsU2cBXeprfkdAjalgxbpgGul2KMet5CEH5U3ayWj8sr+xAR7vJhy
ru2AHNDQhwOCZLLmp3Kuhrt93p/0Uhq9p4Xo/18kku900+7pg8S1jhCs4x/zSQZLjAxvwHZ2X3uD
Lt/lbB3l5zfpKEO7kYlZvpQhmkrOrfk60jnKQ0B7IgVZakKEWNbVS7PvLoR3d6a9msveOn84++J9
jOsjFuD4zHOI+UZJcTBgRXVCgkpEHO1thFrE5pzDhSGM1xc+bPq1wmVQyr/8Dqj2ThmSvz9oFuQ1
yc8HwFhl6mmcQGDr4mDc6pi4sMa0/Xj45CohfxeqgR3r9ob38ONc2YlMr3eSsu8rwz3aIiYWzgM0
A01uet4OTAt2wrLYU4fOcmgnG+NUVAmxu4qiXlyKXac2zu76R2yswuDLMWVMUMBkWDLh9ibHuHUC
wwy4ojSUGzwwD3I3KsGiMUbu3SwIwqKoXtKe8TrD2H/YBs7Ve+6HtNPjYSdcYyZB/Nzn/HAg9IcZ
8i3rqHuEhNAhUNB+6zCJKhMhu3iAbyIl9BTCgLx53Xm0nkhW7oAsbHuarqKxl6/JR1RCd+BWU9BM
gKJ7Um7u574KriWcTRjLTsdFYTQ/YsbWqRDVvqPCkXjaqO0HnWb9OVeP/mZvLYTAXcs2KswCGcre
qTGAbuV4x1U1vTPsPywJzoOuBgNjkiAXycBIJxA9HG4aDuquFG0KdosnSNGYyh+VxWjjHVEK8NsI
A1ybNzyn8wsvy/Ins4UNgh7g0re5RFTS32k+UJThCXkqDkdQXqW23/IYc3xbirPQL2AwJc3CmRrC
dICI8zcyplk7NlXmwuVebjls83caklFhO2KRe7W2XH5mh/FOmMAE/y2c4DC7nngZkyHmLMF3cXrM
MlVuO4a5vl/nW9zYR/n7nHDynZEjli86p9+DB0GnaeRM2ugfvSTxvwWCUCd51U+auGubuWrSM0Ua
EfgyqNBVF45uFN4F6l9e8YsY0NgC+NUEsYtEtMquygqSJ1QWnvSjZZyS43sj9FOe+dq9HqCjhEY/
x7wt0p2gOzYjwANCTTRNEp3Zx8IMwrRsmc1rLKjh5AedrhyXDsHPXwwKxeKYxARYEAjbZCYXyl7W
sWUFPTF1pcRnbCaWLoYjBNE/EH6I/SjFeIZ9OfpRcqeAHg1nHVbBg1h3GwICG6S7dZ9apm39rnz5
OUKg/nREiXgeS568jJGpxUXowxuYCw+y8Yzb+aJTNilasTLRwZXQ+ZSvNimb7zQkg1k4/84RF8Wo
Nw1p8fMB+oj4drT/MUSRMqzuIXQFzie/lXmaEvuRPZb1vaxmdBFDByPmrh3QyPqUnGXdi1Hw2zZE
No+qZlk138WMj0Y3hXB7NF3KeOApSIifVvHoI+Xx4NAclDsxs6hdc0MGXJCRTcOsyMydVvU+79DA
wqCdZG76Fh4v/K1U1thAAElmurbmzGVKcp1d1B6a/7wSdfGA7DAYrXpCkUU5g6zyw/X5801COUrz
gtazASPzd/HZ2cRFWy/b4CZNxgyNfP2+qse9RZKhOIWcJA4ir8SWiDGLMaIdBUAFaqMM1FiDLNz4
ODmluxzHarOvyEZmhF2d7EJx0uIYYMRx4Mot7bOOPnwTnOoTW+1+mlo41/x+MjvC2xhbg88yIvvR
gPDLelVVJ22Ry/qFjTGmS9FfT81DRvm9kcJxcgpt90/ieuRz9vL6cDXV75tFIYdmkHB+1tuoTp/6
HhJjHqdV3PU6pCnGwoomhDn9p+zbczoxazw6vzoPnxmjXd4zHkHlPnW6LISkvwTkhNUPqKqrwcEk
38Rv+vecFHSRZ8U5Mr2761WYjOOdsak4eb1bXG6PhpiNKTvTqkRLSLt2SgyGAZPSH0v7QrwBtmSM
DspJGHQhTx5/DMpd0BhmvlV4Ym2ifbKRYePPf8UDdo1UJx8sFFFdy0+q+gPHQpo2B6LVfHmgaJvH
7cTp4tq5nLBiWpGNaGrKiHFuHg1fxDGEmuGRrgfq5/0K2I9OE7+G3MSAnRvFyR/LMMpxuefenla0
DjKXC7ZeFZ6aH1/irDp3CHrna7Q0ntYdr7pnT9TIeOE7oZ0+ZaRHjN1nfpbshsmvhECjJP7ouxhA
jFBC0QIkFK0wlbbcNFzNbj2w2gabF7BIQFQTPYaOTRAFTcmJoDwn6/mCnVIo8XIGi5vsdiPNZk5/
BbBAkquOABBgoQVKNHlEcgut+9yjydngnesKx45Z5stuDYHloipGCrKr9G7+oBBsOecsteLUtMVS
7JYT9MztXMMV8liyheBJxPxq75AwTlO/8keXTnqlgiEaantbW2gJ0+a1T30srC/S0X4RTeEgPZC0
IuekmMfYu2GwrA6DdOup/i9WYmaFYan0pLa11ChI9Se6OCRzcdb79+sylHglI4DCzZnQJ9o2AP4R
Sdp1plPz/5ukk2BxPH3Iegn9xr1ZaNpeA/3Tfs18NoMTwqS88xpEHqo7Yz5pW1t0mRArJ+js5ZU9
9mWf/wKLl86uGX70G7aVoixCTFhBTV598L4nyiVDDAuhYaD9vUjnZVTyYmUgUyum9ZXsTpSce0Wk
eLjTas+9II0xasQb02Zy2SBbMF+u1Zeb3Gf1QV54kh5VRR5MEAi/NTLd6YygQfy+dUKYKBkaIoit
d23qSWiT6fvMbNhL6hgaLrVS4l96C6FAIAdan3wcYXpBNo3mqtKjWgV2I1HJ8bSa0bt16kRa3lk+
uRS4DyKI7ww966ULojP0iWeYOOsza+IIlCvDXAsj85cIC8tDpe0TPd9amXTL25l/Wl68P3hLaDvU
aFEhesHtPiY0qdDBANrggtcpGReB0PTAi/IZCGSLg4Psxqmhdtid0xFamBgmpm2KiDY7zD7VhDwQ
kknz+FizeB4cpXKMskWEgzCoo+oQad78OgYyd5pjPe2RddRfEVoRXoqB+W1w35wIb1ht9598iSTF
bLY4ZF3Em6yReBcippNhXwdkbKEyGsSVwj2Qv/bcC80np4gA3Z+c0cY5Uw1OR6MTNoUFYPD8NTLP
+kvT7WsdByHjgWpVhr2t7gdWEgjNGYbutHBgsEnKXAfi9npDgXPnLyhuESE6qbOIsMgbDwRjpPJU
YZJoKfKoXjglQow83encyj7vmaUNcHCN8MQxBQYIdW+qabKQwb7Yuc/MrdsAAH4H0kFwmyC2jKQk
d5i0l/4zFRaVRvDkL6Bz5gnsEbhSrq8FYf8LiVAtU9EKecYrbXSEyeluUs7pW9r5uUSOMG0lfHkB
Et9THeYvuRab51NRPCyYriN1B316CLZ0HBPqYzISPYSKJfi1UZhl5QWSy5ZSGEpj4/SXsNiLZlhH
NFo6oTXikhOX7eHjdLmXYWhPhN8n2PgHuLF/uMTVfPRz/6MoNhw9AocbwgKhtSdOilCQx3blfuAg
a2nEXykVDhdKcOCbByduxc/NdjBQfPGSV3BzpzxB4NzfpomuZvgiOL0u4DoEE32R4S18EU7Ws46w
Jk60Wt9TNwbjbVmRT/KEwOZJTdbqyjrD/nErJoXLha+ih47JarWi3/0izB1nHy4xkzI7imneC/hJ
kVomx1KiHFqA+9mXDKi1QLmuL4tQWepsrctBX8d0BBfhXErGGXqmaOf2ej+SmToWvW08MpfFI85d
wkmRPeR3aHr6VuIR1rJPeDnFPsHkoE7/vaqRTuRnTvjfCp1dB0B/rR5s1j5mwzjiNC+LncGUSSgS
MO/tHI3Nup2CgpyEdceBWFnTTPE1l8823elWo/lTA93HxKNjKRVDgeADou0/GgV/pJyDDSW7fu7F
okW0m0KA49b5gj1NHUxkmKV0NdAznfht8ouWcOzSW7xtLOQ9TBHzncaVBY06y3Kzs2FwgeV4rGbm
IAnhorOjjNlsvMIYqJvDiRPzmQ/4G9xSD2nvTgij86wZPC4fdC/fqYursKncV0rxq5gl88JzIKC0
agAeyW/2+XICOHL2y5E8IuPatXeFnNsAczuDtO2DnUc7mjOKr90yIpIaiMrHMkD/iCxO8jVqc5oF
2kMPQ4NPzmolgn6l85EGSOhRQ6CBGOaJmWtN0lkzKb09ws6swSSQuG8A+c7H21a22KZ48dXzyL94
I1w8hRalJPmu1ZsKzQKnjAtkr8Yr3fhOxVE/yfDOdrixs9eVCPwW4jz86Cb+HtWASppXyk4UhokM
vV8+C9tZP7B/F5y7mVfSsCe7BkaLw4srSuadQDRUrzxf4XKi2HrKTp5A6cBym0/fMFZbtCATerzA
ikHr6p5mu2h3bRp+gY8X+BULLebUzYshWBZ8siKhdvy3KWoIRTIH9G5VLSUCKdjx/VIdZgEYpUBt
rVbKFEjMxhxAr6wc6MTCCjqtOzguyzPbdiBT1R5POi3gIdak/DD2i7vO0NwZikb9guAKYe+F3rdb
IoGNnxTtu6hHTL0766xjXRyeIFohtsfzaipuV6zvmxg9rW784wWppPwVv7FOr/glyM8kcIw8Scdz
jDpPOibpzQf6LD7ASNiWZVpfbxTwjpiZi+OIRDHi9VmzsISzrq6s1aSOAQtIDuOtTnzcgsPd00wm
4cnpVronUQmV922S+nXJmrUQ+rGfzgv4xDJseJGcM7OmiU4DYflv9vA65MwPewfV/ho8U17b05Sc
83ZBD7ysHsN6JtupcTAnbqaa6lszQNhzTTRh+Ppx2beRg9m5tsvlcltpGXxK2E/9gvnaznQmMi8i
E4aiAJ6kjNLwoaMXYttmAhDxn/U3bPXcmlA1lklAPptbia2vSBsyIjJM4siqppH/2jiQHb7NJrSG
MoBhvGsT4RE2OCrxqxiux+RRiAQE3a1q4xfznzBK0gd25AkpzIEBH4b6KDWJXm8XT9rscnH45ui+
vOv1/Z8VhbGbssp/eYuy4MuEVLiMbZk4PI/QvCvGRQ6Lt+2UUimit/0ulLFyL155z3dQKpuzaFGZ
q0e/lgaRktiOAvvwjR6iQSV3hr+MjFgiJmaza1Kl0cjZpiklutR1CmE670QB0Fhy0Y2AuuGPlnsJ
EZYl6XGPSMCrDrBq0hZdFE4zucCd0eJGTIwEGRSuTpsKJDtkKfYOlD2gm0zTkITCGN/5K9ZT2/Vo
nczxDeKxmxvKwkT/oMDmbu+KMI2uLSLbM+3JKn9wOGM56no7OLvXwDhN1PK8cRtkkzsTm/JCIciP
Ku5HeqWqA5CCq9wPs0gmHPGWdbPQ6UN6q4R/tdi5KZsbTQSqP78IHIAclFzFFX0pSZKXDgR8RCCG
qAep8pCUGy55a+0BcyStYy0QGoapR+Y53kyUZGLlHHIfeEMSnQVMXt6gbSWjtfHOe6vvhGxaXIfS
vVyOh+g32Q4ozmEW/lajGHn5wRbKaJTALUh1tae8/rxEg8aP92YtTr0JfZhV1CYlFRoSWLndVHo5
9L1+KlnRTNupAMVrexAIxOBuPpNT3994aYd1nmRXj6/r1SoKqU259o/JYoYbT5vCF8g/q6YtQiWD
2VLzOer3Pya0RhvprdT+qVfDTSZmB0D/+4x6sHylGGWXsDj3C1S9OOUxGEInPEyEw9zXJXbuwL1b
5sgSCrOoLRanU+Ta9RgR7eSuDucCYU+MqpOySu9RFpluoWiyqLJEXbC7a8lJ4hgYMMa7vokOZKUI
X/qOKIzvY43s7XC4UUl4INx74vz3gZJxsLlV+0yPKhXefFqaXFvLz0MZi8+t9yjD+eAUfVxhbB6r
2wVYgto2p5MwV7rui1n+mWy/Kkwm2GIosc52GsO/Zre9zddXge2ugdpvfuCBrTBYe739Mjhmj9VO
FzR/XMYnwb6piZScErxKBsoMB5oQhcdZab0ImqaICP7pMyfR8Wi3AXLRq233jLw31lnY19zFxTYW
y8ntrCtPLu9yiD0tHBMMkXlanrupIyD7lw+bt3VMIYpsbyYNP/XjijRxWislP0KROU1yKisMHWHn
Gk3QEfUKqRtcghFAvOTdAKAkBFRaI/yTMJflpH5t3s6W67KG1nczdYt2b+Rpn+yJrDE6/yEw8wfJ
7aKCRg6HpmlCMePw6Gi/r1ZjYL9rE2s5BEA/D7m/KUbnEJ1T9vxem7Mx4aiU7plkLsmCS7BV6YgW
/URokNsuCNHnfYTpVaNMwrU00g99aspCZytPapoutpM0rAd9kI5HeEaw19ZtrpoE/pxiqF0Iaybm
I66Jzj8zNUQJt4trKpW3Z+QjTVda0MKnUbtULAHTQKaanRHuHEVMBPdghc1KwCWepeENzXnBSEWT
B6dkeJJlkOVJBsPlds5naWE5UOB7KDe0Ihhl7sCyLLpCIUpgqeYEpByYA6JdbMUOPPSJptTu3lhg
+BFn/ezvL1AL+CT6+w9zZWCw7u/13XAYDUI51FKoSunB7hlmHuFtXtV2R57/GjEbfd3b9hj+7L9p
jgb7EBnriTUE5gxow9Zhulc3Uy17l7y88VEZa7OHvWgyPoqufnG7svBcYjmBxIhkii3uFPBoHmrE
+EoI8UiXafgI204FEKAjezpKtYt3yb/E1bTWtI43E8abYGopWRxaim6WHcx4dFwD2J9HMYXvrErI
SlaVPZbrvrVmEKNWeNW76mi6r9eT0qF7tSNBc3KOqs7OZ+DZhOtunqDabMpdxx9sKINZKv5WX7UW
KPktBLeFW4RNkMIPj8mNomfZ1K/dzdFmzCSQqJSRWCFZI+JIi4z95C8SaanZgA275FMEUNLG19kL
b87R0A4dwwbOEzbf4njqNtc3GUUZULeQJJN7GVHQIYwo0eBVn1Uc+flkU6Lzyvi1OTLnF0i6hqiu
eJ1rz2dHVbMSAZW09bgVtKtt3D7v9o5fF8FoSHumsanyLp0bG6tHyAssaJmSkX+Xj9CK5AH5OBHK
MtFa3DghVb2zLElWBaCsf0v3K/9ZJJ0KkvEfeN0vc5gZ7Mr4r+98FLsqAEvLXOACRGsQkwKURiJ0
F+BWafeSKZ5avhyuTHOuRB2A4+KhT7oaDJde373yKrUTqFYKc6PEUKGMwnPaS9cBvp43udUB3731
OMGzpBL2aD87S99GjRQcJ6oKqE/flOvA0f3mNCC0AdmIHnEIKDJxNBX9Dz6ozwbAuGR82LPscQvt
7sX9w3GxWX4fTv2w19/l0tZyPONliyrKV33rXHuR2X/4Vboq57cOH+0SeKo1G0Q7kXWygRVXJAQm
GQ2lFHPxqM3CI4caUo3rhkzTtp6N8A/UG+FwHCDvZoYPIuiu1T4uLPaTLCBN3o5vxH/W0kXIaaoy
7Vbi+qjgl6IaW7u5RypESj5BikUa+kL4nha9Fe1BwnncdGcGeZu0EI9Tgoor7ORB+tAM+Dw4aGK/
TGrBHo0topfGEDno50237zZtGoRzQcBRdf80rX40KA6+v5JGDwQjap32W8bmq5OXvHD+btobwFmh
6439vWthOBvu5F3GMATf6FNfbV9RPg6afkFT+6N4PVxFU4BetvtpK20KnNNRvfpcbV6f+Sun4TcV
bo08ygW+7iezb1aqHNRrUY4bLhcMH/83rDVbfDZ/yLiAHPa9/8JuWQIfcsFzex6S4wmjk74j+61j
JlZ4l35mHqV9Yr/2frr1alXQbaNnnlYyvZNKR81gAL2gqFtB43Mf4z5nLDXlb+smwTZLPTCGxj5+
uHzwn+wKEUIx53lbyDCyAY9Dl2CsKDDKz53hlFTFqnTTFQb8X3E0/kXwETjSPlFeVgSZSDUzJKRn
fG8ib/3js/9JsKVgtqsKXIZ6OQ2hMtYggOUM8KCT4P520PFbcfTupVcX7KxfxjGmY6wYpTK2EEVN
cYEYL7DcuSmDwGWjy6kEP9CYrafUxbzsVdeIsCKxI+QueUnfhOaSQWlczG2LXlhKLdrP8Kejmwd7
ShW7TuY3vdFL9aOrvLQmDq2MuNwTnwPZgliewkRwJ8e+EmjzLoZaVdrKlqq2so2ABAkIiuwqAHzp
7XwkhhRsGdfKMK+swJ8xgUZ92ynDlZEhLV+uY0+29G3TMdYAcwzNY+yMgpd1S6eF50dPusJzJcaM
cZyoXlndZJ3W39dqaTUE257hBciUkHUAVbM8eA6nBdvIjPfqdMtmPvwmoUc2xT1zdyfaYA77hf+R
YultqwWpqK4ydD995OfnVxzGjWlCfPqKFe57Xcz0MpXsdDplK+OVMLFOWRqjIVvMKt2st2yO0sYF
RxjiV+Cu0OplELLrC4/GIgmSFoJoQ19sxqTq9hJJxvTjFlJsW0Ba+nT0pO8aztc4Td+2mR0ShTpH
qvCoB+gg6XBeNOK0Zfzq+fJkvNLsecXa6YNYRog7qq5Fn/ArjDbmdQwBHVULStBWvvyHsogNrhcJ
YWSaVidB/i8VqyD2U/03mVPDAj32ww/htfG4af/i6UtrEcZFpwbnBseS17VBnQfJzYRX6B/95AcK
SG1o8r8Nykd8V3ka2q8ZeKCyvCEr8uoWP/waDu0PO8SNd3Rkno8CvA9bu34HuvgW1kBNIRrnUE5u
tBrDQbJ52uj8GVYq70otsA2kOhHZgIFC9N0PBgb/qpblBZ6v/fzOzdL8mFaU/mgLwHITP7Oyy4fQ
0Nb4s4uS9byvL5pAjV7gB4TLQyLf8VvZYPI/KrSzcAGAMpxqnrkVctTL7bDQBQvAfl5P2MmO47M8
MQRmy4KbfSSCxqKZRj6qu1MG7rEIXYobAjlrooF7akYWd0Sk/zXdIpJN7X/eXlDivuZWeTDRvQNx
+qicBjlOlkzjnOgN/I89TevLp7y/9Kb3yVW5dz1jFgLeb5h1tvo5PC8UMB089VdZ1cj0A6eQbsaq
Mnw80bmBrwaU0V3bOdtQAzijRLGsrbQ38IErXFzPqfK6THpkYqrhX9V3HBadMdUDHotfopM7FuPG
T0sQ5WUy6eJmTo87luiAYyGMl6kfhe/AuNlBcjPEZ1LxDCIR25uqFnkpUbLf8srSxVl4CTnJy/co
H56UoExBaEgs/JY4m2+fPNMkEh9Y0k7PSPhe1knnmc8Pq4RqE5KJHjNqYTXICXxx60ZxLhu842IM
vWQQefT54gPnebnApUI2anS2A9OFSRxDpxpeJ50wVBHytVOXot+x7k5qQxep6ITGC4SfGhKAYyqY
G7F1OAxThjFmHFFS9ymi5LNF61bUUzbUIRaFYHA67ADjSU4CmVOSHxXzchSw87jVpeZ6Vue8XbXR
QvjQsSKDRNKfZMibVl15wbpZR+3cxS0tglV6LSEY3o4ueaRJ/YafIx2BByBVXHNiWbpLbP72j67e
x7tzAohnnU0hPh1J1dn77CLggSy4XiYPXBSy5MfevNT2AU5kOfZlwsx5TXZi8ysmj82GaOJ77e7K
2SuM39jG709HbLBKWFwZBgGYgjPVq0MJCGncwYonmsGskQa/8Z0qRWpi65JtIzJOVn7GR4Xl++rp
A7nCK9vwRQwGT1/bZ4pxORTakH+zxmI3Cg3320K0n7nuQMghjcn4ev1H6YbbWZsGHidFim8Ang+e
B9vfU5erW67ylUeICBr9riwsTleO3vEIrowWHPVqM5EdlAaYb0lZK8RkyvTmSXG4+NSpmziGFhi/
1ep7BMUeFvFUAbGNRDvkcVwrfIyfVcOf4OTx3ZCudKzt4k+LimD80V2DugMX9d99ApL4Bpv1H3Iy
cf43w3jTphh8SoXxNegAbCa0wRdAaevoJAGbsVVvmqzvSOmt2vtGem1/iCOM3EsgOH2Yeaofy/Tt
zADyOQ/4NJra+Ukj/NF9l/yklkk2drSLt6JLS0/XL50hIqOfIpyAqXPjDrJPyzc6KW3MsphLIVMx
ZII32I2chqH2fiP5gxHmfxwRMR+CHqvXEBA4564hpKYCFYhZvqXIkwgephGLpVxoUgPo2dkBTnsd
pC5zA0iI23F2Vlrt8vTPWgzjsydBnDW4HduTHLgTCP+JNo425q4JufMu03zx8NNRHriPr79tLanJ
nc14QkXXCgnFgZfO2ukdu2EqBRXU1R0EO/wtRXpXOxO2zbIZQUcVkdeDs7i4UgnrvzlirRN1PLgr
JnTaleUGzEZ6ZMPIeanInRhe4+4G9NLivXKhsVRsFQow3nFz51ofNHDBoq6X40/YYXpJUTq1eSsz
TulXcnm2p76+ZSgEivXdxBHMW+/k78S6KX9aTPn49wCqXd6F8fJ1g2JYP61sP+XTT2YWxZX9o0Tv
PW6pFLSrbWPqU4v11HlvMQFR7/XJehQDa+4tVjUiHbJ/6SeZbhxp9yQf3aaQM0Bt/Xr6i4TfkVbu
clBOf29RF7kprW/4ed8amHyEtU7YSUthHiurvhyIRWa2hFPJl6LFDD3iDAWFYfaxljTwdrvVZd00
J4Frf1vM1/t8wfyw4p/PAvFfSNef1M2/9E6H8JOHHl3BTk1NdxcIE6r+6rbJiohz9fofQelDKqBQ
v9kxdIfq6M/tderZLZIUvvpL8fkKH3wMQwXgKVEbPOkdZ34kIejd/PFyBrx5rDoWFgMFG3+fS9vS
d69JwJPbZVnIEHrEpKXi6SwQwVWcesbyfKhXkVpi+i4k3DrnqtPEN5T0XbYjUWvbkOSTm718CQZB
OOYbeD017NgcBTDMZInMceAnUWncJ5ceA7uHbpFdTKaWutNlDR+yRQ3q453GOgvksKVWFqAIW8E0
3Y6GQP5xkflRNSXTnT8vwgbqAXjc3IuwJpiE/MANOhBVwTZ5S6supy5jk0g7ME4ONBKY0fEEBqjA
S9Mwbra2/EME0Sj/gvw8cMBlJlTr7rd8JO5tE6XTrNhqE4KUTMqpxAdwPkJqzoSrBMQmvr6L+Tkz
H8AMHR6BpiKDzqB7Po8DE/NR0dvasA+yKam15H2nz/kjt5Oir8B2mUhgwZ8DwrgM2yONMpf+JfNU
V3MxWxe5YKk3PMcUJd+XjUMijoHK+kZJzlQ5KDvZRYvYb2Z8tNBuWdnaGpP7yWQ420o65WnZ2LXL
ybkMrW4qu774V9WKl42WRlYAMKcpYBCl2/gnvnJw6Ft8+rvgvdLTVZXJs9ByXDKEHUfyD2eRway5
5pmBwQ/OPC5EVWu7cMx4naeEQceliP0KEnuqT5Y9SC6erhl/PStWHJsOezN58sX5bAio7tURoJZF
jOQ0veyrLVk5mCVtKFKUC1D9x+kYOZZQAjcYyIW41YyocZm7wF11qdOm+kobGgQ7UUzobTc1mF67
BP1N2qshPTyb5lxCJbjkg8wuiwvXtbw1PKrnu/f9VkYlVZqkcqWb1TaCPJz0Oed/iN/1Z5DY9TCU
mdw7TrOzGTPVFPQE+fR6UGPD3P5nHk2e3EOnWUkfO9OvWpcBi1XkFT4WLF1ZZS183iDX9ZZ47wo6
eZDjgzLd+HtP7Fbqw/buqtotRxXVIQrZmW/oe1Th4LM9rPM92m24NBJ2vvYpOvYee8mtyMWKhXQ7
8xYTFLAvfm+6KQ4mrX7jUZGbqXZ4IFqK36xDCZ//qCTIKjq/9Czlz68+Fkjo12KI8vzk+VQU4BsS
ZpsUdMbzQ+eEUYc2WNX2qZrA2WDkIsGbTsSDzHoUp2Zfd+VjveBFtlrlvscGMD/v41x9JOoMd/gz
/RexT0YOiwANUmJgNn+rNEPKz0UtH9BT4KDonnJeRI/AQXQYdgBjPFMEr2C9QmzhvbR5a3GG7YMp
tuxnu06FO7Sey8X6mbChEqD7s7+ZVwIhKD5JnQ+SV/4w35KJ7oRJtWh1rf1TfNXXLN94HaCEpvW8
23kkIpiRveuKJUBvLdFlzNR3rrVYwXwaNogAWaY8bI7WPortqH5gaVIyhzX+ypGoYi3nkjdbh0JL
w6cIj08XgoDgDEOirBAv3/9jCx6WQoyPxW2LUEq8TG+qGV5zvH5W1I/dYR1NzRN3ffzwSh8JxK2r
JcFlG8ad2aKnrl1VImrYaE8Bkui2ZIRh1M0ALogFk/34hizcWmvocekCrf5wziIT6K1L4I5dMCJT
ZiR6EzG2FvQY5ksBSqTu0nHnSiphAFd1VLrcsX+aGkzor6rrI/ZVuDYdYZRnoKk+NMiYoPqwItnZ
XUfEtLHHTYK0PiotC740WwcUxg6iTtRJhuWclXXQBItvKEHAdwWH/INxf30qJKkhnxUjBDqB6kwL
Z11WWOcIALkwvLRqvkNaMopK2guueq6h/lhXnXE18YXn1CcnKJMZNWP6VM7ORhAACNaaR0tTtBqR
og1Mc6vv928qcaa/+ucxZ6nV3t/Spe0j8wflkdxveJjpbP0OU0Wha52IkofNibN3rP5D42v9Oidi
tVnLxgU9V4QDVW0LpjjUwkO3E5WmMPwgoP8NlfaXLlFvd2ZYXHjGxlPGsVKfEQOrU2PGMKGm8GbO
S65drl4lrIaVDoszbbpb6sRUZd4S63GDdesqGu5plVaVzYBhGX5+6MJr2pS4UdcXRZTi8QOuNrvs
dVE0JVKpajVKPB1xfpruIm/XccI0LkvqOmQWaTBy20XlH25t6A6ZrxozncRMGDQ8Oh2IMCNeog5j
KVLtv4RHRkjSdHeSSujNly4QcgYaNCkwDvV4jT3lXU4B0jtDuWiXqCB5TaAuQ1U6PngvHKyH/zNv
YK8DvxpDzMMglVqdZhIBrI660FahVH0qxsWyIJl7Ex2VgWPUwjD5mzZLj0XoSFrwOHj+iffv+Xbl
YzSCl3yZfxlwJkm7xXSQsR3TYo3IdikZvqU/alAVD7w7IZFQgx80wTW7aJLBwo1CmlvZmvcz7UXH
CW9HpTXfdrqiUvoIPNJk8kqRN0Axiw2D0B4qwcaiuY5l5u3aQ+yuWRSzqFEEdqc+b7PNQ48DWShF
hERA3xXn3073tWWrna3xgZRVIsJ60E3djBca3xOpwOQBsKO/jNu3Zmu4QAqlkNzGxeWmLp2KCVdC
Iz+G3jR+FdgIdMgvI9MMJ5vne8YGXy4FwGsAmBqqhnae3rUd6tVD8ywTxFiBZk9EaGCI393DE+B4
QkzvIesmPZFpZBPwAQGN7zZf7MRep05KvAy1mkyGkdIw1M1xCV03+pfk08jb+V7mpUoE+uo3oVMC
5jiSw93pvh5tA0l9P239WU41FaD05AjRt2vEJxprzLT2NdYqt0sxvKmMIXrEqXz0OOWIIxzUrGnE
dGnF/7/svcHMxQBVo9PsXo9ZoK3Mx6LYBxFT7nOhHJ6oxaqj9t39lBXewnEspyHArR9zAcsDZVCz
B1aGbZl16ePMAcrtEsnljUbUD5IMYntzRaFq+5VSGt5sU6Sbu5CNF4+V8CvlNnxSulKtOCFZhmg1
QyDnIU+ZyTEpuhertvtEBUtPpWMSPwBsGO/GVnZIWZ+aG6i4ZO3xjPIWfY5kTK/sZFMwfzy8nLIl
Ly63htz5gsMPH0+UDh02c++bwLPogyjm1qYg0bOq9+GvIhbS3OxqNuYEQXvv19eozye5GCI/XSnF
9hMvPlY4T77ZbJGDUQV440/Avw2CiUrToR6eg7CFrlm6yzTnzhmg6IxSDq6WzhIjd46KNFjiPrp2
Ib+BClXsdAmgjGnRUnuJktqMTO2hBcJGp//sqI+LzVdyQyHbXW+cdsGHZzlf0P58tiZY41avDe4E
BKioimGaKizNzNFMNbCa4tMxwIVrZyDi652opUPFwSNSDo16N3NI1crGV9vjPnCzia/cg7mpLVJp
BH4TSlvZxFcVTwMgvAbFRF+YFtkQlvj/UMvx5SCqCeIHIIA8VxDiAIKOc2EFPSMRqTwJZCIk4rlh
mwWnuTkFLJRC9azvgNjlLVsyyW6Y+cKn3FvCbTeaUJb3GlI3V/4WttR+wLuCDujxrd3brdu+1i6T
Wojeys/ilI+vaO/OL38nLyWEXa7mec7GfNFHcfIiRVHNHTMJknndAWXm7Z37ovG4c5kphKsk+Pvg
kK3TGmrUR1PGNkw7G/Y7Z8o61cBhXXolL84S6DNMtzUYCVti92MP3ex7Gqn/zs09kQ4U1mxFmElT
tdfZ3hixhz5vvJbpPtSAnLsxZEK4qDd/B/Fvw+wjWBogavDwuyuY6hsq73m3IMyHi3OgZ6tC52Hx
XQ+ItoBYLOxqTYwanayRXXcPwmE9GupsLJlTYF0K9sIv1ofb/b+KHgWXNtKPmUEQLspzd9v1jYqO
VZoV4+DamIzS1/RP6Aobgvrk2Bsyz9H8h3pm1T5GXOPuBK40hvNGokAnTGzwPqMqPVbyCWNZZkNh
a+w0sGkjlwBm5ZmTRitF5qKY70SJE40ElxyajCjFMPrHgixNfb67q/Qlfo4dZIog9CZOjcjIXByC
qH29zZqPNSCe4Af3436MCxBNMokP/TGnnEpTfLDrQ1+DH/b3ObqN7f2KOw4ruJOMBKqwXwetop2W
mGYqKpAV5Yl6a2rA0o5BKpLFcQsgGPUu4L2DhW+xLwsEh0K1lHC5Myt4Ilp3Ny060l3fRalnLhQ+
SID2LAKsz4JKcq51Cmb7XctDShaz4DlPFEeZ8lkpyntwuBvJrjXSSUeQQrZCG1wgmEMjBXE9vWG4
78bt7lHghdskPN+xcor8lLiFAkRgSzxG/C4w+l5n9mRle35B0P7fLdSJjLyulSUCze3fF6m2kkUc
DZPWklMXV06s4DpA7O74N51knHdn8z7CoVY5u9jo/qKaS6MPx0cZz57/PeJz63kZDTu6Ggcv9Adg
mdSFWtKWGcTLyUyOvMZ148S0E0IK8ix2rsYYN5C2y+Swa/9ceOsPpvpsSsWMSy4j3OlLzGStlE1S
7lykWSo1AJzCtK4OYLuPIf8rybokgvVOTxTHcWW5mpcW7gBZciO/DGWB92W8gEdFfVBoRklV4Gj5
2Um/qfyQaCNzCY68SZ6b8Ve0BxSV8pGk+6U2ctx2RNVr+A6wNzIczXwr3TJoEiLUEPdcnLUX44ka
Rjra+MZAMOZb6AXubcq5hEYYQd4IH+Gkhws3q/YrPGGpU7e9pBzHdGCCNseP/HSSA4W3CCs2BoCl
MBeCRx2whSJS0v6zWRMyE65L2xeILzG5wFV/I6T3qeiW8+cFqYyg2Mgx3TY55b/R0yaxqDOuin9i
8z0mETcFxRJypdhFWzXJao5AoRUkRwiBDf5wRzqESz4y+VH3IXBaUxefYbbmiIAMNNfpu8MzPo43
5JEaO1YciVJKV54PdTV9lka6txg8dDMA55fHqj8nGMPzlKizkYEnvA7mNQtLYtNeaLGgX3AhEmAn
7v8AUPyqPkExffGMKEgRD1cbxRox7IMfkFN0sr+G/iHkkByE+9oFEC9l6R1DdBYpIP2EQNMYH1lB
x4lwM5ACopcxder+n3x0bBYJP1GIR90CPBvN4drrsoyaT+Yi//XnezknqIzRBel7gXEKJZOCO/2V
1rhjboct8iIu2OTQETuQNcLgK696+ET+LfD5MfkGfT2F82l+4MiylOEiPCxs79DXbW5Uz86Cfi57
XLJbQ1wGAVQNTp3g7xBJp1qxHhqM743gXZWLA/l4MAuid4lbBWBuooNGgTnzISSna4tZess8nc1o
QribrVUE25k4K71096m9WRw2YMhRzMDpEnFVgfQmwwvPj0Bsb9yKAPn40Gn6IN0jD7/kz/muJHhJ
ak82OwzCv7vRBQ1a3HR+ZtlQhHg8sqGdcAqYdjMWojzNrrY4z4gX7PTj6b4RbM1M9kzxmkANhf9B
0KgbGxhWvjRzC3tNel5LaNGkjcBUc/ZDR19nG5EiIxKzcbm+Hk2hY1ywW7v6KDFndhiJke7jIbcp
9/AaH5tjUuAxLIRty7/sU6Y2pe4GI39Rr5bIjr0kKHj5wN1HS4a0OcMWWNpZz3WZ5Dvk4q1s/N33
UMsQ3MohHaTDu97r+mFIebaPOfRdITOLNqpPHl/Arzx1o7ra/Tf2Ap/FbX5qUbVq3pGf2+kY/sf8
YsDxfTkfgnb2N5Tl9YrBV8V8B80A9y4wSdlquExyKJZNd9o9YRs6lfTsJJOrJQ5Euvf8XwIgkOv5
FxnLjiXLY5KTrv2PLd8bpLXEnTDN3PfEsE8lX4kO4xVzLlWN0RucjCdv5hmJLz30QvuD1PAM20wn
Odo5KpZjamRrjcdlD35ONTbQicrrv2P0fiJSiGRXowlKDZuJhLJJ/sGhIIwMrzg4oLL1gKAxx5M8
45rvE/GodQB9PlJ56jZHKnPeBodJOIDAErtghFf2DEHAO1lZXpqQXgJ5JGGlD5C7EDLF3kHrR1Q4
f18TJAb6Ebi13KYJK1/2NGW2VGswv/Q8WGdRjEXW/NJfojAt950S+rbp+fq4SWcv48QGEQbVlIOn
mgxlp/mWsXSaPwQeJughSAMCmBV6acYMdyJ1Abzx8TUq2+obYMaM+l+VBNJBjYEvD4lgPi7TBzJ8
Ozlw6y3GNoYWSM9iVHfB3jog1ABo598+j1fj6WSH8MKzioYaLedRGSYAUsh6q0itLtf+2Rx5k+L5
QQRYV9imz0SlSNjoE0jwZqZ0jBWQoSL2fj6bqUWGyIeaiQTq6+2/J8l/Zwho+H1wh7MuL2ULjqlY
mLKcuqQAcPwyJKOErpLHOXfDO3L3CAqQH2nhSKdgT7UPa7I/yayed3S3u2Junb2mk/b6VkULvtiT
uIF+Pq+98Wk7MmEvXOBe8gS4RyWxekNj8gEtVmc0EkI34IyjNi+8+222ylfqLRhVDQTJoX8m95aw
tXP3/RrliyUnSftRpGpndnCnJWLhXkf9R5Adkf1OhHZkeImSesjD4LOvBvzqfO8dJRIZEHPb+yaE
D+6rup8RE4g3gTl7p+YCqs0Db8eye1cPR98J2ICswaE3s0il5PrvEe5/PVdf1OIcgzfPaY4uibFe
zQyIZcQbNnBes5HFMC6dC74hZuYulvmAgPlMqiZ0Ff3BLqzPox2vAUGHaxXepp0YY2el1O/qyqRH
vDyHaUKN2pj57zA5mT7JmZVUQtePOkybCMX2GdwBHZhs4xpmkVV7Bpko7/xb5IjYX4U+TMaM+u3Y
7IAmhmcyxIhaZ44j2jNL+8pZeiio3oDtvE7A4hkZrxVr8TQ8VjJESD/RiC5p0DUreQlw8M72NrEO
PvpSlRjVaV2nB56mDb/q30y38bQMKZ+/kGwpEawkniMvwGEi27FCD50zwbIcvg6mlpLjlD3sWrxF
yBlimKzhQ25xc8SApEkLgvdnF1mWoXgr1Codhss8qnfz9JYUsPeniKTj3uUn9GcL7j0sfY/Tp/0y
NVSXB6Uqo6PAX3+J7RxkBsVmjLrxTxejftxWEmfnyyUH6JJ7AxyHoUSawhDqat7ngbPCYcwXOOBb
9ripG8d188dPmhCS7vG/F0u+62g9uhD6pFCFvoexXf5FS42FVHIvekVVooPo6/gOXIMFUwBMWv/D
P2P4vqZ7QtY4CKeYvi52ZJgHivCCiYdtsFy/5I8MDQ8cHLwSdy5072GbToTeR/e/mDP4xL9eJCzI
uL0oIDLH7xAns7Wm2emk6kLAAWENuRHGzgDqOd1xJNNNKyK6Rie0E3LPVbMWbue2knaU8GwUz4qb
KgQh+bOvfc9eByGCOt/MvUtf8eI2zxXOUoH4Pi/Ryli23FyH2UjDWDKBACqy1WW/vGx7Q9ryFwbI
cdUzKAcqoLQh9G000A0kppUo0Sz8P0numP9NDCkPNc1ncTBsXRsd5VcBMRAdoZonmNLEaJ81mf2r
KA4WNsgphWUf9TMRybMebuu3lZU+q4knxnERDIZMpEZwMsBVJqV0X2LCseolD0zBDKvzXcVoos2H
v9oItpVNrXonnBDxLmQLXYRuXJ6iDDN0K5HtzIFZdtAo4ZiNLGFRsxSDi4cEYXb+Aam+C01xwhCN
jbhwPsWGIPLc4X1CA7pMVdyR7DFIRiZUX21GLSfXI8g1lZLsUQGaDHNyW28AHhZnTlpw2FQuY7NO
RkspMQo7eqQHtJVn60ebHLC2lUFKbIheueT1kM/GAZSqocnWO3zyXY2BsWs7NYI4HdRg92hjj4wm
o/P/jaON2gHjPuFMHhbwd5E//b/Uil3tQqGAnhpHN/cu2sLxOCZpz5HO9xhodeqabgByp37bc4S8
fNfWN5W/2JDZ6Ic4+7M/LtoeropYr0bPxMZN8Utda/DXPqDBX+tsPuvtlx1gce13foBdT+g7EXQW
hTlVoRuXtFGfyQGEbVY6uCKWVl6tvL1nibj2hnbZyND//vI1nm8ABM0SET9yFPKAtUIl0Dl12NmX
pAoaSc2YfBSHsAJ8sOin/Foky6pJ6AtazAUIVKV8vydDvC8WDnZEupGS20U5gT0SZlxS2qnNOlGd
5Kh0eBJVci30Oc/U696ij3YM5K9o45EKHBaWOZKQ2fICNXMlDkdk6VNLx2VRJMSzok6dZ4JzPxdA
cJbRLp7NhFMU4WVm0Q8NgMVL8CKLFOtepQas36aYanQERV3j8yHov3Iu3gA2OrxqIhZZoidAFyaG
nFJaHUmAjAzkHV7O6kXufLoGlcVLLkBLTW/DjxBRXkZW3QWia0llAuSy87Y7a0uPqZxVKiTaVHGj
PfOAor4YKzQ7RB7tN70Dl5s2lkTj1b/NN2h05zUQ4RqevgTIfgr9OlGrddOtP9Tk0lgTerOmKUxz
RRFEKOFwVQUptSLqKagUpwlp/PCqowzndhq+EWy/4dZtbrAXx8Br9q4UsoVoWp4QNlyEh4WHZZEa
6gWgaL3dfmLsRaFBMi9etL24eDqM/D2lLsSUd2zMPMRJb+ANG9rrExsR8Wz3oT/1fY59S/0lgwu+
A3JwcbCnKOVVjhyuymqqg1jTb2bl3fcle7rnzTQRDNhDkn4epNPt7aaHTNdcRdd1EKMwP7UlKrIq
mNnzZTrtFuTIzqjIubnsPv0qU0WyLBFGIfqC492rNIvGch4z9r2zbbLj9s8ssfudqa6BmDHY/e6z
Zzh+HVAyfojcYI3rqlF/19TCFGXYVB8pnLAHBPitMpO6Y3P39a+uNKLYtJnnPSuX6E0KaWzJvU40
JOoGaguALAK+0XIjZtO0LepoUmAFjXUyKpvLH/wbrNwKZbxX/4ED+YKjOXOe1P4hTdNbpy4JIObQ
TwLYneXAYR6HVXX5nUtCK0F8YDWZl7FInSD+bWSlizJvlosQcwIiyU8tZ/2U0NS8aGXkYBNxcGv4
KQGiPGwCWILnRNTBLX1Va71BP9Bzm0yKZgCGWfRHIirxVgR8Bj4ohuPGLGlP2OgTVQ1PotlcTzoN
jTlFvC0TD6SkzZdaIZDtRHkr5nxzPI7C7LiKbk/QZtgDzVUfqHNI+AVA+Vg1bF0z0XoJw4SZ/4Kv
QZN8nrGZp2/eV+DwemisjpiR/gT74eFWCJMEhai2hS/9WW3bKbTUAQd/vwLDJSXVeSkg4v9CbB80
Q1UkFFjVzPjjJTFXjpwxh/KIRW8MxDGt2V8nmBpFDk7SrHhZKsnfjyTrs55l//7d9QC9Dw9viZOn
HIWsNgap4flFzAE1WW+WczD3QTlfrWwnvyuJ1dmxWWUgnj5htR5lydu4j4TNHMpa1XpUd1xFb3Qi
ELSKe2K+POr2LAub4UiXUEFdReV3fJHKfJGaDED5kX+NQjgmpcuXhi9RoDoNjz9zuSs0MPyJa1tL
1m5f1OwpJV6HKQJLcb+ctApF65vcXdXjbHmJKL49unaao+VMirMRGWBchLm2QcWZEW1/UNrtjdjw
lcuwj5emvUWfaOz30FmUEL09OllFS38EwKTNmtHo007SWSi+gNklkkjKMAnB804evEyuH+ak+wIF
B36b7SXuWkzHXxOozvLyBO00dBsGyMcprx9OktsR7myFe10CReD1btIHVLs6oRSegTHXChNWFBbw
pGrX582LlVAeJqraQJ0fjJKc8rNg85MvrBYBPvJUUL7B6Onh4uVpjjhNxN6K6NNtyDZmwnozQeSv
ar08CefgrD/qdHO9axIPWekO1AMVcPlSi6eW5Ef0X+J4zB5PNLSr5baBASc5KeJU+bO5xjCRqtBh
Z4n7cDpaZcm1ErP1JZJWpuB9zUva8vJzmxhElnjoZhDXuLdGMsrKwG1XHPDL4uUTeWEiWemRBgkC
ocASQcPsQ8xpSHOdS9KrlcD9gSprGVaAn/z6iEIWDKquCYHe9cGaGhu8mZYbWVNaGI9tcg0Rs0bu
yivpTHNsLGUMmhPH/P67KCkyd3v72PzLF5noUIEnZFuyWHyg9YGfkgdocbdQWdFD74DoMxdh71ue
V09GBSEyRUqNPzBcHGz26DMMLwQwhYOkY4t7xmvuX/0zwPChi4/X05yvnka0OD5Tozqaz3WXMK94
Iv4C3A8o7MIXIjhKDKF76p0Z+nQk8Ed9lf4I5TBvu5H0UCzrd+mPlLDqQWRj88/ygkaiqvS30mwn
4IRVGOcqkJaNIngasshOimdzelO9iVnBTqZjVBZ3NunJrWNzpPmqNeYt7m1tqyrfk99ewNb+H2uo
jJKCkjcb+GUjOhA5B/LX1JLnhdlETPWuR5NjiJ2r/XuWxKTFUKdIGHPlIwwdIvMqd2IYBNkU/HS1
EVHGRvvSsKHftuSC8RJvfIFJpjKYEkAP2ZUBTwZk0tsue0Z8IQewIWmSp4remVzBxMfBDsK5g++N
ekJXWoLYqNcDg6rPaVCd4UdBGoo4bRkmfxRQNAyTDA3Fwqs1oJfyzlnMxGAeXWvJ78h09VzPz7U+
YpNW5H1WZCv+2zI1QavsiKUa/Q6wZerfdwVKQFgS6PYvCvg2CYEaamOFUemo2GTbs2dOoD7mRB2e
S+U6rxsH+9rVdwXUh5mOAS2Ct9gVtObPIZhVl9RT146LqT1uZqcgfYJGjT/VmAEPtWqAVhv5ar7K
osvQvIkfl9xvkZUEkstDRGp+kpnwIYnmFS/eWol5GQnom0n0o/+CxP3HZ+kUwjy54jI7QqeAR5Mb
kJvv8zt7Psl/0sv+GW55RArzmh/NxW8u/mQekV5xqyuOj8/govLSeWNZE/UxIGLiEhWI45Qvmi+F
QaxAkfSZy1EWOKtACrg2Q40Z/4rTvpyKeiW3Rn1M92iK6fEbByEzJtHqViMjBwyxFTPCFPvWRwvr
V/l7K95C/quWIbC7kxY8P9ccSjJuyqs49FwDsCuxDMv1Qrqz2dqeSvZoJd5ROOhMW+8opEqRaLJV
SowpnSEMr2CcKzMQiHkBn153H+zN6sjYn4BfUymt5HpQenv1CefYWeg6oROdeZ36f/mGYLNZwS27
K9uhdHdAUfzJtwpzpgAKhCLAYCPjbJB5wODqfTq1bBa6zAftyAr2fLrPmxlG1OGKp77Fi8r3Qpr+
lnX13DvN3XMeiN4IB5YGlVj3TZB2UKnEyDRierZsiA0G6nd8I0vOPaycNiJvgirVmc8c+aKJSLcn
xopLd5p/1oNooyN+YeVibP1UU8Q7rsm3fTID2Tv7cYD/La04q3rItyOvsa1/onjMI9ZKDw3EJhn6
j2JRhwIcXLMCR0sG8eIYzch57TE0xkFS1QX3rMcw9R30s554IJLlLpsgfqAWCPyBZqVpc8cyMbvw
yWLV4DQkzeLXSvdTS6nCibojouQWJuSIX1CF5tyPHuXKr6JC/5T+ZueP3SB9n6AGUs+O6sBUh+49
uh3Pj8DCAl+knXkuw7Fp8hNHEmpaHpnufru0hCdygUid8kBYn5kgZcuvtgBwKVmcj3c+DsdQmPUP
5+tHl7WUrlz9qffZRG+DhSfCT8/slB9IzInL+JECBVCcVcQUOty6FWDTZyx93QJBZfTys706a7q8
RvoUZcOHJdaVdKGVF8YeOuQKvG1NsQONfFY5xRIzJEezb1RKWoSDGKK9GsRT3g+pBQBaY1mL+gA1
SIkLldYHVtlHmqD0lSVonFBpI4h+5J894rHOOF9G5UjxypwDk7YO5TjnTU5BwYgwQ+Ar7BL96XUU
xXtYx19J4zMjS7slx8KHT0V6VzZn5FWHUQzm9oPkVx2xKqa+i24nVmQ3V7Do7CzSEY9PytKgDNMB
Y9Kp3x23zVo3T/05HqmeZejxZYBGWpKOq305PWPVFc5OlzZwM7BhHmyd4NO/bjjzkpCkE/128Obd
8fri1clQzs4EJKAanXm7Zh7H+nQLOzx8asmfb/oiA3EHuCEYA4s1YIfZhTqHlwE+wkK5KUL0sxGa
gabnvD7absa+pjzNNnII9jVay/aTx2W5ryojYS3LxnMN3DVdhVFrq7m/kKRKPCdVx9SPHuu6W6My
lOW7oxScWnpEzlZx+gDmFzgcg2NF/SkXnC6d3sh+an7WUe8hkqACkXrjjHs2Kg26PdMuj76Ynl/z
IUvK4uXsSxa53zCNvW1ni3EpXLPaEQjI2gvYQLnRHVeZxfnubPKRJNId0aHaQg2aGlVrWaAK0s8J
yXZ1h6ytZtREHW0D08+tY8FC6Bn+Y7mVovU+s4/6STqTT0nqq84y05xxRYRGwZ9KI2fZKaRczCx3
c0ZHal9XNhESW6hpJ7aKj0+p+YfCmQBmAjeW6XjD2yorS9mc/AiDo8oqTZxryIy478HYjfCi5ui6
vAyhKroTIqpBBapSzeAN8gRd84gwAnygR62nQYl3ABxRofJ0G4VtdFmEfOu5/J8EMpikvwx2dWwF
PFQ9Jyg+E/C5qR2L+jh42WwrvPIaOP4tx0s3kCX14mQ55X8N5CBKxEZdz5ScWJvwkrHK2fI6Gf4R
Zdn3LsJfV4tJtRdko3h22ZSCwrhS/JejqH8I+pGeac8A73tlUDGXc4uxgTsDfHSnlOAKwvDXAdR8
/ttgFwPv9N9gK02IqLBlffpydwz075OLw+FoTQHoJhakpWy0q2jyq8R+sTx8MnXgqtc0NFACAWSo
zVywh8hP2swYR3AY2yxagLZBNWLt3gjaFzkR/HUcTXo2DunbtRrYi5OI0z/+uyQAwEAEYK06vqdk
tykuTwiR0rDA2kOX5KUL+CbgJHrJi/IbQoKtwqMbPq0o3J5EW0wFQDmpUqLVoXV8QzwnhPPK5bge
Rcsqg9EXJ+pIA371OA5w3ubQLpDxg18HETSZiVTzTJorkVk0ROwnMtT1445aZR0gi2hXHA6bGWsG
JgT8qMdGKv2sYpUCbl4/iweYRcvjqv05bVGIb1feutYHb4kQDpdKXAoGZ6g8mXj4Q7FtWn0lx4WD
ILh++PlDWxaZXIrpoAhgnXg/XXMtmMWciSFb5eeg/pwHA6jydOOP7RNJJKgn1tfCpouu22G/rAMl
SPEkdY3EtI6fQHl7vbNsmptbmEc82sR2q1a+FTaTAeCV/OrY+srn4SU+ggvGSG38dC3bV5YdmyVP
1rdvC2BCJPwJkKPhrkEHiP29Vhvy1cx9NTnLORYZexRH7E8PZnn+6JaTpiWme3hR96yl1QDQJUrM
rqaSVPWCoTVTDKR6FG5TLI5qZZ3PpVwSTAvbQwTnBH7+sVQabYh0FtZ7pCWgKvTJIAbeodeH/uCt
yZQFFyI/sZKfBlSi+6bZqV/uhldF/3ffnZRI9ZVCDJpWKe/g3VFnb6ZqSaPwGk2cXrC1CphGhAdY
cBHqk19oGmM+O2XxNGPkc+a2Jz7Qgim0f5omM+2pbnHvevPUuUFkAXfdh5vIAPSfXDvJgSuuDNCn
SX7+schI7TqMD4gCYZQYWTvD3SKsrZoyc5mZ6KVJZrHxq4Yqyzz2mQJu5cdUKQXsaLyO7+qdMuT7
FSKEB3oAJb+b0qo/GiPJqOSWNaxFE5cCrseIxR3TVy21ulUQRnW7PG9u4LEQ2TzHFot7m0e6zA2T
QYWp7VtZU6bwgHG6XQri89M5ef8fn9/YZPNSmtjODLqhot3NU617wKNQvJVdVA2E/zTJBtwugk9T
b0gIC8ygiWn5mJ1ecBDSt5W76OaBprl37+6h97L70H/uomQmEmeYwCbH+nnonURy+S/qam3vyy/W
8jyDEHnGRCNuajw/qTv7QH/hcJSIVewaEB7fEDAt+1/0GkCLsmE9RNflJvvkoAWzfBx/uOnXIF3Z
BsLJOtBnPG/YrJomo7Wbfxl4vs0tyamUejlOUTwLJyjX9uZQC2FKTlR1ccai8p3usp84lZGPgH6X
wzGWWNZ15GSoArh9l7tICRloTbMms3LPLjH1gsRveVZwOh/paMHs/DpF/Y3weEGW8CNikMlQHyLX
zATU12j4teJ1n8878FzR48kQt6sQu+F268E/5LkD4laChVfCFcfPd06jXWIrtM7iKyrtyOFqmGbd
JV1p13TV+cw+xSw/s5OVqzwapWiQYc8zsPADMfYa6R9K5gepP2m762gPDu3uUIfCkUfe/DiMQtRr
GNuDK23zb/m5jrhYLp5d+JpBKT+AmUO8uT5EJnN+tuLBwvOkaOjHTorcg9snNZo4qXQa1LUJLfen
ZoqwwpeUcPAJxlPjJH+wmDq012+Dip/N0PsdDP9Ik1QXOZJfNQ/VKLh3b7K6DKE3aWwVILtdxIJB
URfyV2lORSINOJMFQlSO86D4KPxpHs2gpOEEgUVsuHUMjBpN7y5durmmI0p3bk3Y4562/xGvNSiR
2FoHU5Ji3EBgmGoOmMxhjMQ/yol2ih+XPS1+q3XQkjr93c0MR4pLVh2KLWXLQ1uxXLnTI26/46mI
bLMLNFOBAMPZRs68j04nvr2aNzuRo+jlJiY8CI06+4aMz6ptrXD1UiMyyfwsIKySwCimhaImLMwA
DnFPk7PfHtnGxTp8Vl9zMp2FwCfHpjpPRC/LklTXbKYMmcg/JgjdcReZAlzsUbd7AjYS/BiOZout
oYp9h3agZbuQ93uPI6ruC5UUx4nemvdRvSooIjs+fCZEBMmbaYQTneT9s8MiZGGatsnTtiRSaw3y
VoBrCuUD23dqaqYqM08I1ySpm9Rzpb0E1svN40eSVaVRtL1uJxeAEYdrFJH2c0uzv3kxyNc0QZA5
SCwHYLvaT5lz2STJSaymO7APAZbulCue0c88AYPp1mxeOg7al+rpCSHnHiOqMeKthFNxyhhsnFjR
QX4lTw3KhsDoqk46b3k8FF2QZ9s1CPzQD7tt1ehLsQrNujb8t+MnoX0HYxLgHBi4WLHnvc5oUhZu
oG3G+ex9hMRoRO803GoaiofHolIuA309ocPEPaQG0R1u42jEeCMQ8+JDciIqoYZekMBqkg+kHHuh
C31q2IK6jGUUB4qiM9olo3bVS25THV80TlqJyC2pg2DjHvLFvujmQumz5EJlWcK9QMKMjB5u8ldT
CPySAKDtZkpe7q0+XiwraWNworNuLB8f/I+3fspeuw0+bVvxLpdyzFpH0j/JDtiyC31ueBP0fPZH
wUU8VnYdJ73pf9lVikUpZFXZG0SrP+lFcy7dBjhuKrP0DNm2DFYIVG4qkWTeEQmCg05D8Ap4ad3j
Bmc6UeJdA+F1BiBlx4v+HDGBs6CM0bReTP+56UpRYZM/pXSY1wkdZ1EmsJP9ZURQlb0Tb6AK2NOa
aCc94isq0G+VwF8p8x5NYpHF+n3MAbIroww6TIA8APDqTFC+Ah3hFTy2aZiwyG6IlHvuJMUFZ3p1
s/fGrzjDShOVChUayUqDujQxV4NQMFX2r+jK2c83dZ7Smw+eNvXcqqiv2QQsmyQYBoeRWZG6ME+r
34mfk9GIfcj697UqEFkQb7QbZ3yaStlJ1JtYobsx8XjbdDp9qTWgq+8n46MKs16newayNlxR44yB
9uLQL076D1uczmMhES2bD8xH7zhep8crjs7hrTh2zP8//z3gW8CTli9YakS1wvJ4n5WALfzlYf+7
yPwekOgYnJpYdzWU7y8Z03HDt1j1ajCn5eMR5YzY6aZI1rWgv9TemXRMw3R7dIGNXRX5UIBdxZVl
J6KqXZ8cQP7wdXQSwzpF3X8GrphuT/mr3mA5AM+Oeu6gj2efjzyjohEIDGxG6SGgm1GdJFS/M3L+
zxw74/AAJvRp9qudFsHerpSEZo663w0Me8fL7S8tI6AZioRPgguP9P0O1XuY5gz/kXABXwIPseew
RanKPyAb6cz23dvL3l+5vVBne/VY9SoW2hkCKiv0WYn3QMDdQuunPdftu6RKXEOp7QkZf4Qybt0t
o41+noXHICfTWwn1+UyaIhDtPk4jnp+O4kyXDpkhLKVDHnptBPtlgSvNy73LHQqHDu36wRVNSpR9
z2OuTgS+w9Uq0McIxV28smWAZy10aHxuwsioof++HJYdop7UKhuan5iNTetq8ji3Xxlcmozs7tvl
mam38Rsz1yJa4K+gEfT47/9izEiHNAlcn1HKwNgGDDsp2sag/bxB2j+RPFASUhSD9meKHZMQid4B
8mmAxm1Ot10YR43+gknbkAxRnImJ6YKWeu+u874mdhtzwwR3dUeSljy0hjLtf1bUevWls6ZGogfk
zetsbX5UmRBuc+V0VCQiDCfemLKLPztx6vdXrRlyRTr64WZdfhmfnctpDnqzHf3BWJE2qvgo7Br0
mjhF0VwX6J15leg7TduZHfn5p2mYdQQwRM3IyQMemtkdjllPwskW5M92xljQiL/1xi7ObL8qA9LY
FOnWOWSrHgUQTL6iED3iuj+QIQXnXJ5XvvpA2p56hUoqwSn7z5Ct6/1MKJpVQP6t6UFITGGkkkkQ
tT0TjJawyfzr6t5iAIFdMHE514/2sT+/KA7GeQlc25LVoFpGgB5ZJppCnmzrx1vg5Swq0V2aigUJ
CxMoLeHvQB1OtJHQzjQ0fWHa6s1BrvzVwbyYbnkpEn6RzBet0ilRID4DecVuyRWhr9bEXyvsjDhP
J56UFjia0vcjA7ESmV3G3MMScACgxVOkrq0JAq7QNtevLHep2XgqZ9Ew/MQ2f5Sfe0AFchmO9Yjd
uPQToJRGOXuu7q+NrOg+S3CWifP7R/5sAxHkn5swykyjK/68Q01boF6OrrSI7eFBTxLKPQFViAz2
uMyasl49Ti1LKr9dN+/Nx2DUDOIB2+mXr2YroHvrSwL3g6Sbn3iUMzHp/GqHy2o2hyetfCZObwHd
6eyQ91zQa1iez8I/edr8g47ivGIkT//LiabNOZwXxdNHfHGzMmDvZHz3v8oBMmS4gzIDZhGBt/i2
MwgsCpky4GMfw907fdLs8siGEZDqf64ffTmipcJXK6f62Fa0bg47eh1r+rLobjJzyIjzJb8ihqb8
TWoE6oTS5Pl9oI+5FduE5XN9efONgKyXmMac+bPBBOL4mh4gTOPeEFKwhBku/lnoOfdM30IcRU4d
LhDbz0TbwiXmi+wE8L6WuH1Zn+VpCEjTSFqyPoHEtVw/kcMxGuunppsX+WQojLRFio36Vh6w75IB
ZQ2hOZgXJu+JNLlfjGZ69hTu3LZFGk69th1+rcJODDDvEoWGxNQD6XEmcdRKVD+ems4vNpOmg5C+
iGwyq+uWDmMEwPdKXqma8KL8Eoe4H1MqST5Go6cYMdvrzEB3FRvVkkTX7f8Ye5JMZuwY09ABg2XF
A9LfG6j8tSxwgZ6PS2g5yzh5HVu15x58Trd8AckyyhtC54bqjkyfKe2qKvIfc7V8LylAoDwaOUjG
ElBfwWT4YQn3XAaGKilE0vN77Inb7zoh1wYjwmxjE8jK2efz8XpMrmeh/cV60J8M8HIsF1rei/uy
cPbXV9aeL3cW5r1BOQ9RMru7H1vSgqVsb3VVD8CRvCKBl+/4EJvxto4520jtRDpB1HWtpuwnu+IH
CCf+CSJGmSXWGaJkdbnsUb72GUgDD1f5bcLOBeZ+dislqmOZCo3702e17uag23WBdpOON+iRVOp/
TqBPVnykFQMHb8bZMcSMtt/4YwsTsNUTFq1BQPBYKT+Xler4ZmHDsx7n28VTqdCuzHKyUSn9iK/m
Af+yGRknOmoBZUa1F0DSt1WXFHn6tFkGGrx4UMNt73vGyNyAWeah5MBofkghMos47Fx6YBqEeVjh
ncKaZx+BWp++SHL8EalX2K0DchwWO8Y3uoeh9uxFHMGrSD0KfH0uPGLJFYZa8xc/RGsuI6Q7etOi
vmQXKeZ+e749Zw+X1YQj+Vt/jNHLOD3yeLYruZKq6MDPqTzvElnFvNZZJvSujcI6hc6TONaLwsul
1W/tawfdig2o7hUVlPkAH06Nw8CCk2qTshFtPTZfIbr8yBpXfVUPTYFL4iL63s6IoN5BZbQZ38hr
cSONO1QYK9jasRHdkzNPkz9Gm2taYcSSBvjs+ztvW6o8HWlc7/FqBzQE0tAulkSrkm2f2eNlpHNX
Boz+mPDF54Iaayj47LZOq7Q8ZiIl9W7gw8yTsqVyBq0tQYShwIf1voedtIdAuD/T08LVKl9wt/0V
0wEt6sZO0+FOFjG/TzxZshmlyt06rYpfLH/1hl+5OxiZCsJsQbthmo4J2e7RA4372LRP5SUELV60
gv4vge7jWn4IU2KVTfjpWguS4v2FEu9tsm3jJzOiO+9TJyfsI+6oW9aymnU6XUcwFRdz6FMSAQNV
cB4Pa8eLPhTn/x+9T2vhAxoOjcRw3HUYNXeLe/O57uw8QbsaBUQ1+pybRAr71euzrmFDSY5hOWji
qwMcpoyWz88NmuitrKQ2/0eklbwRzudu5s+BGM1b8GlJZ0m8uuTTtfVVNceIxUTx/LmXa5DW/buw
uRtBYpfj8qwPbihLjzE71FNGDd58CIGO9glrHi2yn0OgYvVtGu584VNBk0rXQxYDYWa/nJPLsKKh
lTeNQS7/w3A0fXuVtXbeNutBlhwo3k5pwPUW3nl7fqcZS+u3MPCDIEFKsaJj3EDDSywPg4rGceia
ppOANwgwHl5by7EmT+HH55KdEOncku4jQgOXgowWowsOkEudSQs/LhUxwxo+RnVUFuZ1oBp8W/Or
H6AjIDGDWQmR2tJc0Fa/qs/qW+9sGLHTLaPYNiQg9xrj/G26JeZn29i1mEePRY3jXX2xuZVPw2aa
GF+Fh968bk+8oVOFz7VVO5GAeKprDdeC2MIIkcSKOgrrqDEtlIBduBJsxAm2AX5/aYLev0IzTjR9
jCTEFL9uIme8S2i7NSNEoDecCmZckW5iBFpjaF+P7i7lHlIqVwq++BbhMFk5PsbUMoXeNETmM03f
lJh+TFNzP3cUUWq13RA3piudeAO4t8yyHCWnTTCvWrHTgCEn0peiMhTXAIs9z8HKOYsSymwTIuNb
A+YXo28RVDx4a0aIEWSVWXDThpS8qSQI34nM+/AYzs98hw6JW/0ZjpkUGsCO1ikwqV/aTG3nDTJI
9EzILMVzzCVf0YD6vyoe1OW9uDbkoZn4q1Z1mhqQXQ+asI5VK/fvmqOPd4LJFt4jiWn0PjRHMGia
aqBhPkx3WP1p9Xi28H6lhoKATxlj0cJUbtbspORG+N2amVjk3WTyyxroQk6i4fnpFxpF/Dvw1Vd3
snJ44D22oEGI5fEc8UthkuuVuZgJhg7Zi4yneP97Avv9Bz1taiKsCoauFFWf8yVCKiruB3nmtjg8
N7Lcj3b9MkZDXxoaKaKYRv0zJIFXhFKp9o1o5fofEw/syTDAD52RTMEp2YAZpvinW+QE4KmU6jON
TOrRsGgu5n0umO/f2NtgfHdpXlSDIL+U7+N29sluEpfBUjYqJjuDeHrJCv3PZ+DPoGXsLtQmKqGA
DbTX8DKsUX1nMJxlVYIkwK5ifWAf4TFmFslPL0042BqlKmjQrLxpwCimXUPIyOqq/z4zkvdSq5rA
tdjqKv9ylJkyqz71RFSSfc8d1D+LBIoaLOjyiNtTJnOnk8P9AlNL/BpdzwHUid8riECpD6MRwz0O
R+PIBXAoQAWLGNbj/50xlJPiKEd8hra+qim/QRf+TqYBWABMEH6YD9xfGJ73DdtSZxDai9ptBfu0
cyxzz0bQ82nDyNtHMv6KzgO7hIaLBrSz7dq2+kZ87W7B8Ipu/SUylECuoyGO1MnOlbSAulLkxoYP
wDJkjOOXb8Q/XUu79eO3lrXqUHcPOWwg0c15dcrJ2dwA8c1qWwTuybwo/zWanLmuy7DP9IlYnHG5
pKsegW/PR8h9XaMgY1tePyfsKtfq76gVlAzGcS7ENwW2UQNjAx+5XiAtJn570WEuY9gRewIZTBWC
OxkzENIKXeqgU11bk/4f5FuJFsQdm6/1J742yS2839H9qA73ZktPcZewtbaU28E0wvb/jPVEKING
IdK+xYnSncNE7Y+M0qxSouVjBuVBpRyTbich0TZhaFVxmJGLqZd+rvVbTpvK5Diaw122LJT7SNFM
7YAyaJMksyNN/eeKuahWHtdlT0O4bl8t7Tt+d/bnxrVuB6PwtxWymvkeEPqPSsA1SxGT0lvyIRiI
xZYaBuJKXwMXQPe5Jn60/VOfqDYvO1FXzM/I3E8X9FABqRRBbktiLHC5XgFVbf2j+qWKVNoS5HzU
lohngn1qkCUK5NQix+WDQBvN5Skr+P/yltFlrWhcvgM1/aXi194yccbwvZE/dTy3j/s4P0a0Kd+m
2BVAsYdWPMoEZX1PNmwfwXtYDet9MMmDr1wNEtDrpeIuSFHsEdcDODnD3lIA3Vqem00MKyqcOldY
rrGRD5yCI++I6fZ7T7wWe7VidsQyvPbbrODGhYAYiuXFvjPPHnGa54Qdvml2tvxgHIMJHUFHSxCT
eBQX9qKxjRPAzvvkLxUPrqYSSfgVKnjLVUlP9g+rDTuZybCMT16TDvapDOXhcCd5SwFxtJfnvumB
o0P5ZiUVJ+uefdoytudhQbUZDSvQY4dedWMLpf15mt1VTpSE7385jkHC1Qa/s9uUrA5Xd/4WEGby
ZZMekQQ2cFV+wmpKXAUcFaLav4f7qjn//5paWGeSf7Iv+DH1SkN1s5WejKiGAE65z1v/wLD/hEmb
7ifZ3V+tm8pFPgXgw0JL8gkNcR9Oif8X7d2uC8bMqD+1eOIfIoVXN86By84pC/g01bk1qZMk+wyM
AC0wUaoUs0RAzRNtTB7uNYwRCXRrjb7P8yTRvh5+UIBnLIJiEFwMtFfvCHNDdTwz5G9Cx/u2Ukm9
o16S590S5ZXx7S0W/9DC/2Gc0pa0cFPB20Y1vhCqBN5S2scC9vVqZBF1yDeT+cC2zCNJqpE6cNmG
HDIxkNu8zY1DIvlMgDwBxFIq0wnvK96k7iRXbxy7zY2CLZMaph3ANz1H4Pt+CpQvTEAJ2nVTiukd
fk/slc79hUBWQRez3Ru9Wscjfqj5rPH+eSEWGnnCb8RqDVQjNKC15BIrtUNP5ATcPEgdCjmlIbyo
4rVE/MboFIRUap9I3oH7m6p6Y3eR6lQTSn4c6zhmx+C4nf92rA1xl58Rat+XiDkd20Y2JID0HM7U
wfCyEM8MQ5szlez101P5VvZASaqh7mO22kevqk1ldRGowxEfpiFlSB7F0I7Iq8KQR7fvnD2LeaPA
2glVSShkuigqYOkRg6/fzJGCjYfOYfQrS+4GFE5Dv+FHplYLjvsLK/zmk70eI9PpCmQ++h5OE9K3
XYeXxfRpmT6oy3uBNg0BR59YNdnv8KiKRuLgbJNojoquuJJ4WU7sQeCI2Dm0nzCmCbOcAbgQ+oSg
5OYAbwT4+DOze04CZcwTNCY/boMxxyKBIXlnJe5wOdmxw7xQm805FZxZSNZ84dHpbwZJSWe52Mf3
WjdfozlOqarhJw/veu2rmi5kcuaG57ZOXiwa4obkdnjZO7DYV1Kacg37ThhFA4hwTwwo1T/L8SL2
EwNq4R9nEFwJMrYchJj235hloJ9H0ibTdfeW6sHx6QpcpOs256y2St97Fct7eUIyr3vYblxfmQ1k
EGjS/4vUbUGBSAhCN5oQL4EDl4mss3CWQaa3Ao83YA+qbYUlpi9R3WRN8YvFLoTifbibCBXR+Iys
QGaM9nVBMy0pIi5iZBaQeesKrJbPILyCmXK3443Gfmoshx5Zoc/+YxiV0Vbpj/CWPlWdJ7QrLeLh
p+s+zg1WBNVvT9iu6Vc0a4j+U6QubE8dHXC9rmf+jsH3p/wGZk/GNoRRyEQvxDxA8e4xfHut45KX
lIcIHItSO3WMyPPcXhkIFaWvgiIS6t7cez9DT+OUyVRAB1ZQs85E8Vz1Ngzg7ulmTCF/LyrZ5kXk
5o7r4JUrLHrZTYv6P2miJYfWdT85xwDKSJyNyUUZPeaE0oTE+/poKciMW1s81RJBp2Yf42RSEWpc
7Y8eOKUhW+A/962WdMuHzj/WbCmGnRMvZTNPoUUo5jTP+8Ok6L2UBKiWRzK/s+jsRmJRYpm8odgm
ZSKgPyAlBy4jK8g4KY2khR+rpajpQ3rtdjzjUiJ1GfnZAlUigYhK7jG3nn4TIRWS/FDKdDbLslpd
CFPkzu/pZID46hB7hf7mCvbYgQ41R1qqvXa1IlEcsFjWj0jAcgLH3YkTb3j9+geGypbbkkmxgYLZ
pfx9x7cldINQp90z6+VxSUEhIa3IlNwL1YLJ/HwYSnwXcHJPN+2EAbqKiQ0jn/xzd2c26UbgUjyb
LphCYBA87ok82egfKCaYIF186Uol/S15wG2nfP70DukMmAUxoFj1sNy6ox9mh76OjOh2RuIfoHPv
Bv/bRxNikpiY1gHxJRIomqXr1A71D1NPjWe4qM4jYuA9pYcYMj7kSM82+hOE5yIyD4cM0bF3B46j
9voEMopLD1ly7PlCBvn7R0zrPtZxLvGMHOnUL42zXcLTsDdOm9V7yAHoyxegYWqyPxWnPaDH/S+V
yrUxFaxVEkh588TeMqLpTaXSspGXJw5j4fuBC92B+X2dyW1wRP50J+DKSmNgzYtxvWR13VkWy0uR
b7V+z44juIunzylRimBLjjgI4e/jGOMN3xHzkB6mU/K90wMii4d5wXts72SAOdO/zCPqEcSJSZlk
1eeMQHv7lYsh8qzbCA1dY3lcjqspgf1f/TXAsi4VLYO/R+YPmkNkz2yP3e+Btks/GgzxBHzXmL6O
T95zewrQs2mrdW0gWw74S56/tmcRycq45Hqv4UwTHzXyv39wTCGBXAtHwSgNzCbFC4X5T1bHFl5c
dJu7HWm6xILoYD6Pd+WGOSEfqZmBiz3KTIWjLNQ4xjDu9GkvDZulyYtF4xg2Esv9p/DP6+VSMR6j
fYbbDrPaPXhpdnmBew7Xg9xQwOa8aIA1YYmXV0r0RyCD7y6afwVJHyUCXi+RxrH1FRpT9usi3k3O
wKxhNSs5ZFa0taRwfT8VAbJZ8DDPZUqmkSxRn2kF7cyXeoZXkOUmAK4PW+lcZaa0dwr7cj0YyqP+
88YmyjNix0PbLe4yIJgyAUVjd5rK6jZPG/fvIcSN+AB7HiEnPEKXqG8IMRriXSNfRlaMnmgikp9E
xEenMvqWIzSsjsChQB32CkdYwi5O5mPDPPXUOCV1hDnT+WPDWeWMGZHjB8R08SZK+x8VSU4kUoPR
yvmP7Vc1b/ce+Al51scRarwFyUIV+FcLzN7txLtvC9GyOGxHd85zdTNo2rfJFeFbB/M/Oc+9Q/Al
8JYCmHf5S25T5ERLaxGz+Q/oIDEt8JvX9ebC3MU2cnJGHGxg4QJYpStjDdkXvvLBT5jqcSMl1LkK
ytw9kzs7uEe8iIhpe1+KLhSo0j3tMXeym9aPiQghuyTRTIVIvKS06kLAIvYeXyqnndyY94z5kMKz
D8YlQiGIYDdgMjF0Mz0ukkepxwBZPj+0boo97yWpvjt0fn7Dcf+5iyP1Ogy8SFkFErbxh8EQsE8q
prL+ulszjaDo7X+v30Hgp0Oj71GYeJ4f0vC2ozNsY507YFwDi06Vu9AdWyWlJ3kyotZTWCTDLpdO
HOPKsO5oA68Z94Ac1thYYh9xJkQUEoUkB1IxTp0Jr4qCZwMzBmPm+wtT0mqXAz+coHw0+WTxzDBh
ViLs7QURzXvL2R6mTiLXQedmOKvepGfjph9rosv2XpInSCdlkGU3y99DeaOz/wQKJU/i/gSCBeVI
nHzndYpvUs871bFyu/nN590K1qy9Oah/819DciF5szF9pKgiCxu08pBVhl43DWdhSCqEokkjJLSq
rKohtG6n8+ZpVKW6Cs2pZj0bK2SPPeviXoa5b38wfb8h0gJlGLbZNN+mw2wF2n0iyO/Hlc38Iz6e
+bNoQMj+5U69DB+ofySyH9pvYPOAx0Xtj7ksSLoDouiRJD6JolMczrWMiWoI+3g6lDLep4rLw58m
Riay3EZ9V7F6gtomih/JRfB6uYXkSyG5qTjssEK5Ke+cS1rMddVXowFsrSTaaP3FKl+LU325KGZ/
ohKOZnWWjONINlPmlTC6D4jmPe+zBYkZqc/oX0x2LxhMtQFaprFaLiUqXsUCiKKycqf5HjQh5RTx
2JpMWYpjMY33O+Wn9vH0Q/0uccz3iWIhwAssbG8kdKzetZjWQPHv4UPq72JpMcjCPFwh7JarEq+U
WWMvoihFPr5G1WSnBoMboe2PYX2/Fzb82Sp3/cT54yFtMSo0qsq/TMIAvHcjMGLtQK0XveZNndSX
e/7pGzyReAvAtjikUPx1dlmCypsT9HRZEtEu04QrIDKBwVRbGpzmngvqRcJZkbV/QXWzXZu6tuKn
F3aOCRRep7kh/+0tVIfzLTVPDj01JCtIgxnGPUYT7GoPHcJHmE8MPe2+0oZLMZEEAInkhKa5P7tE
ibW2X6c/0ERXR439GpO4pCWCOcHXw0iQHvGwGaQJfh9ppH7kMZwhgjJz9/BQxGpHvZfWsm6XITlb
4mMM4hZ6wTyPgXJaOezPZETb7HHkl8LzExzXt87S8CraGIi+rDDSIHlm1GUuQPzu5Nr8T4ZqqYLq
WSbp+xwU8DpkBGeDwADUHlvMFJeyw3oujJJSgOmtnVwfGTSFPajSUye7DM83DRxU7FM3IaQ16N6f
5fUxPgCDEIK4+yh00XnUdLecN9sywdFPRpKD/XTZHPuldYdi2P5AI5hxUR0y0s0E7D0HAKwk0bV+
+/pYh/6/DtGGGImb0T/zY5EIOYu0PG2LUZPqcXuI52rLSPUiIlZ6ntrQ3QNTgwMS5Rbext+vpIz3
G+A3LSklDOfySrBpBbZIOem9+uFuFFHvAOCTWFGLTzfWK/5FPzboanQaQTAEoOwSeoU52pEeObvO
tYw5jQx/i74TaJyIleyraHR8XEhWwZUPyJ7Z4pu0jgeXGZxCSHR3bUEVbHMaVeJurddczEBm3otf
aYGdrLj2k0MNETVkM5I/9xGWjpuB7bmMuSO7NH7CqxyUKLDAjHTYnd+a1NkvjvyJg0YwZCfUpDu1
8T8jwg09eRbaceem58pC3fQeVl0aR3Qg9fS/0GORgWO2DrW/aSa5B+DzO/0brpFnWP0M011ljbKo
0JseD0P3p5jnJVkfKZKW20ejmD/89LORN/Ggv444zf6nPHm89ZNVurmDj6euJLRGoDMlsItthFpm
FuHxfhk+ZwaDaBFxWBsYUrE4tT4zEXfkHonPaB5Vu7DlVzrvbJpJgItoDcq8Wercz8RNhDzkMJ1m
ulplzU69HidecKvIILmDqIymwrT/3XevDY9cusMQqo7CKY5IkvuLctiR5g5ZRWeR20LWpWrdU4qV
UoD6vEGlmvJ3eBHS7A1EQvpzI+H62x7EJFxLfT/JFWxdStpd24TVV7b7j/UQHby22kNbgkcwOlp4
lafZazqkikhN5qqga2hihzBWAhc2xcbS2XCat+43FqkisK9wpAaYDyxoYeN+JtHOfTlrduhPFigw
VSd6rHSJDaGo9NFz1ZEx+XntiJQ/w9R+pimBmVWgywytpA8OPigHprnNitt+NXQ2k2t9g8O9Yrj/
yfsbZ9HMjx+uz6IRK53VB83Q7d7oZxgGvgGFWN29GLCy8pUUuN5C7os99/45rrr//1Jq9kiQ8fFj
Y66/jm7yu4eCJLKY2yxnUkBLyrrNpn1T5XjacwwiFu7ntQ6ASTiWc/gu4UGN5yxh9tZ9+7ntG/sC
J7kk/xQz4/pucM6q/6x5nQ5G5+QHEZVLmz2FWCnzg/MAtdPBcKRd90mmFrQhHQTTcdRPx6ZQvxrA
btXgwDv/vhozbZYfrFZ1S0TtwHTF82FcyZyEqfjyeokgHI2gzHS7IrCw9t9hvB9dRA/PgD0p2Qhj
Je8dDW4vwfAIY4NmdbsOAfGj0Nr04ETURDCywj0et4rs2kDOmClSgDNdPxTH5qLt/2+qO0qMtzZn
pvr8oCYIJeL+7gswBqnRqdp7o0OQdmRTu9J7w0UbpBU34FGlWjfIKR1UwiaGrv6sQk1wcuWXaeIm
GTEA25K/c4IHbKySPNK/7hoh5AhLEvf/iuyAob9iQU90pKSawVhL7oaL0q/5piOQNNmgJn7S7FnY
HyV2TrGIJskZ0LO9NNaZMbz/ASxnMdDzbnrFGtlYsHowW2dvVIpwoERhu5NvNZxMA3p2iBy/ElFV
kgX6k5rV0SUm/9geOB0pOXN1Zbuq7Vdi5rAnkkI6zdqmr3BowThr0iT84+YPLSRn0XJlBSsmNOHN
eJCLJTRKdX1Akn621BVvyPeVznaaAViu2CNOpOkw+ntgtWcce4nJ7V9uq9lDRktwYO9EBLdoRYVf
6wbHgUbxjb+2cdY889U/luyC3ZAfeD7DNZ3mL9VldaUhLlO31y8DRg90pPubXrFaHEG1xQ8+/UlB
tFc3sdYlLcJyk8XJMd2b9s5er2QJDLC8YC6QDC9MY3lBfsU906FggkImhNCbm/EYWyouXuDEMMJ6
Q28oWcNJbqhE3d/Wqgl6BwisZjqZZJb4rbRg9wAqxosVP6P5reKU8QgGEKE4zzvuxjZARJQPQpSw
9SnNuCMu8VXulyUQb9AwXkSOJPf9rseVcPCdT0KBQmq/gQw+8Rqa0YxgaTooK90lLzzh22VV4BkL
KSLoLbnJRGTGFv36yaQVxa0ldCIju3Vv/7iZTTG1OEvxtzbszMow8og+mNkdWdaM8qye3fZRG7y9
Xf9FetInQGsSYXFX7+SMH5hFFILqsKYH83SluR+KZy6l1c19/boPSVq1boWWyNTMDfRAxZMZlgBc
/lcoDFepT+5O62W2SVUkWWmuUTVBpZX0mOTrQij5ygE9+yFDBuEieHL97ce+zyvxe6RRaR3/6d+3
bn1ZzJ+lz0MuUwqhig0v0Co4FQ2vdJbrJ6Ih3JbwFJhGN898wV7VLPKSCBZuc7smgEdGI5nMx1ZI
s041fLOoalNMpotVgMGQVU3K7gWcPpAGhaf5Lv3K91bL9cZjncJs4E8v8ymrqe2q+Gv7Mqj63Fr2
4hfHneJy+evrdTkGG1/UKBCIZqQwwULBgS0ePWO/AeeUU7Ja5Ro55BqtJ3zCUtY7JMaKvh3nrLUS
rgnY3nRSrSlmRObTF7DZnW5rjRwJeeaRmf5t045SipiUtwV/I7QHNAObNjMX9E7IciUp6cWwGXOZ
q27CaVWVPvx7vpErc5AThgDAXD/kdv4Ayxq5o+NGGFnysEjNQhzRXZZlyhHiBZS8FJ5s9XH4VkXH
thrUbLOn8P5JlzGbQagIObHWAQWh0+pQEAoZbbY4VsUZlHBgrSPO0P+r9RZoBO6YgLp+P2mhPXde
mgIEapk33worLRaVzJ3f3q7lI4a6W+c7hMSdX972cZrozwQYlnncNjV0p3kuP4xPUlF5yHkw61Es
deIpDVzr7ct5j7q/PANmmLteQpq+x6GxhvIIPbZMO2Ww0OpJhSVbCv0HCLn+HnjR4wjs/gz03Wm5
Ox27zdeI5qcpEGxmB+8WEhIpVf0rCUjGirJIzuUb2Y6aVdgVlBu5Z1G2xoEDRY+syKMNPfs16vI6
jq/m/h/jBcVc7ug2toqFO4W4qylDU/ndtyXsz6fBIQix9vVff4yMbfCh2A4WdoeLSAP48RByUYlb
IOyuW6+Q0r+9PFrsa0fFXhmQlJxt1oP9gd+KDM4UwuIZqZ51OzlgVeGoXOYG81ApodxyN0RMqk2I
MjY54Ca97C8V+77OjWh028Uty2pKE/cEOGnHENPRRTsmH74AJsht+juV5MZeup9cs3QRjTzUTi+L
VHCTPgng9YSa9Karkf4zYDUFfq4GlLzM8gxvCY5eWtdVajDotcZS5xvOqSdnt1OxEwUPuz/NiHLw
3W4DGEWxWTSbPXioRRHfahDlZF0jy4OBJOQDl8xVzW9t1MtcIFHalsJz48z37Vt86fAfcNthPriJ
A8tNv7Csijkgo0ThHuHNKobobsEgCMXB/mhIHo00t+gTOtgn5YpEnKoH9sYvYZn33S5WAn5OQ0bX
NhLvWvDFop+PWXzJL9P8hGYk1GJ/ielbb6i9SEfgeI4iEcMvhR8JwN2oa0+BbkcMx67oYeRwfCQy
NOrY9tVHziV1JpNaQuK5cinJT+0k2N/bmX7djX9uWcH7VlE47V/1XQzP3S1ROjyrQEBVcutH/yQ1
pJ/VLdf+tKDEdikj4ScoiMVUlb2fTisKmrHxWVxwaL6U4eCtRT53xjD1VMEeNL24AqpkGGuxwrCp
Jj7+uAmBVPF6UBijl1+nPoTJEIJ8QTiwHc+RiesA3yPuZ/T8AQEnlu8Pgt+6FDtqPH9d0/JDAAkW
vmfzMGBSl1BqoeUi5ptMz2nIHtOZ7mByHyc09QJRdifnEKpGp0VPi9YE2w9mCFsWBtWkjsYJ9g+h
JI3B9ne/aoZEZ+cWiv4dUE2blKQS2ffUnOcCscGcPpdCvmZEX4sGPxN8HP3ssKHrFpCHc6X4hdce
EucS4n4EdG88hioZHJfM3xpmUAeaTNV7xy4GF/H8WnaXRcbI+u7rDtK47xPy4EArZ3z0n5VDl/cs
Qh5g4rmIXNT/NrEVDSHfDyaHDDXHU9D5vcc2yyr+nqOArfJQGOYHF04jbxdRSc2FJytTfmD9ECwL
wA0XZZCO5FCtqtEz/n5wxHAI9Ig6NEn++vi3cnmiVSOCEiRbq+wqgjyi/h8jVI5nYwRoBzhRN32i
05xWzLpgdBFZPeskob1JCfIP3OGUdZqfO9ZH/ysijpQPtvmn+Rl3G4btLlxExRR3enEASbgPkX47
VSe8Jkv761pO3Hod2fcOaTKMOJcYIaAhRSniCOEedxYqquQLpgxqThSwtYvWAzdBRJ1nEs34HLNC
gBpNmoHNHyM46VriHAu2twQST3jkLYYS7Q9xaja7/NslZsJGKosPa2zrXGxnzenZKIQaS2ZZ5Vjw
EYvCBWx4iqaOHmLqAS4PvJZEWKcsOSUP3ZXQZnI0VI2wDDrhhki9k3bg7JxxV0iuJUBccqxYFbvP
6TdqRgg7zZGnMG+GRMhK2kuwO2cDXAoF4uFZoo7UG73NZWl/DX/ssJUrtftQdu96jPkJmE8NPlGY
bl8q5uOFXEXsadCRejUDtfa0afuWm5Sfx6xQdckorH0RRKJlxrMaizO5gUf1T6ggM4lyk2FfWF4S
uz58UKS/a+3CRW+sIlbOllraDBirILfCKYj5WeaDZv6O9e95fhmBeShagOhxzFFOF/WYfzpXgnuy
2r40zaL88+LnZt1M/hW1Nk6LtUMtay3ivCtpCOkJE62jPt1oA8YAw/XwmJkrgF7yA0IdEYHmyb8R
ZHLNIdOUHc9Q5i0etSG947V1ZLCDBKyH+B2R99kfIBMtJVwMPXHvcc7UDcnDjoogOw7N/danobj8
9KnDilnZRul6x02vPbbedra/vK0aTCHKxeRl+gB6XRgTP+eUkKXUCet/942f+uDsE2eCZCIefWpA
GgaGvA7uuiPtO34Mz1v0rj7iQU/Cm5joO4VAWFdgG/00bSKP5I0uZ/q9YQ84Yg0mgyPGqviuxJzQ
1oYzFKJ2H3D/C15UlERbjNiseYQbGjNfOjlO+vL09uwZZ2tehU+mtpU14g85bq4XnxDmaFXm07Be
xVG4HoBKGt6bp5yFsZ5YGx6hTlea+89JOhl6EQwvwph8odZAvzJeQAxgJBUOKPiUMqnB0druDr6J
hDpEbgGjd/fM36VIWPfQaFpVWYp2LhYrkmanc7HLBU27duhdKGETMdYr78sSyHvYYrOyW5B3OmIe
6FPWMxAwh9o3yhuiiHWlWryALIuKsswUEWYAHFDge12SmVJtU+cIN07g5Ep3XOCmAfdGJjRj77VW
FnvstlZiNYAc4TahKOCQ/s4tXs6rpF50LDDMtEA6AubF/l2jjhTXakpQLNwu/IH2Bd445IE2PIX0
/mfKjCn5ei673uU471/c+cCi/J/LQsUtDPhZtvi2Qhj42lORA1w7KHEp/KOAyXiwrhrmpvXKqpFp
AQ+28FUUZkiePzQevQ0d1De1hFJzJ8O2vbKNK7D7Z30rxwgBy3dvcHb15+l34ZNs6pzGcZJbpC5d
vHwKIMJJlXniBd/X9FwiOw+x66eGMmhOLmsh5o80SOCKZOudb/bVAdm5kJeORPSntsRj5x3O8q+k
t9SEqQqcb1tfJOw76HOagAQM5CYwYHiRgmwTqTjwbyxgLiVfEKvbmDbWUyMD+u7kFztq2UvvUViA
MOEzzHmarLDkS2hHPeFOqUJWT2v6aHHLci5q8j1ctdmVgGzGtVQ07yRzsbuXTbJ0M7DVfZ1oQOF/
KuLT0VA2srh3zP4cqHBMnA05pS5CYSw35lSlznzpaQWKd8LfedHGSf67gWRest3mdQJyhqzbyAIh
hXcwSdGKsE6m3ptpCESNorkQEeAa779MnJAyTwCXiD+ODwFJIP/HRV1U5qNQ/8AOJvvIMZ4Fph6w
2QX5Kp2esGWDgNQGaZS437Uxz2X6/EsqZt4/POto8hqIZGCF0uOKp3N4x0/MVI00PPtmCUSGbN3m
6h9q4U10VLzfoJx5IYzfn3BDrA010i1okFuI/LuomsBeWrWd5Jz+BbgjLD2An8lBIPydOfJQAiUn
+KKV14TX6zeKUtFO7NsME/961gW9ocbVc+V43bHLdlhmFc1ExDZITGGaSvxTUu8Hoh9UwlJecFcw
rfa2JN09mn7TL4gToErP+lp3F1Azmf8YpuZPt80FuFSyKPpskM2dJOuz1j+SplAgWoeE2NJm0CBf
UwSkbqs5Suu+S85S0gvq2cMOB0jBrHu8B5YSsxZgC+7Q1wIEqPqSXIRnXG80LtRsDYn284B0EPbG
3fFISJebTtTTt0RY2Nn/mbAEdXwOu9VqGHIKhEI2R/vw1h6DBvQ13awN82SMUyTQi+IS3qnqoa5e
RN/O9dhxYHw8BSoTnMKwLq3vUUx3iPLh/1YNtEy/jdaY32F7CfGQIWzOkMWUZhJ41ASu7u8YcZYP
+o15IyiMV78D68aBS31VbXycllhOhvkynwF/KXMj5wLKMrqnWjlCEEaR4qGa4KHtoqAIithjmqvq
5zMr0Hqi14YUncbrkNYB0vzp3KjjR/r3uWgHnA4vClUKSoJ9wTsJ4oB621PKhyP4UeV872obwWKw
1wSSuBqPMk3K8yVkqP0oQOVNLnAyHboVklJJig4g70coR0vRYSNhAqBMZrxiukEZjv4pyYrFSoLU
rqPaQdllu50zpZBOqiSYVxoYjCoMoKTaTwCnhyv+CycU9TY5SXNfmpxZQ7g32imirm1kC7vBAEgl
/Bk/5vu/i/Yimup5UlM3Opbzs1bt0+uT0dHa70elFjH6r+6jRicSTs6Wp+Jl7f5+PmKi79rbp/AR
7inpMSCJViEuc5Vbu59shd6Oao7LWJekWg9brXPOWvEx7rAWQ/yuhqh/cA4jDOq2D+bCJwx/mzw1
URhxCGxN/IdJBzQfEsFo+nma77OEYdPHtY6suvuvNzpExXisb/nWfY4ZuQB8+hlNjIOJgXYvtHZN
Ao8XAiPNv6FDGAGuqLkvRc96V9ly2lyl57F1jmTBC3A4uIRhiYaD/14TbYAZlBJuF02Ldtgr5int
MRPO9wZE4SzqfeDmxBpyLl0waMcDGlajXZLC9g2qUz65fOMIg0AbmAfLd/mkU+1hApcf3t1LfqNB
uGWoKsFG3QyCWJ1i3/cZTn7xa44XZqnpl4fNwV270tvb4skP2ojZQWSNq5UJWG9gLBan/6hA/0SU
vO65Z9lqKhx/8IXSe3HqfbqLwGbrPMc9FUc6rrGo7vubh7yIep36BVKHsnDkrkWwcJpxflBj4cGV
xQb8KCV0VIY3zEpPcfyYydxWbDy57w9L5xYYdyt9WM1PNCzBn+sFQ6Xi8VB+nAt/z56/ALCATRMF
k4C+lilmIP0ENZ6ONpkfBVsr42rqa73QjD7wyXTxXm/8G0FUUSCdFcmTCtUm75OuFA8dgqij1cqp
MVlVurBg9PzRcdOOMKe2lc2pHrwiXMeUd848vZ+drHVDsMDG+mnEXnaA78NOsJtDbmXaAcStCPYk
IV3LrSC611gc9eKka7ZqGOX4LUJy//TcSP32TAO9S6ru5miAcuWDQgKYPDjoAPi1gWMBanvWgIdo
muA+3OKkTCsYjoq5H+GVhewnPyCXm9l0NAYg+kXBvX6YoHzoxDlCt5+cZQvfvXh1IQZTD8kDBZVl
CxxyQWNavC1vMYGT1zUtuODu1r86tDfV+jfFCMXS26DbriInA5JCHlPJ4YmFvs9sJyPGmjcDYIqF
oQM2EQ85q9T+JjygBmwutqbMaAemAFvz3hOYbU+A52GRWgD5wMN3MjBGuHvMDjsQpjkXpEALm9Xg
0Yruv0dQAP0fiNVo6WQupn0YakoxOAifpvYS4Zn52NWYf8ghNyTATOpQ5hgfgW0dUmvJ4RluI2TQ
9F/yMK91gNgxYmXIVrvLtsaUhsTqcC4Ov84s93HC8KK6FZQOQBcGQ2bODn3zvEyhP1n9bpeKSOEl
z0VUA/GeuwATP3sqFWI364An2ahw8GNfOJXMeupco50dcP76LaGAi1RkTsefGFd8VgeJxij76Xuf
pL7VEH+ccZRK20hqLRsj5SIqYQ72PGbStRASw4XQ+LYnEM1sXEW3LJfTnlu4i9X4mzSMYrqrmGXB
1dIjBXe2iLptqu112NPBwZZYoewUFN5Vd9dvlaAs9L6qHEkWeYayio0t7+IOpHVd2sgXhhN+B+x3
ddhD0fA2ZSu9M1upJL8WuOOmPs9mpr2anmuEo9ZhtM7ksBneG+6/8grG4zyj89kLqGHG5Lm1+AHk
ARckG7RE2BIuaSroH4mA5tOlXyeSZBJ05bUzF5XaAb+RyxUCbgBZiOJk5fB4z/DEbNXKrc1kJzM8
jPsShPKoLiQP7mHlDdBbGg4UtQmlH5AgilA3upkcRsGEi3B6KSrjzn8FnR1aQ4A5dzC/P8Fdyvgn
Cg38IBBB/sdSM2VTQ91g6v+gv3Khrp1YhhxI8vWOsYM31pjWrnyZeNeqwPf6pD7Zp267fWGX5Dn+
lVi2uO2nX6i4KpgoOKUs7LG6SfILQ8vzgRcgK6o5UMg6qsWcXVeYTrfOn5ML7ADr4j+oCUtT6MnH
NLkHBjZ5pt+sniMjtG6J5Ka+hD2bIpOPalVARsOm0BiF+70UysXjGRendzupdfo9+4sT1s0CKKKx
iyLpPN8KeVPWplTLIZyKgHBt5oKVGlk8QBTlo1hp3TkplhWP32cE1mKaSHnD5wQFaZ/3ovTqSu49
uP3kUyySFMWe0qXKrch0trxklcrApQmn9QUL6qxp0qhMhFjQr1CKVV8gKbNBkC1PvpQH6/ncMyyA
kUv1+z2/jAEAXN82WoX7i6MmgxtYafbveUA84fRgfuItkVdGyh8vp7Fqq3Tt3B+oUdaqLYjGIKd7
v4djP7LeX/7ptUaF7+Z7718oWGxc6wzX81rOuQDrhPTwFf1Ym8zaS5jsaY1JbRRUNulzzS9gSfjq
yHQJB5nNBQDX2FTYTgqU7N1elGf9JEZd8xQA0tCKIsSuB/+amSWkCbYSo9g6r0t9AfUwpVGmS3LZ
xoiM/3vO4cZSr8oIUT88lu3jTOvqiyRUvw3/dgL32mSw0iysnY+vfZEifXnavBV5gc76g+Id3t6c
vYdRtPndz104tW+LiwRC8c4RfSycr97+pyTGCcwo5XGYu1tamAHEoJMlaP3RS20jB+/gpmmv6rDR
wS9kP87rMa6Z3iMBQb7QhyLIFX4Db1Y9/nr3T2GlB0AL664p0OOoqRFUGZR99NGO0G0uV5ll0S7C
lPdfei0dom8GRV+jpqcV1m8ZoD6cyNb31EgsjolOfz60RhX6rKu3ullKJqElxxBvXy0o/TMpbNi6
uQM5CbJdlabwmN3NTfKlUJsJ4xW2ZEL/lLxmis+m4WjG8ujL//YZuekwm2mVdPVHr0XS/lKh8Yw1
0UQ5gqqeOiXstuXviyiIZy2wnZr3EGcIKFxcAlQ9IFMaIVKQpoYOW3u31ZKhdN5FjzqZXpJcRiZ7
gChvu9kQb7HwZps5C/njyrmAQEW94uxTjkt0Gyv0FPq3ym1NA9bEJcYxlLnMk7sCaYPbmtOojeyc
gULe9EavdxFDINsnN1Xk1OtbrQaWtlPE3eHPa1jpMFO9YONyVdQ3ECKraiEdIPNLmUv6oTndT0Kp
59zH7lIpVMadC1hTR0UXXWE/0Xr9pjK3ex5Bk9+tRekCdFCR0OXuvi/zz6h8ErA3/aG3ICPAgqWH
B/GHYnYTC04hJajRIcwdi5AeEfqXTzWoilbBLfVmPO2vEisOQhm7mbMVH1qH0uKRkaR1T1a92TaS
zsAQ1DDNdLAylZfb1pDcTLIG4M4TcCHQDBBrCnbfy2QbK5A0C7Kx0nX2jG+x/69KGiItZJBbRQmt
EvVonn3xaTmppa499cQMQyi0anDFZ6JllMEgLVbK8oGuz7Y745CeeIqHR1ecS2JB+dESWXZn5EN1
XOPs50SMMc9yUzN6Q1V1xOOB447b9eUCaDKGscoEpCjiMqGSdJ98uyGp281qbyhGEFanYakievto
D9hVAs13oS7FsXKuOW+d6v9smbXBuyoO4tf5J7b4KFB3+Ehs3Fs+ySPMpG98SK9yRUjLcyGpvMkZ
axrN+8260YH/zcjumaOx7aqzoMdfHXwV5Vil8yvH2d0d7RKDd8FJBehCAOf3xxpywv3jZfIiM+Rl
tkhsQlHITtT6Wawx5BNUQ3CjbFusHVo05Q4edlz9ZB+QLqLiryQR3ZAXT5SBJw4ZUElSMD26oOzr
gXaz12dcT5YvXkiNhNGXELbErT56Pqhg/Ufeau2xHLidMFoxOFMW77YdgfktW9NeMEkaYG1MAjN0
A9H/vwt04RiJjjNa78tJBCT3kwuKr6fduQikJ+h7HtFvlhVrM7IJQfCxCXbLI98ryDuh2/xwXFZt
akgEv5xR4G38DzUNW43LoLiI4tfAIiitS90sHdw/SKuYNQ1YBs7FH9+eCkUaxxoDUKkGjun1GiPt
AEqgSHLPqL2tor+Odkw7q2da+sksWKudVHtWJfKGqzLFivCF14Q05pPwyMOq+kwbfCbqXKl6ImP+
Iw02abQlS/Slm0gGcWjwTmYY58BEKu1ffBrCUZff5S5CN4Tz+LCE8THVWXA1BYaJSbcZfXJBRQwJ
Xz7QgtytU+FneZ3EP5CJg3qYI29HfGuMhT+YHqiUwyqyQW9sKn0kbaXTOdpElgRK923m8ebziYVy
L7e67Fk4TVGu+NCLuOC+cp0xuDMRkHJSB/ut0CctB3pAyzPWwpYNTpw1VgCiaiLrRMtXV8CbtVwG
6qOh182ZlLGza2qlzh/61YhnlJyDNIBOeF3AWyD/Zxv9OZ0xJGLDW/nggMMeLCPtNH2J2/bX2hME
4cpfAMSslAo8KhcOFtUVxAuSxOIKU43A8/JnjAT2MknLSOWRo0a3Nfv0cGZoX/Ip4tBe0YJqgJw7
PBqm21yyEZiQLQzzmscuFboD+itZJd5pKxQr7Edn4ynWSYJlfU36TK149mBGVX7d8WdB43uuef5m
xoXXKSRGUUSvtsYqQDnjyQX/wLEtoF765ONyVWpgggyGvevoN8ENrRmHICyoy/mtXwNzDX6+IheY
vUGAxk3v1hIk4p9Yfv212EoYLydyOIRNvb8/LJEmXLs5K2yX+zWlMG/xlOI7cqUjTu46JeUYempY
VG3lTJZ/poStgPCtGDZKccghPNCGD0XmoKdkdzoo4RgWO6SGOAPdlFlQ86QI77baV+6YFU3+vBFm
2sRnUeWhUKYL+YE+EqO6P3dzJ6DQf3gXJbiEG1bkIAFRWRzWOBbNmSH5UBwxdR40ZQqcSEl4GOaX
QZRX87ziGqm1v4WA1vMnxIjJKHFP2tmgxIXQjOivPpc6F8Eel8laHAhnTcdRHOIfFfSIw7YRTM97
ZD1ZOxUBp0SeZWQjKaCVYpA5Hsh1Nks80bQDnaqAjlAsDFegX8eDXTRnYypFJKTYcHICeXzavyG0
CmlphAB3eOFCgIo+DBltTJHevCWABTadKLQgBkCC7ZKjyrszZNJbNjCwF7aQy1HJkMIMGzfeXg39
I2zzyfA8pS7tT5iWlUAoH6Aja+A6G4iR17DBXgsjX5v04qwCupvAs/lBj58N3PUJPdaOfcDWKHXZ
qHGnpFrAt3LooKidCXsaxYSealsPusxw2tDvM0cP62yZPvdn+ioQoCXhQpf0pgDEwelOfd11uQWy
Iznup5rsJ+AEWL+EucfQCYC4559T62wbWowRnTjH8PP8ihE+eOOUEp+S4fA8reeS0fGuoVd609XX
fUpVu+iCSeOJFHH6iZY9cn9QzhLdSmZhFpZsD3XpePGSNwH0MQ0h4tzzwURsJMBZst2lk+I1Ao1v
1Gb6WYwTfre+qzi/4zDnSG3mlkt1mvOvfE8Hh7wUwpHAGycbCbDCKHloKABNy1CWUIJdgFUrBCIa
o6suHLF9TwHJFMXROxKjICElRceVQ+lhKC1A+tyUmXUPubksW7H67NqL3l6tF9S3Ss7e84DWJV+R
HY9YnOOxIqXZXbfLY80p/8F4tLtOlgLtxEiH8oOyQ+8OpVM2G/brWu5Z9Nk91q3BuMzHRxq3e/cB
WrBZyrKyJ1B/11MtPj3FrTWzc9Esa8qmQMW4vGE6PEhDtTUgjGxDGDvg3xrYlciwirY5e2+wUin1
aehfsQrAqqGdUQ7cPj/4fwTpjIvKMW5etrMtSJZ9xImCselbGftlT36tpBykTaeKjeC8qXRRJlrX
WMjbfw9ei7eSyKYG85FZb8toKGKISLxljERpR9N2SrhonZehdz9GYauI21XAxIqE5Vd2VKpJUznd
I/IBCNYdA8sFJvmU/tz12tPcCASBpXApRaSCS57hWeSfoNMoXZ0On2zUy/S5OyPqRzhWr+7nc6kS
sFK6qkFYMOb4Bw4lK0wg/suJQ8tVKMKl5Ly4eH5bZWdSq1ccez4blsusJcvVo8uK580pUEDgKNRV
RPqORMEFS8JeT9NLtXUHlNEdaXA+ZReqw0OjE6Crxwhi+tGE5+Ao7oQBLOcK3LXmPxJoM3CkO3lV
DeKEXDkETfbAnbi6U+ckuJnPeCDqILITHxtBdFoJoPEMILOAi0N16ikttpWggRYfnVzk2PIcXSHU
/fb+tg+NzWTHR+iYWuI/iadHIeOA0H5d/haD57r33YDbHw2lFyGSW0m2ebAtM03YJhn4F2L52bJO
St5gKGDCI2F9rD/5PVdsmj7YUwKAkXIWsGsleQ1pxwMVlhvjwcTmghxmi/nmqPyte5iyUSiXPbMO
C6uCGzVBa0jgk7vhVQhsSkyMgJSvPB5DXXVKrvHhTEkPolshHBpC7UaXrsaZtdK7uMMBv6hdGyuU
r6Q2o3fkCEXc7NaY+/zsLFdRUPFgbaVxfHv/D24ewpRihWsfcMoazbbR1o5qoHadjO2w5K2PG+al
R3h8/OyHrniBhruMeE6TrMVlj/Zx1y0qq/xB+wzjW5P/RUax8+NgdObXePYiYTc/w8LuJH3qguAV
5EFOdGRVPVVrJi4rUdSfsqkz4GbDtuWgPaF+tjuf7Ibdo3qibf9iFyKf7W46D5jFd2qPUmOgdNUr
BC+UlBD/ppNxkJ6se7V9l7ReYhLtXWj6WB80EFQ5WZXaF9uPfgBQrRV50HTFnI7UtArOF/pH6Fe9
ZFa891h66fvqxr5acddR0w53DJO3TIXoYTeknUe3OXyEGjYe6vPQLdU8q/zXAp3iXv7O2nz1nUaJ
smh3OeGAUVnTU4UHPx5YMrvpA+QcrMx2Z53WaC1aCcvyGpTLXGnecOYzp9lOmewj9FwhYVNFZepI
aM9jkV3D31YSvtZYrP/ZpfHgPk7ors857t678rBndU89Eesifk/4axOOx3c82LkKWTX9GPXHw06b
AXcBcCOPE2kJvl1bcDX25XCSz5n87SEzh6tYrmUEI1c7GWYKW4pl3Ezc1jqMHVO8xj9jBNE0wME7
Qu7YWG4BAoFBmGvrlHv4HCkCasxFRLcy2kr0OUkrgUD92q/co1xxDsuK+bXVsSDEbIzYglWykwaj
JpnyNZvdx5YbhtcAO/T7hGJZ/vgamq9L/4eSW0m/xDUNae2razCy5xyiNtXiPaEhaTBOy4vxiH/B
amBnPCCmt/eOePHwOTsKuooE4SSEYds2BgDzhY9/7Marvq5JeARJErQ04yxWxNtKrDGywWPuwn9b
pVq2G7FcQ/Rrv6ryY2rTSTQB4FDYTLak+JWXAGLwZT4z+zCUR91IKRcOUfh7bU841fmx4OYca22X
85bduEeon+ShR+7s/34tVpGBoKeRyV4jYkhy0eaBtGGoqn+60ULoxUhARZ8sFuMWbilGt5GQqAIE
xC/kwahFXI3dzmp52+BldnxTtdQrnAiS4Eg+P0Dq6RYYSQB3LjRYOTSupuceIOPuL5Idk/UGQWyN
26PScpMZGFgknKGnWL0kc8nOmw/682wxMewRFT+2IX6Kj+B2EXZXnjw+aFf0Z3VPQAnMQrhu6U4K
E7s6aK0ONmgkXYaFVpfHhkvTnZBMWoPpId8+wTu05Vz3mxTrhtkjAJ3XtmYz5xLySRi+z5IYrvl0
43DvFTynjEn9S9Fd54FQ65jBEkgVqo4hZAueIOchX32zX7XYovpcky2Iy+nLrqjKuBBWMrrUHrPD
LZiBI1nncPY7DIgVTvD2on4JHhe0w0MKBSe1rbsSHDSx7hMNYuCA6bDjVNhkT70nVS6h1yd1SQPQ
VWwEWBjlwgI9fcpb6mUhp5+dmuCMt7qGAOiIbBzpC0IZcbKsl2t11sP7rXdGnFbPUpmkh74IkQIA
CU2fJ4AS4YYPl3CfdUQwP5nLUrtu5Yy2xPTFwUKEjrBO5Jf9YQDYFe3TU1HXUtUeOID78UZZG/0j
W39PpEPzfYqo29CB7UXRVGQgzTAhiSRXbJTSswQtKHwXWvGJhmRWgRr+DfdmoWm+Y3+1E0X/s58M
NLM9Z12Y5pN0F18yVReE4wU6pNjO9c4jBpe2AtFFh23NLC88KOl+IZKJ7Ye/4bcqJZKOd1hFE+mZ
ZqtkTZ8CWSu+6Z0MN35lijhm6eWAdRFr73lZ5xKtGPIvll1CI3WuYdDa0e7cvLb0zXhKJ2mKmAll
hiyPoqooxHIlRMOB+WbaZZDYwXnHc/9kcAw8e1Pk/lD07qD9zrR2IuJuutx7+xTZ5lnFHeIWljkO
ueu3kwkap1nq9cjMkT8ez9xcupYKQdJ3CZ5JEqqDpy4XH0cX0P0lTgRtRqzDLZGv7pjrZSdqwJo/
2DmqTjIcK5DPGOW9VgZ7vYt8aGVqzeR4U+FxkMwPjwL4TaFEhFYR+/tvYpdCST2B/Lb7nlbRWHG9
vQIlkArd2DY7V3xiSUzLaoDC5t3o57lEPV/Qhr9XW2wR7F3cnsVamj6jq8HNkvLzeIXI8K8uqIvN
0ScgVnKG5e7VTmgGbbrNLJ1MrIKAD8NIwuetLyydnz1hflAS74s5/BIFRjGpbA+CAhlIuU0nYGPl
WTwrWISjSqS7ZdxTOiptoIxD6oZr268uWSKCkHheOJtog7PN5r+12mqc0xDGUyRQVyjsLrKWcWO3
OCt1M9G6L8fwhP7HjumB4oP8bSFUOWAT267JDkxMoXi0WtbgOm1hetOaRGegQxcsnqLWIbEDK8WO
ULJbbfB2+m2MdA/uuCIYUmssWt8rYbHXfmF7Y2ZvkM/HQ4BM+lX/8apkAidTPlnGP+5PA5F3x7et
5RX2hn1Vr4YsR9cVSSMzOsB7NM3JnUq/5YKFLO7MoxkvFef3YAYGIfikFeItHpYQJHc/3BHFkLVo
hRXSmbCpn5lJ/QItN4WCe4p2vnyGj+f6fXGiGxmDAEb37EXskyyB9L8zNcwy2ZFvWXIFtO3xsoPu
gOZLGNPEb3tsvvy826JkWq0vtw9cD9XCUh7d0XybXVXxYSp6elx2z1MgQES0FKfwFjoaesaK8JDP
OZPNe5RVTiN8DJsIkOhuva4hi8Tpq42vPNsD72flD9WB4s0ETbDaJsfLu8OeLJtuy4keEIYwMkLK
yfDFwlqOpcUUXFB6tOp/b45RUvvno4aNa4EfdVTU9SaBwdN2fq0EcD8pyBze9aVeCHifTkr0czPj
TVtzbNgdDKuaqNlX+IemN9DrLC+5k9s0c3WxqFEHAHl4TJNkfAArj6hWWynllhbVVOK0KDmyvgH5
aa0uouxa77Dnh0Jc1tyfI/oqGqhiET97bRDP1JtqE4U1TGnsfTcnBJgd1EGnyGZfrtS8CyqFVMuJ
mThPAkLnbim2WOyKYKFA4wM14nRxpUfu/QuOlXOAsFRJEw79jLlL5ni6B3bvlUu/ieyg1CSUZCbU
svLxfK7bblTiQQ2NhWZmkQKgzuu7SEtMYLhgXQf3aO05MPG2hNqVLproR+NrJslO0MVNyB9zzy6L
qetmCDXmHD6mHsPtyHfhObUdQLBMkOg99uivwoRJ9twYjKRsvn3IOdpZt9b1SOGuUEYuDdUXeR44
UFT8sbA6cwhpkvnRnI2lOFsTZvSAkWsI9p5Jh4TKRzZ1wKO6zOtbTc9TxXGGdZuuPQ1O3t120cSS
xqS4Q5cNjYCqUwbX+J1CIzZrL+BRACC90wrtdKonM3VGtdA5Qv5BSJya1f3nNVRlBH+pUSQFhe0u
naRIE2ix/coU0h8OAeK8tRaZp/R970lBhPa85LWEIwLVtCiDWVsUTUqoN45s89UdcNwYnGCQHt9s
+acMFaNfSHreIcA/K/ZzmlU7LKSopNB8taAOHb+hAgjFum1xmqL6RI9gh+AojcTVRuEDcTPL46dZ
miMoavJmps7+XBys8wp3pqfHcwLA7CJdj+nnMvllFe63CyZIDRaW5+wywbbEzH5AZgkcTngSnz0a
VKQm7vg++lLDWdLCr43i5ac+S3yj6gq6kINebjK/Ace78TdUlmKach1J/ZaH8LGkEtrmwzyQ+bPm
LPlJTFs5m7fMKzONdyQe9n8Cjk715pLsY0g9qscNdUmJqpvVP9ghW9kUJkh902Yiu1DKPOzHob1C
kmGsgq8Sp4w6Q/PiHrJSZdJYHkqJ6hzGQcYhl+KbO+ugnd7SHraJmBV0GsDVECNwOce6tFHrGxgP
X1s+6Y2dxWgUBnkPG7b/bGvy+81Mj1g8wauwghJbmf2jXgn+EQgCch1pYJjRC0NpH89HLJqCWFHL
nWU7O0yNLRFmCm56owzuvgRD+X4zJJG8EnCwvKoSPKNK+LHgGb440yL6Oj1+iDOWnuA5iI0lmRLQ
IBDrex36Xtf3Gdb0v+mzOuzNpR9S/b3GeY9eHzsYF1jvOhIFE6t7/oPI3XrkUPyGZj8ujGmJzHzz
cdneNoO6FJlScSzbgq4lRpy3egrDEbp/6EJooK62N2eGNgQI6WJvW8yVQL/EWq85qXnzy9GDETk8
wBZo0O47gjL6oaEYBmMyNdieCvaIfHRqqI6aMwx/RH7L7XVpGL+IQQzocViOyr/yH9rvjbBpVIr7
k6dYN3wTv7wxVgYN9Doj1C3enz8ywmY81hM1vTSQhx05w3aVPwkgtYT4aoPYvZkjYellu61N9OGN
tuMSNZ8EEnkgYLqkVMJ1lWYR3Ej41Tp0v33B9DmlwYfrXTWif56M7P9C+4z3bW05tEPRrrndLO+q
ARrWlWxcXVzIGq20GXIrWAsZSRPnpHXB7F8Z9ks6lNCCbH66XwmYdl9QWeOBsyFXDnEcB5FikpDc
Xc2DvjZS6FB3AD6EIsxsEPkrNgwFHm0k9lUgDRnbRzDcwFxxfa4yNkBeM+5vAm5Om4OIcpfzJabk
pPNuhzosRsuhAMmpi7Tnad7x24YpSQrEUfJ0ABrMhP94G+a60stJH6o5gFjEsE9V24NICQtq05/j
/OAZDJT1KF3mBBXFR+gheYiAYj2kEn3syesQo8D5x9jpHjprHGCs+1wHlfqqYM0leozh0HTakv7K
mOxQKu9TEs9Ntm1zFpClIPsz7KcZSjlo5s1lYeX73b6aFu7d5cKoXJntn9nwyOOdHorOxDe0OL+r
TiAUFPCX5s2Lnrispk858Egj+WQCRXwx9kDmn4t6XLRKw6dNQECjT51ybzPrJZ10zppw6l+wCOdy
XXKgb5Fi5WNa/gCYzaOl6nCzr1wvuu1DV/4UGqDi4VEFcyrguJ+j+gk4jyTimsa5AvOH8yFzmVVl
DYxUx/hRkXxALttsqc1da7QZ5hmJRKt+1qeTyWEU0Z254Gp4K6l2Uy4mTja9MQCzT5HrBj//WZCN
/4WTYJPO9Ohw3zRCYZ4WJRXRjJXSs6JwCZyqKqJk4eeBZSqAhK6eL2sJxTHuxF7zI/Iz0LlSUb9Q
4/6bXr2ObLpZeAu5OQbQM6LvBNcukiKd3zbZn/V0kdCPcQ2vbsxxaDOCMmhn1bTN32sqo93Nm0QS
BtZlhlEwnqFYYZtmVP6dec48cgR73I0/82glWbUbTS35e03nqeF9kGYjH3dIsHJwV3bzhC5XWLTQ
YcMcwmLZ8MBHLlCDgSO2mi2t6sWNZ/mVzy0dpsxh1IDQNFwhUz3O0j6BGpYmZFq6CzBqnWSOe664
Ai2xxG3NLjcagtA910Jb2EPzakCJm6ZdBq3t0YvK6P6YTgl6OWZuveDAiGeOixW8vQnixa11Su4n
/RR3NfXLu1no08bUGQdx8hk+z3dNTBTimCbGSasU4K2ymU/ywxyXc23NLjDAQ9nRLcAm4DujOc7d
qdaxUulyiMoUwj45Z3G1Em22K2ZvlGHv8jB7M1iUX9GeojKzNClt+ang4lDRkAP5sC3AK4zh0DPN
VPrn/QcdtBPgzjO0NEb3181ku2jnLiEnxxXy9VfSfcCPFYi6w5iWR8ycozODle0dPC2dOkeuQEG3
3w+c0JCrb5iErS0gWNpyejV44c3+PBXPzlO+lbDbyBGpWqSpRMm1wzm+rQMU/l0Dzz1tFPCICqAO
C+TR3MgRom/9x48FInUPG6NO4dYgQ+QtzyPWCXl+fmZKw+HtibkIYvyj+aF5oXjhORBjflCNQ57T
YQWtVWfV56DYU5h826ZAPRKO7NJ5h7HHzIIra8Dm1cpC+kHZ2AydtVK9C62Pb6OEd8tNylMazsRj
Q/1ArkmZDC3VcbC1jw8AN0eTe7bIQfFLjyWOFcFbyX5r4IwLdjaoJA7315TV0JmYqjXp4hrghbct
/LsQWlbu0Hxl4OzIjGmS8EHrWQgnvBAZCPwZzssSbOS0heZoaMrvUQ3aIsbnOlvMDap1iW+j3lo1
9ANUbCFak0eRfI7d037mnC2msxQ+mwo8V4a1GcZsd0FvPmY97rwuHWq7i7LGz1SvVBqABydDkrr7
mcOQuN5iyJlNA6O1koLnmExezWezjfkddlGoNUE+8/XYZ92p+kxwv0pishZkkmOBwA619nyyPFD9
rSFOt2dAN5RWHeJp2Pu1o7EVAt9nLgd0EP3L1JMzAvnPxK5/hLPj1bWLD0DDXy4QafMehk9rv+qk
8xiPQUj8oJ52OCAoxEatJ07Wp5vtRq6pUA01DJyy7qQ9ix+fVlA6PYCGbtk2BL97uYh0aToS1FtL
k8KF4/KQv0HYB8M7FQGY3xXyKNupfuKhprR9ovmepktdw+RSg07AYRFJP5TQz8ZBzMkhnb3act8z
AsKaQJJ8AM0AIvhf5ChgwfbxPLxy5fobn7rhIAJMqPGW0xS826BHYhj8zdeZJKMYW/UBz3VlBnO3
V5oW9gGvF0izDKlSiPfWD+kfWipe5ZJW4zSsAPuZfLG2pDDJmOH67CR1lwLPsCDcc40u/TRwgAWx
yRGX3PTabaVKN9K3ccmArDylAJViL4KPAb/hyJx9s3X0CAsdEjeLNO2+Vfexm5zuEpvXYrmWvtbU
/rAiVQhpO9soClQFDXCGxJ9tPzP+jGu522d/9/ohzB/nWfwrZsZGJDtOiSRbZwo7I/lgtcpUwlWV
Grtfsk9UJL0NEDBCgEtxnc8NxhHy8Gk4x160Op+gW0Sp+WPLmX8DBZXqrLNmI8F4NE9SX28bJ1zD
tPo3lsrWp64quyidWYE6WLl+LTKq0TeF76Qd3U2IIb+TI759Cwpv8aT6Hx/pyAL+NqS1zrdr4Q/5
vIaYXY1XaeHvtDuFaQ9gunNZYemV9tJsnQXdyD9jd6VF1K33N7WxGNX3+Amojc+L8Dkc1weUmzpu
4sq2DV/Cd1ovuNvJp3mAC7yuKieE18aBiW1ng6cRp30zCpx6LJz4C9xgkudbXMpOYlX793RUTU01
aSA/e0Ad7DnHW+F8KO0bgOAHWgF6KQD4VoefbbgVU4EiGNwL/8a5sZ+aqks4NgzKCWDKLY4qQzA8
pm52UZtdGb93zeBXVEcr+F9TWa5nykwGHHFCgYALfQWFuwnIhoj4uQLZMGn/VTxbYNXFbwk1o9Yn
1e8mbPvVbc9Qmw6rqTjG80DTrPumzTTKtHBXJQH8vIAMnLVRlGgSotdXgYMq1D0cmGRKJSXJqsi5
vPye7pgNfZbenApCG2oUoyb/9N2KzJLwkn+DXjNrD9swH5DfDBRUpLIN7/ssHF6MmQkFpRyVmcn0
7zCIzBSr5vsZuLVJQVFu7zG+W5HfnC6sIdiUj3crrFtqDPsrIPae9b1SHuOdroAcxQuh6DKtcDcB
jzYJiTLMMau+t3tygfamp/EiphpAhTQ4dKPsSOt41DyAWt+5IHBqq5YFhqPULZ/4ISv+N5RLN80Y
kvbQzGLGUhctFDrc8nSXV8QJPpMO7x/6cs385E9pw1Yo0L47fJn5QiaJZfDIrSVaa2VQUiEPYGz6
xrvLZ04nWgR9Gg2vBSvEYhoIW1FsKnrgGaf9b93uuGG8/EFyl4eokXUs5i/XhvYlQwFt2bJ1p5m9
+EnOpjcpME6oGQShSusyXDIJMfNU+VqfOvAwwKT1eKrIVE8OwSiWbrzpZx2pArgxxMOyrY14sE1F
XqkqsYKeD8CoGBpdUBt87C5EEroZa91HmMmXWaVz+ZMyiGnbo6LBh5L1A0/lWea3/LMMhX4MVopY
GlY88w/40Tb7MrSzG40V9TOy4V8Rh05rLAi2CmEpdhQH/XABzzP357HpkmqLZud0KmHVouW351dA
fIXcl6gglFzXAcMM00phvNEV/+e7y6tPwJY6kHKJ5FIqjJETijxdvFxYAIPhmV2AlsF9ZCnNQcUm
7QhqRpCJJoh/kf0N6xI+kZ9VZKn8iESb1Jyjxb8t+7bfmeMKrHPppy+bnKuwqsbAPtRQfN3lj3mW
ernSYtX8DQgsvWS3MgBJuaqDGskCzH1LRI3jvEk/LuJ+9kqI2zXgLN1aeZjUxo6Af/fCkJYFjhrR
xmbo/wmQCYj9y61HkyAQqs53n9PBSmc25UlLATitgZ/mDyLMSLKtZS/nz/8a20npxZnVevwKQuB+
6IeI6LQNRtDt/r2+aWCkao1kMoz1e7azwo4VZJ6YzUysYkGy5aL8sJdrLJiLyXb8BXEU7dZ1snqj
4LmR6+hOHKVVVK+mk7GqglunBMak7yWWdzNdtuqm6xikl2D2ujltFtP9Y70+/K/Eik1bMA7vb1zc
3nj5ovvlhvYmWMgGPMoiEkd5FIcGsEJ8jFXuLpChhsGyCPf0Cs3z9+bi220r36AT2TxvFPZdhL6a
z2VvdXQU3asCMUec6qDVWmPDyo9oJ/mJGe8oEu6UMX6I9YYFn3oXA1KlgxtSOEe4UgvZjVQQUGk2
R6t7/GbZhZA9FmzH6mz2mHAlrcpyiB4NprI3U3Ur3HsEuoXOFx/qAqFtHxHhsc/cnkRju1RhD6vL
fIl3RRxYaY1qEgeQLYbjpeyvrMTRGJSxbOJDaMHCA6zUlhgkshKW12EBj1AXfg84PjTg6cGuji/1
OFWmSc3pytNeTyc/4v2bIiXcWfn22Y0KMG+8sR/RGMTmQXVAKyZODR5AzkqA5BDKnY+rxn0wGC+C
KwwX+X1qrl31B4+Rish563hc3VvRRkqM1AORcIDOok62y2VHP3WWrSLL+Qf3GwmBd1nnvTwyYEst
0m7o8cqAyswarqfoX7FTc2PJ4ATvBjvZ8jwc1G4En21EHuSB9z5Lpkae1jniZt3Rl3qAaMKVN+sA
7kqaDO0RDAjERCdqIDPU4Nrb1vG+kadKNrYyXpqIB66v5ZFdH4q2G7qVJ52XLndqz/78/rkAJvkA
QIjY4Xbi6xvkbZhRtj7kGqPIfeIZGC+pBT3Ciyg60HgNXR9k8PBglArkY7rd03/xpbf6/DKn8tVF
fpkzg1wOu0GHxM4j0SPGSzKxvvHu2rY2vsIdrP+F43Wadlt0UUqLjQcTsu8iO0zMGW3Rce1HZkW7
CCrMU8fljBFNSWneBn/YLFSLnr4gjBemX1MrPN5NzGNrA+pBLjQk8+Vdqy5Bg0wQSE/qg+r8uBGQ
MYoIwcNuPMuD7ItXCeakfQFwjV9pmuktqXzJ83bF9oYoNVF4sSmadA+rLXeANtN63o7D+Eq+KXmj
kUJlBKDorTEYovAQL2HHd76ybCK5fd0pbRGp7Ge+roQY8KcpKbBDHhrU+T3iwC0KQMtQcsP9CQfG
yaHkASzvMT3mYQRu+adFrUXMtud0TJjUCT5D+e+l/4Rvw18p5XHsKpnjvD6TbTnfR6eZQknKE18Q
BYCHT4ZV9xUPqzv9UysGJXf5PFol3BgDI4ltqzFR0l5jcrKwxEM75ywpqdr0ZIzCg+WUm3vjiJ88
si6FUFRIpaKhAiZ9Ade5GpFGr9t0PZ/u51awNnH82o3ehSUGwqpjepxwwKiQggxu5dgvawqZ5G0e
gV0NXj6JFc7LMHVjiOAKuWgONINL6Re9XUDocXlFaxQuf+BNU6wpnSOcHv7s3WxDzY0QPLzilyJE
IP/BizsEYGp8Dd44Oj3HwtlkPCLc+u2PPo2ugD8pWN4Ihbzcw0RkscA9JlYzFqje6Nz6NuJAnft3
Dz+kSFBC7LEvsa5j5u7asvRC3ngZwFU8be2N5tM3LadgzHIbvAsGOQQs1cweJWgy0w6aXBj/ElG+
wWB+3/FtqOUrrT88hpKr737V7hvJBodwsvtBPQmBpvOmYDfrE/eAOqzWHbPYhLMHZIsiYHfJKohJ
WoZxMrd2w0VVqKLnGMyTw4i1SguP1rImI5GRVTL1VLEHpyUJIBEpbPpcluSyYe5CEGyeQfTkFxX1
CigsNSmVesmHbUYTSCIU6/BbSt6dsg/nHozDVAl83zq81HNIWcco6Zkc93XQbdTNG8WjILgVNa07
vC7GXnQ1XTjOdN4NiXwcp1dNpR7x+KwBLCb1FVTXFnbyepkyEb/QVCF9VTz/LkYp2T0mRhOb/Na0
s12kwiuuwe36EHM1T2Fm+r1YyRqGylyuTx7KFTvBbSYOaIxpuAMsVUMso1DbJoNEkduIOwa/Uk/4
RVS1Y89xcBz/hiy0xjkmnYGWA7/PxDi9iuei8UPy5vU7W8+nvnYcYPo+fD+t/d9ZiMYBVPhgKV/m
e059BzX64pZ4DSCGdCL291THKclXmed4BnZVfFmkGjJI8mSCGDMw/EGoXdd25ngpjfw3sKKlwQLH
5d8Fz3nnwNv8CnVIonbyWuCNStjoMV3d5cQrk/jRr7XkIK1o95jO6Guo8tXA2Dzp60V5IwB5jJsl
1Mi+iR1mTviX5PJMahOoSDk7vZrOmjhJDRHB1izM1UqYVgnUtnK+7jeFvlgIUIAmttMO+fmYpW60
QOjX0DQDi2R/zw7xj7p2ImaXz411cnDtYK0Qm47UzTxqkqwvjElUV2EUa2TSBFZ4gjNsuMMjh01q
expsqPjVQTqpARXGHjvSOljmDSOGiZEzMuRNufPBuo8+R/MtIdpZv40bzhkSK0qIXfae0Ze3sLNy
0hOXFg0eJ4naid6ZL5GPTNlLuYvKOcnqykMr2MjRwOOWckhCcd1zINtRPG+cSuFxZlxmzeSTqvUg
W05P0d4vNlFQMjALLz1feFpBXoIi3yv0zriAm9YlZ/W/6nJkP3bWojEx37tRdA0Exl7YzkgAkBwz
FB0zl6rJ4gCNOyl3ObaAOH/qr9mZ8qwZx2sCfvw3esc3lzGlcvV7hb/bp+fo2MXHUCrgK69gf3L1
YiMUjz2jyRw8CpXTmags9sfPCioQLx2X84WE5T1xjeINpwX7OwIEUeCp+ZYtEvk9DmkeW/G3cuau
DmWSoWCLeYultVECXfoxgWT7jIGLI1K26gGxE+a+vD/Hanez5xDhzYa6a7lyDuh12E5kcNXxeqMs
Rq0WFjU5ZTjAmutjScYgze/GeDjIl1Hu08wy1KKPns2/O6da5cZPI3rLWYU1ryuv68nwvJfAeA4A
eqaVJ4+yn21k7bKaol458IygONK7AzJ9GmEGw06YM8j9uocNPRryi4RL0yBwTuNkOORKo9bKcIzg
qpTspqzJX41tDWqSXdJ1ElPux5m37J31xuO2gmfSl76Qesri4vugHADEcO3SwBWHq8+FVN/ZE+fd
0Lm4jRJn+X58O72Ej2tXDlNgO7zWSrY61dx/OVydW9/gY9PVPOhPmV1CDu6UUsqAmhAf6MYICvNt
mGfmAYT1C9M1ZwKJJ3NqNUE35QnLPHiKIoNJRyswNuBYJauBkrCVyLSdNacnA5o4gHC+F8z6qA/B
RW+BmpuMaMcQe8srQhb1wfPZqS6tkzBiU86ZKc9eZouuug2Oyso3YoIfEFDTzDRYkhKoKXRnGUJz
08Tw2uC3Lu02hD8OQa/yPpC+mmNAKhOK/3BmtxguibeT+uEhkXqW8MqKZBx6WBlLl1kslC/IfRwZ
y+VeCTQ8pxKcfP3peWNuNhwjxgCaBFg8LB66YSSKNJT40Tc7QAWPlmrY0hfcPUj/b+rfK2jEACyf
+nZy2xj3BXRltPjr/AIAJ3PuoX5PjAzOgeGO3nMfC23y5chYXwbCOWmyqClFMQruP/RcaF9aE7MC
0bSl46+8xDCIBE0vGSIXkPP6LK100eDzJBWUHKwozdxjQtlaatLS0qbXAGBJjIo8e0JjDJ0Dh2SX
8COoP3tNN0NbEeSmlrO8ZAUZ4B8T3LYO8xQXPvnokcyvR1m/DblsrSmCEWx3TNOl2RxD1AaJ1Njm
eDIRMwu6OxhVdbCK0h58xyvMKvKdYPDGzWQDXpEuVSThT7CHiNe3d/5e9d9S/CPCsyVVHUl6S20c
bqhgZ8aHq/q1qtP1hb5PxpvE5YuGhc9lF8MSRptY1/T9ciF5XNpN4M25LOSjpe2tIVSVy/2/1Upg
av4GKrffMpcLvsvhNVsdiip+BsJzLpKkdBkltw4iZJI1ySqsqADWZtdgIc4RMivkSiZxWlkWT//7
hOXnPPlYI6kc4J12WDf2brKJxEAmrR7b2ucqaoRTSbeY5HXCF5MpUcqY9KjI830caTcQ20Y3VqtK
lUOVMM3+b21b3QUsKY3WgPZCvd7UHbDcGOYs8ff7Ug9pYZhYTaT1Uax1A9YwxZpw2NoRVKrO0QO8
miUo2njSTPqZeoKduJFYvi6MnU7dwWZpysN/iHtQxX8BoADkFMdVTi+HK+eNCAdt4AO2zu6Zj7Tl
gDkvTEluEmsKCJ8jKjVn+kNyJwl64LcxudygFTzuDBFJo/V2q+e80pdZmxtVmuPB4234JDMQeF1c
d7ZYYR6FIU+4ZhugIGWz4Sw2f/TsI07W/OTuO01BDunJ4NrUqLkRu2c6JGtA2y/Pq9f37xWSfxNY
ZUbB0fIaa30ASoGru26zt1GSZR2vVfkG5QgVQyxCgAO9ZFckKdDlgPx+mtXqgIq8Z+sV2Zy2YT0S
TbaLsRYOpSmhL86bQk5oVxi/2GMtqHMe0fdTFBhvF/12jHvvjEJgKMXLiH74h4stgz6tJDNvNLYq
1Yg+C7IWnqmAjjlEVXiibcCcVEu/Pgxk8DFITvsaXV1rcGgvmTxBeenDxM5Ol17RPA6j8P5U7ZHS
IETj90A8QtGa9VGDxr3Qpj1L0p3U+PpLzrkIj1iAj3r4PVU7Y5qtcCP7/Lf2na2kuZhN1au9ESqY
nJPySNxoDtIduJ+qjPfTSSs7QLYlhfx27mBO8LrC8oLqANCcwNDFNseB2zwxzj0XT5P5LGUFG1sQ
3Ju0nKDtdpqfjNRgjtP79wuZ8MCPxnS4M+lNaGu+PCDaWbEXpwJblTJNLAubVJE3v252AC0EbV45
QE2MwPUJ2n6olGWjz1WJ4LMQOVYpaTgMuNfsEZee3Jyp57HAjTK5rj9eY77l91ijGEaWNYWRfXC+
t/ameIrYkNiG2MHhxBbMSeuM2iHJingXX0bJ0k1LNeqh/g0wFMpqeCL+URgwcRUIkkiQZGBd8VDv
zZxz2TNTI7C12sh5UAZ5IjI0wokzeCT/SfDDANXXOY1ieARuI58R72GgV2E2fsiOoo50aeoXSBl0
GCyeOctjBtn5yFXQ0ZwnF+4gKMhoG3HBH+AdIxsBYCaa7cDRLmdK7jVn6z39aLJsm8Z7GrGUYRNc
SuW0vYk33d1obIhKhrcDozkmpNch9xED1adWWp6ds+X/A7R1iSrV3z0eVr1tp6fEMGpTguPSKqb4
fbI5Zc6jYm+t6NItrNOqhItsBDHbwUUI2g1J2uTtY1YiCfyxKfjUYfM8jKud3nHDtOcpxLOfQA2p
u+2DTqba58FprY4b9b5GSgpHWkpvDoYwHWVP918hGGLnx5EHnkhBy3gnqVuAOGkFs8DOrAzzbgaU
87lapCoGTwsc/GWPEgADkOF+v9+owejFOfe28pcYNarIffVD9B0tIhqV1UXFm3Z2pwJli1bt3NGP
xgEltf46z0/zvLLAqDioY56AGUF+mExVTpvukYnRnKvtohRUC4iLoondnKkc3IOKXOO044kaa+Sh
ICtffTL0TzE6sL1jhu8fgTlDKJf75enx7FfzeENMLuz1vNVmmqBdZ4pHRntu+yOrCTu0hr81+Wyz
Z3gks5aGzhruV0rLZpomYaY/+9mB2i5zr9IpWI5cvBJ8z0/MZrPeTRxWEDqfATMlODm4HQH8m9C7
o+zHnHLU2F739yG5u7JnhaxY3vnMuVaR/dbJlfB9p8adFAHh4Dn4ik526MBHkAaNLGmCreIv1u7y
I73hFQ3GMcwWyIHmMLEV5Szm7nB2wK5mm5xbtBaQTSgDI5wTCSNSPkU6vRSKva9XAIoZQXFrmUzr
a8P+mgWNp3cq4LAGR46EG4W5v023Cd1ZljNhYcAus3XgdR15Y/esE70kgKeHkMbfnCg6M+Pcht+z
GKP6ppaHMQ5CHoUOKqlpaWBYOXL2p+xmOPbzGDxp4UUWTgk5kpWUiF+xVm3aVxUI9y0EH5HTBE39
NsMX4Nx6pYuAjuKN2sKv5YkRbAPNeEgcFaNA28+xDKoP0MWTkpfpRouxqV99CqXPHk6IrpV7gZ1s
1+0c0EWjHJtkVxGG92+49YfDT8IYKzWoxgT7hJkJofY7dwv9bZfwKBdFo7umu1SP79uK7khg66Mk
9fjpcE7BGcf41aqC7HlX8RVHaJISW5GuIeJs89V2Pad5AERwBkhKT6mbSH/2sBp8hbDeAApGnC4t
8br5smChUEkoMwkiwFv2bn/vd1L/GYQPbWOdYtJq+/rnkBqJCTvIDBFW1SgpqieEhCNW12D+QZX2
A/SG2TBahQHF/fSlxJsf3WHc/itfrPuK7MVxKpM7oc1OsM13vF22Xdf37YCUnTdzGMRfBzJBAbVd
HS9tvdULQHddxTWla0ZEUcZM1HvbJKW2433xPKfcJk86eIqfJghJ1Ll+gS+htr04RqBFUM1Q9Tht
EmfNxr5h4s34bCDRUNua4w1RxsNEebfVZjZLE6+gWClYL4yQz5RtNV/d7ijy8ROCKGMmJEF3drue
ItGMcWjokSMGaNk7KUp2du+fE+9roULrun391mvC99y/pBkG97Y82pme6JSIaf65zl2NRt+n7jof
MZw4DHB6LVVw+lsKnOUgYy9nF9aYvcLR/AQ5pKgbEe/jUjh9P5BtZdeEgGXk/e88cWrlhVC4Ukes
EtTj61G/xYJxTeDJ8V1Disl6RRJEOgS/ojDICOiLF9OtsKEC6W/jYKgIrLh7JZqVRJXypMs1pimf
qdiFqpYqpqTVRgn+FimmCj5sRx+utC30TSSujDMTi3vJmEABN+I+Gj0IhxIx+iX1XXd+gBXUdjUS
hLmY0dhrK2xd3pnuAeyrxYkwyPlDZ1btUI+y9Kwxrx/y9bpCEx4ZRCR3Fk4ZHR1BkMYaB6jNXZPI
xkI9tyfMQJJMtgrSXpiZLeKD++fycTVbSl2KuGMv8XkWIqWgoRJL/tuo/uqq/aO9Zowo/5y2GH43
W9k/A1EihqfQILElHO6ef1GqDJJX9oWQymdh4sUTayubGn0aeOwvyxJVByZYkoiv2Ndd9MLf2yrQ
CjRmF+PoQqJdGYbdFJBbo3h+SEuWanwAEAUFrDPt6OciayCHqaAG7zeULhy9zKFCJLvCyFkLb86Y
ptYuuMo8a2kj8TTQjo1KhrCT+t7lqDsS/O3s84OrCzjRShqXmau1UEbBRrssNgnXxhTna9xNss+7
or/+4SGwaQRcLiW8po5AByKX1SYCBmu4hg40hfcSUPcKVO2kgA5+ipAfYz6kM9YRxn4YJOex2EkW
H6XSHkA/b7HktZQ9q2bTgZNmpGlOIkASFmG4j3K0gzF+vd4DQYzALP3SD1rK0KxoI9e1XhY+klwC
mTHn1Gsu6VY1MV4dD3ZkhIqqWQwGge09y8q9/ydNzfhmPLOOckWAW2HOwmeepCY5vrdHB70CyEAv
HDQTBXfA/RSe2QadVam8/LRbIIEkYQKEHL2c7IzMl6hyIKUZJRj5aSodnzgZgtqJ5VfMHIFlJB+7
XtTVXrMnhkARHW8tk6psonPI6AQBxTg+kzTfO2ecIl74b34eunNFsim0x0Zcet98XpBLa9O55zPC
Cw/vm2Zdyu3pjft2mn/ujfRxyiNaLXw488DsgMsYeqlUmBVqEB0JA3TXe0OIJ9sEhnnloA8ZtR28
An1cCsevBbIUiaTvzUOybxe9+z7qCIObVNeCztOun/NacRcYQcmYdsbvHcvFl8CUSc3mFd7pFHyk
3jSwHsk0gYpZv2S7K9K0PoU99+Yf8SI7ajIZyMPtcuBRMp4kTgsnErhEhXAJZ0s3DjlBhEG4u2ob
OMcjXGaOZ7qmIye7YXSTBC9d13Qzsl8fdG+RRUUaedGP7jIEDwTTJqqqwSs09VDBrtTFVpH325xv
k7K/J/b2S1tsTdjlWmIAfqsraTgRftSzA5lwSu3B3aYcjiq4J83yUt/RiTu8XbgFDEHme0GGumL8
OtW3apgNScGRpaVV9CXiHdykD73PBx2ByJaYWVDZH+5aE7647K7YYVitKQz4WG1GxQL3cghWtZg1
IpuEyWkBkAlJJ0eIckeELnV4lzQpcktiF3lVvX4tOS2YrcdVW0bOXdJqjcAtBUHRBF/ic4h3f86W
frMdm7lXhfmCmFL0ZQOvgRVw2xPbyPlj51XBH/CB1fyf4FjHpqGisfzKZXsiDQlNb/CHbN4pNyGz
Z5Qw3ak2Dy80ruMUIjDzbKJ06c6VKXSP5DDZTU1DqQS31kk5EuHewSlMsyPQELOWPmMDqXzXfC2P
gWjC+UpHrevzv0ASEjujwSj2Yak1YA6NH9b44TXstBvvsXO6n2RVrA3Q6Txd8lKK4ZzTRHV7B68I
42WqVTRoxCCunZo7ss9hb79x2eiVWMQMU0NaizVFNhyE9Lb82sEgoOevLroHqNlHS7v8fsZ8PJVs
cndqb+DLYN/Ocz8BVoULvFSA3+C180xMvsJsdL6I2TAMlb5DsHWQjHpoX3XgnongpH/3moVjRn/Y
+xp7uuUh7LGD5mHIZiE9tC1/IphET+tFJji+og+pLMI+r9c202gRWpZ5NMsMl8IMHcbAIEMvAvxB
tTU4EqRswnHbbQVg+6FdZiYh1DBG2nqFu/CimRlw195HQ7lPexsJ2bfm2q/i3IsH57hZ9fOqcXpw
fPzRBblwZZyNyCW1Yts6BtKgPvGSp9Rre6a9lXrUEXIWpiL8+xVOEUJlfKGXQRCuZKNZWhP8NLBL
ST8IQ6C6WZUYXrZYf/Im6y8BgKw2X7oVtabJQ7XZZYMWg8Fy4mhC6mVoZl1957fgsIQucc5ZH+PA
SnoA73r5I9KO4mUv9G+ftpPxM/h0aYfJWK/IGXz8c46cZDx6S37l4/nML4bHj6UMUw/5GsvnWH1l
C8aWZwoMnEEXryH0Z/OKoZVpVLpyzsp0a93L3KVNiImsebQ4CE4Ly+4nZ/jCoZK1S36O/foxzfOl
UxS7ttfaF1bDiPWpGzd+TtXuucX2M/UmkjSCycJsyJYdjS4umxo3a542x/ZgoK4hqZ4YZC9agisH
S5KHusv0JsQTQYgRVRscC51SGdGyW3IukTzPf/qJUsnSAhBopcxFVxNbp5xMkxN+kcLuNqGf97bl
FcxY8me05uGvYnuPrh/To6da5npix/RP0uwIgtWV+g/FtnLfhpdcNVnx4yH0/NOeVYTyIcgnQxDJ
K68ycZkNbjD45lG/fejevpS6FrD3AQyGIQlGwkOnYyXtsfneTXQf5wZNX6ha2SH8OX0S566xBaGZ
6OV5dVqDPIfaLXkl7YRj4EbjfOsphsbZIYCwLO2s/2+GQxIUvKda0WE6smzyo0XHmXwOOHewXWT+
cJVXbhqaMaOwZ5xIXarRZGXZGbeeJ3QK+sCbZVzdtJld0Oq9dTTGAbkolkh9qn/u8Vj5ZUVkUvub
MMQfXxgzw0gbdb6A0tdZNXXJuNMGnR0zCWQT5lr9xDJuvyn87lqemrT13iTxYsutrLRNdQvO/z/G
VjiKS1y4TnyKZpgLFF8cLpGeLpXRpvtuk69jdpq+VgOmPb5crQ14utfUCzrNZbDQYgNwu8Qw97ez
cXHSCRP8GfHvHgZLQdsQcmuehYmhmY2Zo2SjgzZCB4/uWO/dBTV5lGalPGR8T3y+SRh6XWRJSr+F
oeLGkQd7jkhAV2OuqzADtpMLb+SLOe+DfrX7U+diovYjcstCeNDik+LStTp1ui6/4M+ReKKDF3/K
NlycV4bOYnH3RH9duJdsb+BWKWoqitonbFDnmwqqfwD1EBFaayx5Ddv59ZxcPu1BhuhkAKf/8AgM
ZTS4dirYza6E/s/ZtepPqK/IbABpamL70KNcOf4hJbpoEnp+kMbCOzjLRldD4Lor5yzx4dqwrGaA
1SYjlDUSDWcSCtwBB6YyBPjssLlVAkjOBmKesyEbljxGU86JrHoKnm3CuKBJ0ydo76c3NTbWFail
qOrzBX9lSDvAfTNPBdSyspyR1lJWO/amR24PChPQ0Kf/8ohdXaeYdQBcOT64lt+uX1t5PvtywNxE
5SaWSiU+cSJWS+ltUqHTQRsNL313BcAPj5JOnmTwIRKU49viiSuLR8vwGkIHvFe5gIqXs/CYSVTM
eteLbfvFuIZw4z1KPmtUsQup5d4UFtyfjjxAkBDVeoJKusLucsON1nMDRmltzQsEER//retSx6UG
Z8KJ+wFNJBYvm2BQdMWLnjodybIogN1YMYtp4McACRCjo6tB58UtSKtWjeEHUqIzu0zrILQ8+zjn
b8NOL8bk/Mu4L53fM3TDcwZxDJoOdWvcFTRCqE2+gZ6XoLhqR5fRnoQIdqYksRcxnkOqm4+IRnLj
irdiaDH1pRUG1RjulsfpOeHiQ8MXeCdxqK4b/d8e36SFKWqiFkCkc7xBGCnDRT5ThqISDUBsljuv
o0heF0l7QKCfSWpbcToHgRV/1hw/OPyMwMUetYnlU46toHsulAB9cFIpAbHBbdARksTJ6P740h+t
V1wJyea/W4F2okt1EHyviyN2V5GRuKEgYHguWdGJSzNukbaDIIQf9ObFJ+Y3RgmxJ2KrZeRy6Hl6
Q5axGQVNi6GlFJKTHJw9CYRFuw5y8kgYTPBcIzNMuRMgwEv0XMXu+NoitR59zdvTIjoDdux5Iap/
n47c+/t7o0VjoyW7njASM/aksunFjgEtpap52lObv3tVLqxos+NriFdcCGC8W874RQ1HlvnUroi4
3Rkr9sRH2nAuqQbq+BXsyIiX2xqQJcpclqGoReR6TLex4tJ/Ykfta0L+Fvgt9ENCIqrv4jTksGEL
zx5sPWyxW5gNaypIUZ2L3gNjAutMMujjfAVRe60e13T9ieNx5iINhOrGzvWX4aWD7i0p9ZVqPY38
xjjO1NvPTiANrkUlLxQdVQUwM8pMdftvMPsuiK9ZBl/WW1KuTNJQBj4NvlVeAh+DQH9zAhkWMTWD
jVAlFNTmNM2KzdusWEmx0ts7+ESGGvHl0j/KybGKUqy2OQ0mY3BBSRxm/dDFbRMqh+Q96J+gJLwn
O4fOiACNUsH1YsmW4UVYf4o9fAW9SjLvRH6VN5KR4Uy+eChqTPDcelxzNbuKLbPyro+YD091UO8d
i+9PfL5k3GTQ7lCa9mJMQLsE1WMPL7GuOEZCjlxKOW0nrwlVMEdsPayiuKI+7PEb20zUZLv5Wn70
HwAo6xq1rs6sfygJseoS1C2/azFjAZac/sEyjnEWiNFI81iQOxUd8+L50ET4Us+6NpwTG63043yS
bZQSEI3oUT5G+dhA01R5m1lVzigIImUksVaMUqD4F1J1+SRiteZ18WbIF+DEg+SV6gFaqAmMr31d
EAGjrvEnBQXwBKWgEVGDk11WW6EnnogO5PW2t9IkkRQn6JH8HLHnV/qmiEHNyzQcEveHvk78Ssol
pw3hMvk7ZtTXTA4s1MGlrmggWyoluxjJuqWVBZ19lm/HoB0vgFTJMDbLappf0qz34EnHHu4mJ+oa
qxFQgIohlHmFkC5nfVYF7sEi/k45I2UCn2Jd6MQ7+w5QS7FC8DKCgEjL3DVldAI0vdjm8Jsvs7kU
+XS45ImWIR2tVzoFG87tROT7FSlv7ecalMEHpVNYSrGocPP7NOeLjvx3bqm22V444/ag5RPy7YeA
iKzcMIsB7QF6nycci/Xzzw6lVnvTeNHihFQ/if6bNiz0q8akFsf/f5fH0s1u4nKnAqSBu4qWoIUF
QTagkYT0qXG50flxbpxbj8nF/UbvhUYzyjKdEakiICmcxXU/ghiaRTg/tdMLc3hQ9WCpmWu3YKca
YpK9QTiaV0/cgMxUV0aacVNX/THHfhHdm7TJ0YPaxtvkGJd4LD/7Ps3qvHYCxtbdip9ylEMBrIbV
6X+MrX0s3+sHMa24KgsVKMDFuc8ao2o0OwLgBtoJ7lFcHuvymNjOuKYcXOXpRZ2eEWBg2XcMPwBY
f+CWUZN3ZygB3zuXXg+WUqYK4rWOv+SR89m9APWCq78FNa70Vv1vFBLJwlQXQhgt8Gb2Xa2QuvrQ
d3JqjUwiOpPTAEgdkLmxIfPfV6RtbWrhPnmtzAAnzO0HIclEljIRRxrhDI55E1670NrnZKBGuQOf
YB3w6j9la7RQWJbKxuTkvL79YUh2R2AFn2fXqPy9zWIl9ltbzICV6b9UoS8nUk3mR2muATsPVCbC
oXcylsulf8La8YgitvlobE5v7E1xNORtBpWVweKz+b4bgSf9xsi6mHYWwHUxxkPLmEoI1a6PTsYf
/G5dSjdIY4teFPgOeN9zJzrWqWE5Ud6dfl8kJpeY+TuUUuhgEpg1CYUabztAkHurjXaOAUM0C6dO
a5QHJNUu9cPB0DKTfYZN1Zlsp9BedYK8AUSLoIzqUx3RyL1IY8yhjgZBwVjp3+wjtncHv5ivUcde
LcxXgs24pE5x1A+7cvdCf3tDPFRDFhkeX5cEWAhvl6vbMjHBENu6rHAb9lGCkw1Mn8rWQ0VicQvz
fWJJLCE2pp/OoHQMbtuOAFb7JU1IgHs8xLVPobMvCEnBP1B0WwnkGCxuG4zmFi9KepqBDJXeMj/b
0/eHuIc83JVj0KizvNBL9WRU2RQuwub1GPhYnIPqI9dlmn3vVk6R8mGTj5qyCF+t3nJG//A7P24u
Kw+e6/NmAXYgwZqa7NHgsEQILf4C0E+28+ZFiXNZQfWoWbaKXP779qFWzVjIZ7BJiWFVb8RplAem
e+a2K5sBTM+THQO6di2IjaPza0tkbzEP8wCs183GDfBY1BB33kmM3VbihIyDiwoT+t40YNiJPlER
waieS9ExC6RR06mi6HuE1OrciKDhO1OjeYEcR/3DxIWMhbwCGNOz18UpLKFVWKYALMIvKc7ysrki
zfQL0Z5JF/1Qsob3PqL04Mp0ixYfyya2brIKg66V87S+ebT1FX81PYt85az8HXy7NRoiIWAXP4CD
YDdNLWYqxTZt1Hs/491J/LwEYtudkThIFumI5P5XgMpIl4Czw2AUF/WQf2Zwn+A38pbW3epKxnV6
Omcfw8j5a79TaLU0zBQAIwaheDT+/uNJayTykndXYVx9ETeZc+tLJWfrYc5xKdLlgEg1K+Y3gWJE
9ubjVgN1dsSj6njrtfyG4bezo87ldl7na9EQQ4YIPb9Z4gRllYj26qWnMwL71iyYPBUd0nnDR0fI
XTtxvoC2eRIe+MKg610Mlvu7+vKQqALjP/tECVdlz+PQVMPk/b/K0IINLyWi5onpRUBLA4SAiWS+
xbTNTXtz10cAUQFgS2eWLFm5l/KAywKUHGo6p/liM8oAkzB2b8s1/g+jrpi4R3NZ409oV18Q987q
lk5EpZMzUhhHTm7o2YDMp7+MDSmczjacauGGZ9UlZ7W8p9mQd0YR1ypcrIEVvpNQtTKLqnQTYSSY
fvDjhbii4kCF+MoLzd67qei7I9ZubIlAuai7tuHcAAZut3F+LVDcbTBxTPpZhTIbS9IX5+tCnfvV
4cQ40/ZTy+FLC+LQ6fl49KdflbFJmFyLVRFxP29wkSRQYJST3lppwGxko9ZA84xl+glslmEXorGb
jsA1IyIQ+IPz60OIzJYXlQTj5NGP0IjU0MhGkLn3IW6xOvZ8BBYa/ygy4DbtixT08U4+8fnL3m/G
SfI8FeQkAph2RAXirmGcBSLibyoCwZ5j+Mt1KNTSr+myEoIoeGuUMzR/ZN/JivolcfTIkjQUr0W9
xgbvESetZm/UgtPVQZUn/dpHnt6WwBF8Z831d4Ex1QMO3qXklb/VNNj9JTwGPOnfOgWFPogESvlg
Bh+OdP+RzIx0FVRkrR4WBWUDf7yL8qV8lc9hhmfZ90ZSvdLUcfd+9o61ChCloxPDAJ3ABWokF7pF
0aOultWduAHL9/6/kVxbwXoKoZs4x7QJbzq1GPWtltZmiPRCCCN104OkaKbr4IjLa6wIJ7i58SCc
zw+xN/LRJL57bbbCZfejfHguNUxSCGgYQCHQr5hOuarV4lf6kKLocJFfY68q7ntI4G3wnC/GO8sn
btEMH1H3MO/9/WZ1MKElOJS71fU/yLm3bdaqNhgH/eEPlC8p/nq1rgay/EN6Tu7g6t1mWQAZXJzk
PgI6NcnuHuoBsJ3f5EZ1a64OmH3GdNOB1NuT00mlRIKaxQm1rQ6CIigf2TGp2yqdt1wk6nmSK2oy
yZJuJ7ynfeoVZ2MuovSz3IcXwlTuBOmNJmtje9iO6s3Lncx8MyXLUY8KzgnCaXcB+Rqp7RxpaiLl
NtzqHgvh2uYY85ND/SCR7Dk1LEHZf9nHBi4+Bz37W69v4Y/f9BZMBECPqlsR/pz6AAWk2EfZT+PR
ipCjMrzFKGxHuxIsah7PbkrgkMsClAlwICipshZgospxqCPVCS6G71Q2o1TsEEhyL/pYq1wDp6Kl
ZCpMA7oixTgxGu6PxhbPn1YvDth03Y+RlqVIU98iwwp1bhtd7ZaE0A+grFOwlD0kiJv0hYkB61kw
Gq+l8Ge/jBbF7h8ISu4BbAr/cY/axyBCd+A4qubkWuHrJVCY4AWGB9y3LsF7KJw7536GMl/cDiKW
B7OIWe8iDBpgL9aUOfBLPoxVudKrCUKZtnyPKsGN7wVm8T17z6DrqhVLRfuD5wI1BJ4eb2su/HuG
FBl8TbBEeRXOEDY18jHiS7ky338wB0ZfAQdmNaRnaMvkPT3iS9v0svLOxr2QIkXYVK80yRUcmqa5
gFIA+DRJh8uHI9EXSzN8TV8a4OLAozNRR007ASjkf3qtF4wyQD1Ktz2zjGSDwWXleV2mwiGGw+sX
YxzsQ+j6AutAZ7h/8j+t/QKju3jh75I9M6X6RtwSLUjzTtXPR/lKWQ6mji5tha7XVGgFMVZ7IboB
1oTLKoQXbE9yJsY5+Bq6NUTQILWioSG/9Bn7w0yBQP8XKOd/RLyMfGbNTLkFkVYl2wcogvSQlVXK
qN8R0E9sxLsVaU+On9ZHJ+8RnmiDfNNZBhWNh92Bg9Jqqyje13Trq4OslLQw33bn3/SKeal3f1nQ
+d7CzJyY+aoDG+cBR5afwEBLwIfxTeddaFsABTtaAcP5S1jrG6EICRyEu5N5Q51dnUhx449MGPkY
DQyR4XnpE21yYWE9zvUUePN+XCb9RDiP53LvT0Ir1oYAkjT9zW3XStYsklr9Nk8wDBK0VcufIVI+
5XGImBJtwNLMFWfzIyDRUDyvcwjfz0CND2qvD54ch0H+0W0MMGFFnBu6wr6g5hkcHyPISUL5PJox
4otX7uRsWpU4r7CGDOCNXyLf3XIwC9D8qHjkPStk+XE1irIrsXYPg0kk1MvSgdYsPrwsYGb0jcOg
o8dtbFgEdt2oduM+/+1p3e9fT3LTgFfM09JjzW9a3C6cgvsrh6PdMuBoeeC+fj3+y58JiEXTr9FG
jftGm5O+VJnkTYW5EL3SkaaW7436e8fFY9JiDXzAGOk9rjqP+OEMunycE5sCwy9Xw6rDxTynktMZ
0xmlH4S9Q2mhMoaFHIUsGnV6aMU2Ws7S9q6iKuZzf+yHwH3t2rEO/LJRcqwDhYNG8KuWhikdkQuM
la0MRqO9so3SGepdRgFwcQxoQ5aKFus9QQsDRbYXBg8bF2oEsxl9Ypwz4vBcBURjXUgBYKZpmz9r
fkXZ9OARmrQbnw23IPxaB6rYJ8u/H1sPF/sdbH/FGKWwCTJe2oys4YbTVirohx5RgFladvwiCSXO
/sLRUkPf6NsNGqISqCQM/WmiuoPPPYs4Fb1i0jmDdohbquv8Y/Tqoab8ar6t/wXzkqaB1rz3B4Aq
zxug8cV7Xhuamdo87LUyzYrrqzXPovHRqC8ibuyJIGJ8UubJE/BreHvld+LfVskOOb3ChJ50SUKD
t/G2lP+5jW93m5pcAA+ZC5HUBuLm4KCKvp62/FzL3HTqIoCCzgZZWAMgf2vsQpgzamqkFpKChHPF
lh+atpERHxJNE5UAem4WK9LeLYlpN7RwdaTkS7BcVA+1jFVGl3IaoaEGLRJzTuHQ8918iU0z6HXj
LlVjKmP10sG1fYRZIl44rRQB22Gpi4T3Ym+QnEOlQD3pgJFS8sOszdzFz7brcLfguXECzBsR9e3W
LijzxeIhvsBBvnLrXoU7XRgchCCp7vCW4HrpJUS/lLu8nX/cN76MEl2dKecEIayZWjy/2VpNfPUz
Fa41JE8R8VsnO3WqBKHlxFAxYnNqYe026wOLtbQluXZYZxrQpZLntURBGrse0sN4rXqNrRnxDw6J
UlDzJeiFtL9YVQHw2Fo52bpDL1A2l52wQmzMiT9KE8dLSHmETJQLQ95Q792Fn0qtuSTw3kfPYT45
/7IA82raX+38xZts3Jm6TIh25OpWmdShgMQqD5vtlvOg0/HNfb07YB5iSU71n4JjdV4GZLWRWTNY
YXVM6L/ALDrgJ5P0lBiAOUvCnsof5evvoAXJ7YgzZmgwsb6uwzVfVp5iYMTcn6Dpsk4fvGJ6/ASQ
dH4MITAm/12JIYGUabQILhmjwnySy2dKcnaA9ttIuLp66DBhIiOE5iLSfI/e/5Rcmk+/ZWWslbit
QYEcrW0IXKxWr86/pbKW87fvGDg8PdphQMm8ezaJY/rBcNXiOmBcudiCMnTvlTcRYoK4TJsqHre0
YbW8j2mvJi0bZsnKKjrkyaLeKdibFJ/90Pz3/FRozNTf3uIP9mAgVAaAdgEKKOo58qxQxDKCUVHx
Lgnphd5KXCbM75X72ygE7Ve7tGe0YRRl6CX5OLQbJJl1SUxOCj90v5uon3YOFRSVTBAVIxwW/ssC
I1hymd5pgNazVweE/SNmxvZv/AUoZXyZXHA/a554OVDOJ0saY28Nb00q5VtD8vjKgvvLriw4QjF6
YA+G66lLmtSOY5Ti9+tq/YUQiYUIHMgU/tTR8Goi2kc8SjenLJMwcB0P2oNyvLFnMyiFC0LuLqF3
yoc8awu7pocoPm98rkQhX9VcguJv0DXccXMGhSPTztS0bGRwufpqjI8ZqIlYH1qGVIJkgBEhYBir
dSYPxnJuPStAlHfrIZW73IetR8cdK9YtMrLdQfk+Kdk1r5Cedkg14lqBGWvhxU1Vp5xzRt5tAlTX
3kKj8dLQrx/ur3VMrKUzNN0EIMDB08+A9V8+r68OKhjZ7L0xlodc8Y22JbojlzDVgTD6KZntDMJR
dVeQ5DPGG5RYH7c+GCYR+DbusMYwiEla5n/b1paeO/sEhgPyBQeXssPW78KmneZs0fxOc9zpDUCw
Czi7HMd0IlH4Iu9CySy3Le8yEooVSuBX8U//PTJpqx1pz3uFKH+rSgtA00Wj0rXEE6vFK+V5ZWQm
IWomlne0dgfETpFxeHmD4vO6e6YnmHAyK6z74RfGca5ddZQEdhJPNjvqwhNSqxvZ6yAJonCY4IuF
G53dspUVFMgrfqwijkC6R2211Ke58oEXxHzWbWfGymYabbwQywTAW6g3nA8mktm4obDSI9gJmNm4
czg4mDC2cNxHsTfpBYL6eDJH7sUKYbPVgR0zdXsN/p6e7c71RnZjUra+1LSYpQ4xGlQXCoUrz7nS
auuE2d7WUu8uy3wnQTPt/ffkOH6s9rIllQxmSVJ0F744OsxFD1zlpQJVqIOBzX07brWQY6OrpxFa
kSLxCwbcDFK8c74/qumhOSiPX/8mSzsy4R22QpeAf0fo0uFj1mrgcbEUpewjSJOZy3LUrjvDvdOT
O+/pJsplGPdZn5kbVdR+cFY5lzoyoZHEigZbncYfO6w4Dn2HCSTVfZ30B2qwmvDGk0zVW17EGpXR
q3f3e50Xf6A0QpBR45Rd0y3Hqq3WS3q+gsynBg9e2YDs+p1n0pJXuOpsdVg+L/Y3xIsSDu22y94K
4BX6qVmBGrmrGE8sqw4IxdTYfCvrwZXYYz20ERxKXRWm8kp05D9m+TSrnr5xwE5GxPgtruTTbXRJ
otLAAGtFoNcKlCWGDlox+ea2spBKa4CT2EX54XUZCr5gZeQISImRoyzV5PNKBPaPsYS2xr0i/Uyj
Ub4Yv1/r18J8LbrN6yI8NUSgkjTQUeH7U2d6DJMEWSlZG2WLunbkBxq4UbzREP5StC3MYabu6y/x
wtufGUgYJlWLQm2vcE5zlrUOp+D6zWj5lY9eECtB/Ri2r8/LfkefOy1Y/+ZihEjP21a4uMDc05Vj
lABkSG+qverUieZonhd6LdZsxkiHZ/embEx9NYypAJmPz7NJFSH9OAhrrBWCI/ZUfLxTrwZ0eT5U
HyXq3M40/Ks39j5jXzzaiDmSBiI/bhMjBQQaIvfaKCOFMA/IosjPLSba1I4PXk/TgVwMEDh3sdqQ
kgL+qDEvVMXMkXfik5xgc0A+Gniz7UFYatC9whGQdybc3pSJnzIBdeRNcD96VsXfTv5aguPHK52c
U4/dtVftmlvToMcMS7mL6WBKhJT0xED1rDcIcy9MlVh94kb6KOL3djMbMD+vBE1mOPd5AELiX0sK
MNVDUgxFC9GpxYcH5xcHeVxqmUApV/wM4xwhgEt5nRGJMjuCZI/xwxN1TS2ZMbG3fv1WRkzvgSeA
9IqPvk6/HI4UgKLFmE/HG+zZHWv5YYWAAsIEc1SlqkhYA50TbjfxBSISa0UMTP0kyfI7lutQW8LY
Au2TNiVXGoRrLR0SHktWkr865y7HbuB1bXNp9cOK634Y3WubelQC1TsVPiiG6l6uC91wNMRVfK9c
oyOs2LP2FGtHGSj7X3m7wtDDdGvQTtgbQNDsZ3vc62drPFKSnIbt2CPsymrmKIuJCMK5wdmjO1lF
AgOznL9PfUzXt+x1e8riOwWn5hUeTVJq67twjmcybcUkNifO/6P+UkJCO2CEFRpXVIdfLErJ2TWl
jsHlHAgjX2+BN3FXLFB1lKKtLkukMPItm4JytxKhkR0Hw+nZ7Vm+5+ZsGXx2WpItD0rr5SD1j8Lk
hLNkdAbWmDSPecL1KrPeGQuHXlVWTOKKUpKOEuXIhavbapZ6zuLLpsglvJJLaIyZXHIMCd9S76iO
eEirWqxQFTIGMz+Y2pcg1hM1rGXz7PWKuTXg1bCxdvh5km2SyAfYy0LLCL/M6P+gaPcMLP+mBXI7
xyiXmD8jRl3BuejeGt/wwXLgiNC5EN2qm2F+3HXV9nVZJzzPjjKCvNQJuZUVTOz2fUgIrYdZje5y
GWPnAxh4OWsvgDl2NoS1d10uRwJS3OCR+eY25/7hpmN+4VuvHpuUKmFnKJ8uQbyzfipemjsykkh9
NaF+Bc/pQQ++JvzmXzE+4diQ/QH9Np6+MNnS4/pgtd9VbY/BGLOtQ8bHcx1XZPVckTBDspNe+/in
0rLdRJSAoR9tBLPwWMEFpYB5IvH395tEUJhQIUp+bkEf9CdKls1fSOkXVkJuw8gKdK7JQ3WVDnPY
RnyUAEyhu3BiGVufmlkp6h37cAJY3gzludiLDuL98GllO29mviQLwcQ9rSYDw0eLtJhqUM0ZZCzm
0g255Sbiz+Ip2wLPA6Pg7n5ru6zX0y49/9COF6V3+vhlkzg/vEjZYZISXd8GouAp7+aFlla+hxmq
33WIX/hCeLpFMkpPmv68DIQ58bdCYu5860Li+QvtBNn9VIk8w4w+e/lqWBK3mooaiF+y16eV8Iog
4qe2z2FCKB7roEgVG55XCE+KNeJPkFYPHGzKRV7w8joQHRevbq70oH+ecq8AOMcIEILr6H7iE7TG
zDNmWcWK751r7TB9xAWby75ZXrJXxJ3nXqDjsV4Q0I3hUtt9u7dDtEa5sSfPt1ZPavN3MSlSNeQ5
+gFZmZ1qrlnKGDwPPQDbYFgzsRRCJ5g5oaaV3/BZRwPbv89tSUB/Kk18bv7E76xSEL5WQLYNpI4w
k6v4LpqfDvB3Z4s3Nwwl862wKpY+ZOK8POop7C+AFdAJWPxmtKnQplshfBZHh6yE27T5E13NlIQP
qGpzAU3xAOpGjnWeBaNaV3uuH1OZWSQOec8SvN2axkYLyfa/FgXVKEdXHXTIfu/atuodP8K+wqUT
MRaTbR/OqaDJTXY3a7nNp9SKU4r7vkivOhXLcmN9yQSsgPI8alCWVIbssXqPxD2RnrINPlocg7f5
3OMyy8494Qpbz1Ezcy6ud4/Wdzc6ZMUqt4z4Tc6WtmzX+c9XhUcWKZIiWNqTT3lZsP/26VO5JeI0
K4mhIOfmu8fQmt8V6V4IyJdgqYfcTBZivkr9OICrOOUb+QoUZ86cN4f4dfzfGYl1mZrOsfBecUfL
+RYrvOUHG9+R3HkFtzT3wObESbxm9fR4nWie96GQhDWkK2M2RwdEQT309cYCDuml4Tfz5BPA6I5E
GTGUWn4MmKlBW4oSnwCaK1LA5Y4pqCH8ubVYUkAJQVlXVmXNoh28lgxeo4WsdgPiDB3B8jxSRLLb
0LEhA7q+ljVcAw8XLC5vhJI+JlVlJFeoZBtlKiJoZ3AYe9XHw0DDfW6uhLG8bwsj2qKXdFnTyiRs
n70QWAvL5Sv68TRLbcvWTRn+1+ykzBjmQvbvjqI2aa3+f6OFN+eaalKT20qc/iVvEnnXMmg+p50M
jFFyPznuyHL+E6AQM2KQAq3UsfOTvLnMFREksUPcARKUDpAUDaJXka67RtM/u/FBodVyxawivQKs
dUlNDJ4NimSCRDeEgddLY+OjGizXSayeJnZ1A0v9kWTOld1YPH9VaGqHZFiwOUlEiQPCgBZuBUUp
6uXh9WIDjhl7sKVqZC2QmaSDZzGybhYAgcvjodgi3pV7qo7CqYUhk2rR/bMZ0xXiLwrbLkIlJlk+
BxhqSdIgZWHYoIT4y3xkRr/I+x/bIUi3dZBdn56HRT+Y3qSeklp1l28M5zcyLutNvHp2zDkSA3jK
wO+RPoaRpX2DBsg/oe2iZVh0R9yuResPqgTEXA173DxFrANz8a2aVTqwge1YxPIVgBQH4vRoqFnq
Xu6DJkztKu1CN6P4Z+Embeuh3F+narnWCz2DkxhwntPOeHVVmpZ30hMouiKgD8HkojK+r65q+Uiw
simGqzV2SHBACxS7j2LfgFEXozixnL9XXQ5TgfqUe3QuCIJTjtYxBvjAs+FyeFeKE1lu48lip/mX
XRTkkALHpzbxtdVKjikXovuv5HUUZpmW/ke2IIqKfK/9c2baiH3oF99Pu58PEZpfho8ZTBHrF6T4
l2O9mTZEZsOyIH8iGAObZYK+hjWZjweSWGZjtfjCkwQsIEZsVK8h0x3DIUhgMlnPqYRZQMq65S+d
qjkwVwy2/9zr8qVGQEi0FJD3p+6oiFJm+m7rmfzGlv+wG/DQNofx4f1lP6Xg5s4ye57yD4z0MojG
UtrNkGmqskQt5E+Sim+ic01WaXR9qAnHwSxeQhwoU1oD/4L9M5rbEBMuaRNNvGbolG0/bJPlBFAX
jrp9Crt1w18RpQksuIkRl8HLAGOaEczKrEzu+gYPUOmTx8MKGEtwIHQ4Foh3d9zr1PYMf78UaE9Q
Ci86JdqoD6/IiXvuHpQzEpj7BKiU6Z2AGIeSoS3BJDKzl0SmQTJ9o0ZP15dehpPzrrA0diKCv1m0
rYjQHu73qBv+iNEnkqyBbPWFcWXpJfdfeM8NxHDaaxGtDhGcZrGcM10wV+yX1ZdUJiJxYOlVQYaL
H1b5J3/95qbHRDL0WFnV7cHAIbopCI9FNJTQEbuBkBI+I4afSYp5XG9nQI9loYPt4mbPv0eO+MVb
4aaOtGDS4XCfw+JuzSLiNkcVrepLLROWmvsld6X/QlBr1blT1/AnKhfwS+uT+yUXLbP1wWbDZP2T
l3DgIzYB62rfX79w2DmTJYr++Z2SleZA6tSzSGHDO4BxUXdAO0vlfSmTpipR4gAvbzmjNFOT5BmA
q2qhL65bEixM9M5C0sCwh64TSJG31HxG8lVbqN6jipINQdRegInNdq1zmX6hGJt0fDPEuKKfIAxr
TG9gnj+rqXBbc3DaEb2K6tFF+DQnPT9HbLR6F5W+5HQ9GHAlkJbyY62WRt3Fc9IhTjy0cZIph0KX
OC+aJF2pmKuIW1CIU41cF89hIwFCpz0n7edBhABIEUsv7aexf/KLAcSkMM/fuejZOAa75it7rl8t
w9YghkFQyu/22D28AZjiDDW/Tzs835f/p5YJRmM4KjQzZFIftXkTWD4Z6EQ5ySdpQ/9Zxu9AZPQy
AlydA7niXRjQoEQIPF/AL/ID69YpyhNFkIiV/ONt9E1JOJbXQ9SHNw2MwyyfQU6g9IY7cIs+H/UC
ZQGC2GcCczIUSIYZFHckMTRuhM6bqF3xEcoJ0SdzMl3MyGc1aZj2MX03Cq8uaSXTbwQ1UrZ5TXA5
udlyzWjo71I49ORyQjXdzUTUJsha9OiKzE2qYDaC45woLd8GDu+SzAF9dIjwZw14wyxkpi3yhgse
BYsTlz+Tjldq8RBvmTHhFzFsDIadMjhszSGaRjwPRcRaMW8p7QLZXGxBAQGl3wyLJQ+/6TEBGDeX
4G4ttUAkIbHSEuV35W0ajGJhbvY4H4K6392Q7E1CY/ggc1K3gh6grpEdXE8QQV9L0ABZEaZA2IPY
l1mk5xz5C0zM4T4tnZEERhDAh+iKzXDg8GkPJNIku7AZ/N4aZF9guhbm9Ff/06IbbCC9/7NWhVjf
W33EYgqTk/QQpSgf1LKpwimNOo/ofaZImfZNkAknDe4BiSjAC4CAg7u8PO/fv0NWDoUQvW56lk6L
NLF2lsAsQ1ZXFWhaJdzC7yTebebdcWPa7lmigWlfVP3r1ypTMLOabYTWSxSIkwA56fz2c0FPR+rk
9r2jAvmsYRuakswYh/4vDoB6N1NKVlNhG2h6RZkaMYqYMyAyBgrP0SM6g0XibEr2MjIZO8yyCf+G
mYIeRyh+Q2SvMckaV2/j9tbzAzHDJB2XLPYsAdYCOWY6kyWpBxFQ4j8T1Eq0ERwnOjVPgVNs1eSC
Y3RRu5XLanVPJTYLSamI1AbFXL5sbdXgnjWCnIctxr+k4GP0jMgd1AWJiahcEigcN19IQl0a/wcp
d9Y5UzPkZ9zdrWgXzq6jf3uQV6dB6Y4onIj0aDPtmG4eV2XNJmGUwGWNK0ZNvfg4sUKw6bUdZSPD
PvDjnfPhrGM1mFBpIeMlvVpjNVmvLuvpxhhBa7XgDcd/c6zOYtw/CppY2Yvc+I51EJRydYsv/+cp
sQEbCjO6uMm7b5sK9oXKp4pm9NnF8oORsbwSyScGzYvp+2xwgy3PNKK84vz8SeLlRJzpYg+CQm3y
HVPibNtLhsQDdL5FJUmsL7YEOehTVGf+UDn6LYWuCsUfBoVHlPLIybC0lBv2kvoRCVLQB44sjz8E
gjFgLyvQLHjbOFKWA+9rZb6hhDoEQFVR6h/H61uqsGz5Hfm3kK2g2jmkH5ExyLCvopvq7PCvQNZw
KjiVXe+7IvgPH9TmCRVBrK0cKG3hwdfjgI9i//0jwP/l10PhH2Zy3NIc277KJYpZZHI4JKCU908r
zmoMDvIu9IWXoWgZrooTAm3YXcSDB44Tmt2VUWQo3QQXMscz63NJOE6JmRjHYSA8S1V9US1+LYcV
IuMxBBRbgx8My1TaOAoF5ZnxKJwSwBr64D9WcQnEmz7L+WLqmDU3+5MidTjol34etioCYMQyBxFl
lb8MG74dPT1dJomqNnx5mQnUZKzY7i8A5jTIsU3e8XNVFQQgPVPdpvXoZTJjXaE9+SkjlEffOOao
Xn3fpy3KhXcaBibM6N9DgmpjcKjEsLnNb10/4UzUOW4BiYp5jb3sxKSkuoLtqccPGXU2vhl8Akin
MLNyVrq7rO3Y9Vk5WVhxf2MCvs0qDPdhMw1pcdTInmnVRcHx8cKqPO1QWKeg71Nu8sAyexwdSN0o
cUG+kN54B3mWZRRHt05alezu+MJH2iPnv6/igpDxRCaVINlr9WNM9igCsEQLC6LuskSfd81ht2fc
rQBWNTR7VQsMi2o0E4rlAhmBYMOdrphtHVkU498co6+GIDynMc3uyo5kz+NDqR1Y9VSFwi5B3h1Q
VZdr86Mz+n84u5+zNjgGHLpgdMMulvLc50oY3WwD86CWvrOuMEW9cbz0WyAefNq59ygba8fbwKws
ViMdhhYXrzHznril5cO3pH6vYeFWDASFmDsbE2Z3oMuM4BroGbdLnwjPVAhKJqJUrSFoeH0AE/eb
pf3Gjt6kAw7JIlY1zJwl74kiDJSWGVC5wxxwj50q5Z+L9qx8vxwE3PrXIOkgg3V8jhcKFY535Ssc
XN+A3QI30Ptkd4NuIIE1H0xnYgoOdsAuT4Hu1chwaczaqI81VwPosVwx7Ya9nMMcpuvzIPHgS00y
jGdyRjJ8dI+RYjukVm6jgVJ+KwH9pBUuqMNjJSt75SLkwc1hDAHbpZ0ifVT4I6YQIQ8YkA60feQ6
/zUeEgxB8sZoG3dQ0qjpwGYdwQCZaz3wxQoIeNpk3vUu+VTWqsubcPOVyz3bQEnekLV8gQ8V2aMy
EKOHcFd3RPZ67LU9i3dUEf2hEoyF6heTQCYN3rCcTGY2plt5oyiMphJtR77KchflExAxV8B3bwKA
+gaIW3BErDwgz4bPpMs2hXOMgkeusOzWOh9DUTPMTB6ojYOhGXaWnrIfrPy4Mmedu+MYvuT2H67N
eueX6YslXerhstf/5/QaN8FXH9D+N8ChuJvDf0Cb4L7D10dlsnj70DKXF1Mfv9umcome7GGCnD6J
EKwoTg1ze5c+v7pe3ZARKZM6OibA4qrmu4tTFhat6PR/QdLcb0D13mzRmM447LpvFdByH+uOFeRh
Mh2ljZCccH6dMEV7fPlohKtYbMl5E7GT4seoChbYtElDIF2rPSwLBGIokKW77Q9Zdcj7Ut1CTy8V
BZDY8diJI9xgJZMpltBxC2jBFqlhHVFME+kHSgfqyQDHjResBzpKy3BaQbVqp8/UrxH9xPJknLvB
EEWY/cmvO2d5IUGaj+SO0/e70rS2L5krUdIyvnYMa67aLLvUxkzDe+mS48XM3YcKAFjT0tU1j+7S
mS5Y8nzVvEuejfmHjqi60xNoORCqKTmH/V4FB3vcx5CHf11niVzMoJKmrskuqFHVmPX8+ahWy9An
rEKJZp8Ii8ZuXp4LsHI0VpiTnJkG+RPYFlp6TA6n5VKE4/jWz6TkyQx28pBLcyk1+6Lp8scQaydC
bL9xjqUVEszuBsx+2qGqpYJPHnxKtQIIPPLtuuLDh+8BdpIuCMtoh+gc1h6UyfxAoB0hgVgtouh9
nR+ADwct4r0sciq7FgJAZwGmyiIfvedMI8dlaJuWpmIDI2HYOUnv8/RR1klbsbntLEfBHFjVEhjI
2Kysd7oqcfoTystysZyXawebPFJkxAXreXCe1+tTnqUwEc63KCe0nH3lME6HLzAehr9OCcMcib/x
+VuDTCPFxwpI4Vgf8WFuj3NkCD7HCCjjlscQjKrwejSWh9ZehRb4v/3giqxOclCHXsjlsbBba7AG
ZQJbPojhTTiBT6Zide5NCHLLPGhy+UMFfO/lF+l3qJfVHB1aaYsSxEFkzjK1imBmIH1Xvbv7Jdog
SP914k3Gji/LYFDwLTRZQaasHoFclGHC5ct6n/VjoWbrgaywFBumOkfSWoxkw2eZPjG7T2YS80UB
WHlU9i6I6TaEogouwV7mcSKx6WpTF/q4yHIQPgTaynrfyNQ/AKsuLfeV9gmkhQmuDFv93JRTO5lf
9BgmQFc7JIHBeJOJKU9JF+wpF5/RQ/brSuH20clK9Ka1Xo5zYcB/o0xREAMnUWcNFB06FsTQh1qa
VoMrMDZiCE+T3fF7Wly4EFJiL71+4GpEzgS3Zk53sZL2DxHZI3hJ/c/NOb2slAkuZ092l/+Dq7qK
4N5y1TZ1bfJUZ5ya21FmL1LykpjKUwSNHau5oPKTeew5NDvJOIYXO3tvyr0+S0K5q1vbWOzbae7D
1nb793OW8FTulAMC/XzCRBUqXqVki5gywo7yK38fIy5aU1gpgquLfnBPcNbCLp+PUFeBv8WY94d/
kJwVi0Glfw0XZ3OcLI6+oB+tkAcFCbREp/2rNP7ghqq3m1dqusX19MEB5HVsiwRXOTIudOxcyReJ
z2xWe/VOodZ/qx1eGqK7VgwGXrpghaqrTl9lK4JxHNxVJ4m62ti0SVu4n0ckcCLGH2uj2htCB+hU
oIwl5Ar+fOGFToB5zTAK6dnaNgU3zbdJsytKabdVgN8j9xCAcuixz7v3HPwD3Zb5GA7d85+cLM8A
1uLYKoQVmFxU/JRNDE/jAjpqhx6bCZqE8Pho2e3+1o0r2Iu84AAF5s+0/EcHlUrF/fXuu6cjjI2B
M/MDVuW+WP/N67o71hsQKylPkLDzuhwN+Mq9EiVNHItoTfzsnpuUyAROijZAKfv86CXj0sa+9fyB
5BWbJL8qmHxkbuC8+IeBH89RZKN0KU4aKUfOFiVORnfrswNOv5YtEBPB7wKI2C92QPF8OK6tGKkc
OhW/ys0NhKoz3VwVtrVlZwYyjWtyeyhyjipzsL7MeiJsxFdl7t6LhglGQAS2PGJTIMSwrkqhT/SX
oHEIeB8+FcRpexen7o0jPEw2MBFyCllb5fcp6cm7/P+coWLEHemguSuRZJijaR7FB10GAcccWtZP
FMBn+kBae5WdG90iRQF1Up3EfuBZkrNAyliedgAAYzuRwSbzlebHYtrdRP2Cij0lYT6V4vg0mLox
QM4gQpSfmUsRq4HhcUoTYIoipcn/DmXsbudFj9JIFxngGCt/T8YiVwDja4+p7H3Uksj7UTWHeF6q
ItjADhsBy/jHor97TjeYLhetfWv1sPc4OD4glgkz7mqmX2ULaJrf3zVcv0NmRiYw0nPtDdAuFS90
2Ypi8E5D8dDr0jsPBh/H2LzkqRkLkruBpUuIPfZ51I2c5ggZ00C5wkyPbS380ys9ClnoYq/KR/2W
BGVYzeaf26WTl5E6iNL96XQN4+Rk/5Idln8eBK5uAGhTm8Ien+UKJnrvtE+VJKx8jS+94aHUfwSh
20xYb8Mn+gJRkJcyyJaiUO43YKng7O45aZ0g+7QHOXMbONvdJoU2zUm6bsstVARE2kz3B41VbdJ8
NYeL6BsLtOokItXtOVxZy7oDH3Xjbf72Wc9VPPMqq031EQsiFSmVNrkDG1zGq2u+rxnD0bePH90o
1jOHmiFNFJAdW55W4a8/02d4gNRu8MhskJyyxw41luRwN0yqn0DTO536LOQ8tVK3f7DvDFnHubgC
oNagUua9luJ1OHVchu2RLTlH1QfAvnq/00ueXZ4wO8M20jw3BePXcSVU/56sASe4P7H+t8ylBSeN
p3Zos3PkrIrZkDQfUdsX9u/nO+ElXi6pykd9fkDKHY2p2l3pPshRx719dd67ocpcuHiK19sdnUJB
ixl9IAoHHah7hS4usK2nOlITs+P+6nobNNJk7ceNLrTm9/7iZZaQ6mi9wcxIYJitg+1YLEdD1rQb
v4yTGWREx69MOvkoAccNcwS/IY9BQRpk67QJP41Yvty83E5ACghhXX1BkSGHlrYVwuookz0Bozsp
o6lHdFEZNbpZpnxHh0zfIrZl9Ywbq+CSAah9kWRGMHQCxRit4lsSw3y3LnN07q3xPc88AWeuf+pl
Xr55r8qbEw3cwZfXY+erjAspBoVajzs0vQMGEoSuvIV20ts/l7QUnSwgl9yHkBkU2rC9Qa5p0K5m
JOEcAHBTJS+g2rn2C1yYieryZ6E+/zgPkxoDyajwxUMKsVXHgWKAjqSdAY+evhaGCbJ0JYYLYot/
HHU2oPv92vj+OKYG+UTA8NH6MrkquryI4uO/VNkLvf8ScI7Iz+kWiW96MjpI9ZJD8ZFl2vl7WfzQ
iVpre0TP8PzalnD06kvj5NJ+AbTgigfG9uBWhiLJ2IIY1s7hcqGSzXKr3cEyBaR8dkKd1Syw9vgs
X9UKfbQoRlaY79gtAxHrRBHkvUobFjEGtb64IwUy3ox08AH4hFg5Me1ekxnQzTfpPOYnxqH9RVo1
EPK/7m+jQ+DhhxfgiBfhwkdoJiqLGDmTPurdvB9qSjzaKInEPWrsNfBO0RruLqU2Aa2Ek3EXcAnT
r4ikCIAtFq+zeRxvZ0JqSD7weAweaRpOQ+5lbeCu3gbZwxKsak1JYM2v+dq3/DcRvAAcO0D8elt7
SdVZPB+u/igaB+c29Jr3odyBIeL9wim98q0KTVZDEy74h3WoyvXLnb7L+fGMMF5ylBAHe2xG0DBA
r4kjbgi9ZmtGox2r8qgc7lQe+0i15fiSOcLOV+ffU05iWlTLKnJpYt8/3HGyoGgno+nBdXI80H45
DEq0nAcq4b9JJiUBq0m5Tj7ZItFhYoncScXoR5p1S0lDkk3ZZJiqrvPPLCfmZ2m5S2y6oPcveaVR
p7D89T+dD/W71Xf0MmUhT69Noqp+2JKz/a5LyQTLBuYmlHUDleayPVXztY6KmRkUnJHXtVixOvpD
Ro6OIWEdbcCUb3XIPSFczCIZMccb4DHBYDzdkV8bPTbpjAOQWcZ7fKGv5CzXZd9K/8NWeVq8ZuGF
hpsMaSN1Qm5GWZ1OJ4gHFz3E+VqyjmEfk70ZZCLhXmgxNdO1uKyBKALYD+psRo8BSEJKxaIETZSY
RlVxfDGmDe3HpoN2KWyHIrs67+jAPZFcc5Gt2YatQSparP4DKGirwe+rtDqJl+TnCEg7NpAXbywK
14WkmqrcT0B7EaIelqV8N8BsBp5NaVwvJqWGMWGy2b87tyf5DtZTTNazQCDdXbxMwvUhQ0J8ObDP
wXv8d2uKWcx2hzCsArtGAA2PdcPZk/r22hGjuojk7j2aBQfdnFj7DWIjc+j2IoVaRWwj6waT+V/8
sA2hPkfukOWcPkOew5TDHdD4ymZKFNn7EsUFKKKP1cJL9kcZSqduWkGv8C5WxKm8G/astbmk0gKE
f5+ijeuo3e9iJlVjTz1XFNrNcwVaCtRBEkRl1yblk9ll6mMYFqvXxm1aLPrkJYoUnvjXXqnSI8Ud
w50BHlZzr6XG13QXHnXdwdJK4+SEM1Mx2+m8CF9jDwE1wbYVoObXX2kx/LFre4iAYx1cQrhulrJ6
mnrNXEWiBwE9yEFiTrkQYxJ0BhHR/gtk9zMb7t3V367jrVAgccoyH64xvHfztallOuUJ6AUkUf3N
LRRAU1Q6yYPaZXYt4eCanIFOTOnnhBBfMJXcjcXGbMGKbwUtc1kw5q/Px9Uh3zcSAmkuE2Za0KIT
kFUacDCycZRW5E2XAVH0es1v4yLoGE36QKpVzYDsI9KaiXNIJU6eogJsPUtLn3EDdnM1pu3EFALX
uXRMB+KLwPerWQvCr+AI85APmnbYOVlanJ3LWd++dVtCTcz9CNC5194VM+WHd/br5vPzdScJTOwl
tn7sk9bKW1Ajja+yKVe4HIqgcBF65roUnK9uvXDbveU8y8U/WEZadiFZRDLLaNPgL5NdX2Fn5o+t
ZC7rDG4FMfEwyjhxd1lxrRCfoBBGRiBFEE+gmUeHEvPRPEZ7/dDpiVD2VNT+8tqubgE5D8SGm3Q8
tHjyq7Yc+CUKzEoClz4jUVF82mwTqTKLCIyBpB5U7s1mbZJas68oDHJ3+ZNNIuo0R9INe5/YLIpB
bBzCde0JHqQs2AjEYdEUq3zErH6aqRdbeq/158u+5FikLuin8JWnPMF39ghjrIlWIsOxMwP6rfOz
06Hr+fDGchH8P5baLFZp7ec7PhTvxGkYd2CGCnMF8TvoeisH54Npxjvm3x5Is/zrFvzPpgKk72DK
g1aVocALlOq87D+qBkKA90T4fiyF6BRQJVj/9QaIxCEjIqNEDrXKmsgAudSBzu2UNKqlMhAgBo+V
1mS985s+CfYy9Ng5HtHHexFOy2ULBtpVzZEfUlFdkQS/yCuqORdILhbroDjN3a33NO2c66hiCesY
D6sucdBbu3DMu+1KQOxJWUXO9+ZmGJjJ39KCxwlyeJbO2tXvbFeFTQz4kSTw7Nn2nFrh6e892oy3
ucKnsiqwMFo7VzwPnJhASvm4GmJc+RTqPQo4jTEkEILwKUp/cgvESlmDptkwD7S88lzEsGArsBGy
6JsvAAr0U4pbdTDsaOdVQkK9Ojf1Y01U02AN+2vY+n4Jri+HqoSSbvaToavxcm33zWZKAvTRqsr4
YO+IUxpPLWiEoVexjLqAp8vzrNEkhwfaajpej1Dr012Fkhd9IyCRYo2xBhRqTJl5vK+PltfT9p0n
tF/CD3072ppDkMTlK5SL8dFl8b8F3fLjEEFw58JNNkASNTlq7JS8N/3PwCOIG90DygRmhD1jSCBQ
8JvIcBGFLrR/Q7xIVvh/ZBdIbAkYmVnwBoR8nULpFPAVPV66fJnbq7i9o25rqN0A06ubxTGxFo5O
Lr8FAUQinK4+U2Fofg+8totumTlYZ7uRwyamj1aEw14tl3tGTMIN1UAdFUFxwRO5AGHgJhtWBGeq
/RpYks+Mj87iabceypqaHHs376kUjlQAHXHsf/QEo+plouegLSL/nHOepPAZAOA8NUfwOxYwMszo
75ut6zHPNcGA2ZBcXqj35xljB/xT3pJsruQQqX6EHeVuEcnQmDruZyZ+oAU7IbjAFb+SvZr3CB2p
mgiHG3d4riPjlABX9DAONdzSoIvJS9opDnpP8rFmKniALomE+ZTrUFkPgjx6xhLOzTSKek+gHqNM
tHcEwMb5FTB6W6FMs/4aYsusMCCoWZ5FHwzBm+tYhOzCEPGx+fJM1t799pY7SBX93EnihR+D69qg
H7q52EUjRxlT37C8pyPWDPcopF9iZ4qR5Fc/YIx9oTqiMcrCNAswoQFI6E/EmtusJ0Dn27vkOR6F
tpTNqbecje3lyvhHCy28EA69Ga4L1CgnkUsA0aqqrDzKD3n7xro9/BvK2rpHrFyvbrm7FsArGJK/
b4o9hRL5tIBcOC7oXFY3sdOw10GH3Xksqz4NtH1yla8oeutoI9WvzCEgHcCxZrM7iJuJDrvpog9i
5pjwJz9E316cvuyemRYMIWzvvno0/n5lvCkgsz74JPfY7j8kQpwo72U698yWHhXr3U/lT9yyJmy4
aXj6bDrA9MhYsEf5FLbj6keCO6ACbedWfgfNOluPgOUhbXIH0PYMWKvTNClYm1xMOcdS+u4vbqaj
KBY1DtOzCmnNLY1+cbZHEuIA9Nsovd0j2nk/4N0UzJGJOU/UEm116iHCcw3FvctpzUtDE3tf258/
eeFq+VYGbLmR0DsLw0BLwM52yYoAHMQJX9NMKrGnd6ujStiRCHOiapvzjHnx/8+XTXxLnKPrbxnD
6ZxdLv0Ir3/Qs0GKbRtq20pxwBJCxBU/SCm0l7D1JXzx58LPaOtHcFL+wjFutqlEDPN7t3Qx9yQ/
mhA4fk9dFxQLZ4XRiH0WeH2a77kyuNV1piwDAhsrNp5XrY075YZXaXUJBr9n4u+nlkimGyLUW7jO
zckuwxfbDTu/fKbZz48OFAnAGegG+8ukcSFTnUNroCjdpFQy3mIb/xQG6iPFgnPsdL42I0YY8kK+
mh04Husd7U/asR15V8b0E+72ZSItbEzQqkx+l7PeqRaXOeFnKZ2fb+BESFgUamOopALjiJyVu1g0
+FkRhK7jrPICasaqcowHUkWj9oVGOtuqEJefDfZV/A6lK/V++imLUIdp+usA6RCX//D869G710EL
eydtF9txxr3ccRrFspo/xLtGRPqA2FrQKjj+4+AvzKrbEX7XZUU9fXYjE2qex7vuYcHiFt+n/G1o
48GZd3mGWGkahP6Iy4ugTQ9e5O/e/zNqggKkP2ifUi8cql1ohGcIVJAV1AP6nGFKhs7jf0K7cb1d
JpD/c4RUhnNxtNbqYlJwCrVC0CDdR18guiYL1L7NwfQ6HBbNHa04oBNofBH6wwA1AAbOFX/45/BB
cB063eQPT7MKpQc9oantVopGSeizbOFsUqBPbJlaN/T4hHA6ediDFROoD7swvPxGZYSVNz+fniNp
KB9Aj2DMC0PXC+9sxUvw9Kt+RxQtXznK0x1gf39/ZfZse8DBgteR446JXljMRbWaZCzRe5A9aBhP
dYQZt118JUf0YKiCr4CtErepo/6wdp+EyhIeW/WvH1yVHqSP9JLVQsVXMkQRzslJiMlIrAPNlXIC
byfq8tUTPMhEE9lxFEPQOUEXbYtS/gAlmfzCrNvVI1rRNA+RNZl3n7BATmjhZqtBnCxcziNwID00
e2tiSaEBUuFGwJyTJiDNeEBFeNJL2V6f50Va306KoX73uIGY3mrA/Q6NHynaQ6Fh4vB//nDAwArW
J/i7kaiqLIex7TJd3J0ktv+k/04/m0jRfoQDXk++gqoQ54TItSW8f9L5pkYB8cE3oJMiCWnOZ0rf
a0yylKGOO3U+WI/ZjUWoTo/0IWyiqL9664GQ/xYYjGjaosXfi7CGdhqo1SOvKd9zt0UioH1VhAAz
EBPHhvfdeswezj4P8YLYUU9DtqRVvpt3uLqYg4K1a4H/+rmY/lw59Og4OwBewjAP9QUMA/pQqsuq
Y5aTBLEbqhbIBx0K69KbffztHU5yknsKcUKFCo7gZ+BujV+8hUzx2hDQDLClD89Q1Km1zLZsA8Lt
yrG3Ii+uns7/rSUeXcMrAGQT+cSAdFYDx8mtlm5qD+zKK0k22qNqKy6D8U6h+W8U0GHQ5VMOiaYv
X+axx+ii70j/TyPPtxOPq9+1XBti/WeSK91wzpcewgb2v9U2UibiiIcwqVpuI17aGJSMLi+Z3YAN
Llc5C5po8+0SZKN7/I2KiQG31PRzmW6YKemLfk+XLumnlNxQFGKqnOr981pjXSjmdQD75zolRHGF
IhCjVL89AHAuUov+wr/96zhKYu5y32QvlMmVVS0N2yAo/pAbbOoErAOlLKA7EF+N2IVqncA54BP1
yvC+ak/TuPUhgDXaHarzGFKjgietzoRn/VXX9NjKavhHjunLuM68aP1CEvXa88hYgmrtmzMpbZN4
NA4dMho1Em/mkXbt7hWVG5NL6+AO2kVtJG4EmXMVCA3v/vG9PUYaG5AqoDByQ0KEkqJzJkLOrRD8
7gdqvRp9a9KNOyNhTVQo+THwwdZ+cqBvCtNvGqpPoX9UurhaRfleuLqVRwO/Xp0HVrXlRviq3EMc
FdLklf3FDqJc0z1zIOvKiERvAQSJHKj5y886ljRORXlBG739lyoU8k65Ooed7zco8ZHyYG/WlHP9
nVcGTtU6zBcVBBp8yEQfvgTqtlKaJe9wGe64kC5wT4/KuUAsQxGyJuAzf9PJRzwqP3oUTjMOuCuF
RLOAXHGaLnMQzyYLfrePWyV1aZAE/k1f2d59tbxymqB46tOPaR7N9q3iWx+lW33Q8GoNF8JMk5JI
w4VBAWPNffQiv4zY5TGZQykGzMngtZbnYkPfgVz5H1mMdkM+fgSdMYs0WeUW2GI3EhBSRxLof2m1
Z+DD61ncInt06Kcxs9fUn1eKG+OUqDf2tskoiU0nIb/H8C5VLM69lHiM+3gRKeSpV+tnvW+aGZ/R
vhK6uPHpbNgNU8haI4iQ5Q3t3tKDopp4VzKv/bnBjAhVRTb4bWnVp4Dvxzy1ZuhSe8teeM1xmpao
dSlZKCROVs4XtIh2MbrViprvvf/Y8cjKe67gpJiabNdlmj3U9uM3Z9JOGay5d3rmlPlXYzsdYfq6
KI/+/G23T3lpcgtkS9ZYQzrmDDkFCrDV/Sa883vaojMuS63MEcaJ3pUPqnt0pywH9JnXIc+RaucM
Pl92OXkmseRx1WbRKrCXroV5T79B8V0pvh15HqZCISuKLyGmk6L5YCxqJympIUkAjX0t854UaMcn
BaItH4qWTTigtXlDO2o6mqvJDkA9ekkacKpE2I1nsGoTKTEMAHqWrlVjWTERm0m9juXMXbmukXYA
wTLMrUpR+80mSUBDfMB9U+vSZiwzokOHX1UVbIc5++TwEuz9vVJqc41fyUzjgqBkog3dlsQ8gr7j
CPzDDpGkyW6hGmLgE5EbTPzFph5lV3RuZFa/Qi8QB1EZ9yaQ2OcVh32rWEXSZdFxQe0naD+gOPtp
pQWLRE7r0ZmQMwBPNXIX3dRrB3X/3lSGCvydWGzcxITiHjMXvWfvQU5ZqqqdJRelwprQqgAPtTuv
8W7yXK8usKqZ8Txy0lx0vfYVoSFmDtfioPuoVF27bi4Ir9UhmBEgB2JZSPgfYOCmT6LdcOyHrTxu
oqG/dYjHeNzZ5F/PkcsfFivnH4Xif3I62jyAqMeGdSLJsBhLJmIx06Vkkxsf8MgKFrkbnK4xZYXu
Nl1LTtT0jVac+Z5MU5MaQdmGzS4lAD7uXH9tPUbq7w7cRM6KFgrwgM/BtW5gMKIJmpLTx18s5QVn
bSA4eerU8dCcd9PEFyzIkvFtr4lz3sMdFjNOJnUx1mc/+l03ONnE3YhKEsPo2jky2rrCr3VZ0Kt4
g78SGzUPxwXkOCn215gYrTk8KDvY0ejk/cjNQhqwXxwluo0TCT9JaV2O7DaprqtbiOKhwiYAC1U9
QNOvgHSrzn9asJznTgtAGuuIDxnMpNYXnPwf1p11KrsY2XQVtofdt0s/UPNZdrFTQkkojOacxN63
s2cCGaBZ2PJqjZXFrHrSH5KO67dguU/UNNPup1CyJbwcrbKbDwzIQEkRNKVZyVsBEc6YlcG5BEsu
XJ8zBg5d/HHf741pUCdCfJHDDjZmtqfrEOk3llKeGLEIdxDx0ZA9vMuuZuOS3LMrCm5nxcxxfEKT
tauRYLWvNebDDblwXYYq1dtNjK634wlQQkinc10K2Bi416hq9PmchLokd6mRU7e2LbysdcBLx9df
uObq8k+Xl6pN9bnFmJn/Ip0XiqOK5QLvBHYW/Ql6KYfcj71ckUBCo5nTt48doyHVJiacYYS34zzy
Iq3d4Y0Cp+7l2OmfPKoNwtuq1Tq9hZK4CyP21ngWCzraTVHPa66otKWf6DoFaeuaVsTUJ281z9AO
n3tOCO+WyMwpioAX+aVlJSt6DWI3zNjL5k91PyEvjkUZSlTPlAmcVpONz2oPQydBwo95aKfypB7w
lEY4PEb5qegBRx01S21/ti+w1N8xAxfO7fIFn8aSOFLHOetcrxm4kUxZ/EtFFWnFSQlTZzxIVm1L
QcLyyNQZC0eDwOE3NMUvJkumjMJAqF0J7q8EEPFwbjn52wax20SwwK2zjo3M2Y+HSrhXfwY8ErOZ
C1upWAI8KHLvKtSs/sVuGkyEEnpXYkOVT93zOvMe4ZweY1TTcMVw6/60NqTm8PdArxOQIKrUwFRg
BggkyQS+d1dN99GhK0fvhnCXSkmLYq8805pCazuAcTz7erQ3YsBfEC6r4JC9XI7k7TfrXqVvxgwM
nlVzbKiGyAK7Dseq9d2gCzJA7GkEUcwMVJamxX+agXyordy19CTWkgUuiuohVnABknXYBog5tQA1
t2UpA7qpRNPqzn9VgDx5NDGE7fr79JnQAzkyibkJgi1dAf9En916AwAtKyeij/q7v5wiEpsdSFpR
SdtFgd5R+7bUPJ/AHS37rTE1g9zvz6bhzSY7GL9v1dfegaG31fCKW/OeYYf9mCdVxiCjpSg0/LaH
3y+7Gpkf79nHollbyq69vcvz2fyE1KepYEfCQfHQkVMv8at9M+Poh5CepiCYZWIWNH4eGEYhnUgK
XBQmun1YcP9JjdEdeIVa3jpQtO6S0vhh1tly+laFDRfmp0HmTvN8HF3sa704mhaluRp5BZGrtOZf
axGiWTDQucp5HPbIIlPt9Q4XkNb76UDN/45AAa6v5znz3xvVdOrVQzG/bs6F1OUsqJFLIsNTjqWs
Dk3Ve3dTniMuwqnjN/oxui6IXIAPJeMbscy9YJtG0hAyxkT3ygG9mWJpS5lwH5U6lZDzDVcJ6rq/
DzgYdERKjMrYKFZh4smU/G6UiTP7gxhngNNRVdTWgcEN+M+rE9zsLINmPAq/ziEbh/iI0FLY0J68
di2kBj/9GVojJQN5o1+NLU5y4aMw+maAoAY//gJa5zDIP+G5L38dd09IwxvU48IETixj4yQycEyC
HNKWz5dyTjEAm7WymZXhCu4Eewejmjg27NskIgpVVw7LmhGaYGbs9k9hQP1ZahLYHTuzV0aKpYbg
mm6Mpi9Ccf6IZpfbqrlGOYx93DnvGdNrnaVOHfk14XA2TWr+6m1EnX5Jm4pcMmafLvDF9fQR6+Qf
EUgqD5wMtObvB065noP83LKwv7L/IxQ5qhMqd8IC3rorEMl91V4mv8WdHK+K7seu5oQpbMW6M+7w
ESdOSppQY2EDpkIaQPFlUXdrIGaqHSoNjOJ7vh4ymDytG1+57GVnn94NNdnq0zDNtysFDiN3TzTj
1eqRAGOb+QkhXW6S9rD2ospsJQPIaouczBMRQhD5WJV2Dptpno2jneOpxOOqVBI6HYwXMZNWO8cj
tqMh6oM/95KOnneBK4jw2LsHyyIv2UVR43fPGExHJgqXrqjfF7ODwc2lVQxgY6mIkuECRxOtMrFO
Vo4QMZejxkG58uvEBNVf9o8xGO88JQguOlBUBWvUW/aRiu9c2Snv6J27HSQZ7FurJrHD6hHUzfkN
gmakp1uxC9jNzw463OLCFdbhqlvFKl4nPS/iuik4FFWc4aIinA48tZH4gTdrGsJY8BQJrYhcreID
ApDL+cnaNVOMRC0Zb8rke45t66Mv5GJKEgOsB3IWZro0a/M6wqQrfDF4WginZPjVZ1eeuBg+SbCd
KTGSonkUupfdRZc/H7s7GRiNX0SAKfY+37Y5Vib7ZOog1aRLipVvhOcrkwjWx4wDz1fMMHGshxjr
PKtFNAx80N6+xAbJ36wL3UzyM/Qi6fc6iTqkdPPus3ekTIUds27YGmQt47ZtarKhzlviYcIGiac6
X4MzqvqkPsm7BIPg0XJ9oCr6WVX10ycc0yC91IVXz9O8OZjzjoRkb4lucICri/+QT0cVGfvruxoi
YS0zvRlW8fhKzAWh0jF2AlFv+34a3e5hqLyWYkWYiQWilo2yXNTPy2UqDlfwRv4qBXFm35n0Jv+2
Km9kAceT6EX4eDcenhDyrbjOnHP+kjp9Cwh6JuNNZBAkrvMUV4Db2QN+spXe4LDcdzovabpIP6SM
CZSSoSnUBV7PKo9DWwchNiVxaAh8to97Mccg30iaJvvHdj8RBU7QaGJnqCwo4IFPtTYacI473nIn
kttOPN4CkAAPieC8egevVh3cZLbji4VcHS/DmVD9O1hpDGx20V5jWQHViUApRK2+In3gMrerw6uB
rglrAO9JE82MNtJPC8xXVcI2XoKQNsxyeaUlhXUV/kIT1hDUnJqpDTXGupNHtmcVQ/ygcogmskdY
8WLPdYbgnRFKt3EV5cuf0Lnl2yizgh/XJ+/2hxJMYRmZh60iKghnQcA0XmspdscjdQ3OEIwrZA8g
Ebh0/GgELSLZPun/EEiL7u3j42qZUoLY9lsqAVJ2bhczfY6bxRW8U0r/9/vFkOVaobI15eSwsaDS
rVvMLqR3rFNrP64KVvyZRH13p7KIKGd3fWS+VNXOBtM4uEIHu+OEmJQ10cDxgvpBBUzf2GsnYdb4
L6NFiS7jJLpue1+KbdPr734fD8fy4gjlSZO0N9nVIV7hlrIGB8BcPKPK68GgaAfbsGqY4Rhxzy+4
dWmbUVelvsiZzmqOz8GgI70PmpZ2RV+ejScqE3Rv22Pliq8htWpRKr7whBX2lO+CT1bCWqys/T3M
5KQIuKbkue7HRHQ3Zw7qqstHXbRvU//jEsT3iR1z/3Jjkyh+Grprg5XRErGwiUsARs8FdIxBrL15
Y3GElM5WyMS34mTJbG/GfJGv0Mk9qYwNGn1N1q/4rsqNPxBQ5TTB9ZXSvZVEDEaT7Uhln+I1GEqx
oUwmiI9I4O3+4YTnkA9gQZCXhJwWX4JFN9KUYEYLFWQ9qII1eD+Ckt8o+Zm9xbi2jN5fO+C9EvR8
73kMqskWFpFtipq1QhkjPTLXWfcgb+YbmwaEFuZj0o1sykOn7QKVsMzty7dgOT4EVsr3rKoAhapc
Pi2hp/Jzzr5DNKAexd/cFlHZ/NQrNW2EfyJKj6IMnaAMXTOBWM8hVfeVB+Ij6rICv2d+b/KtrFNf
L1bj6ofRp2h55XhXqSws9xy0sjBxkWV9q+sERaNPQPGG8ndS0zOI0vbItzPHvJ76HE/jxVJF1BSJ
JPAN18T72SIL2wwJevQq6VGea9mbylUgXBzRrnckrKUWP9517mdhsmwWl7VT1fDIcnobyztUfW3o
yWNlnSmKWgPlBs9ajM072GXyujQhsAAkAL7R9UDFWKYKxl2SqLi8BTX1zlgRgDERWVrODq1awQYW
gwcuSyXOp3O8krlCVwAPkNGZOPeTpenDxFhvuuOQ3U865QewccWbHV9Z+9ndXpHlwb53jpiaEuD7
yYaIxPCQrXCuOfpzONi8D/Tx03Y/KbsLv77uAQXczNF6+9Q0RXbd+jctGwdW/gcyNBvKmPw2Ui9m
Iqkw8mXDgIWflzJoa/THPpc77x6maCPh3CzUdECRPlA8bF1rerIBIhO6rMArisRjAKRER1qZ/aWv
fkcI2ygPPec5OJwWZWumt8sdmqgV54SnWeRTPk6y7ncNJ4pwIru9n12AcGZ0t+OARlzlkXicoUJg
IXsqrW3SZNx4P6zM49qDuCh11ogVVX1hc5r+prLIcaf0ds+9Egf0HiKD2voe/058wjFky6w7dU1L
0Nuv1shah3kcp2pU2SxWDUq2Zv5enwTTG88i5w4QbcGLWgVNGe740Y9ZjoVZHz7Zj98xCaqZCecn
yPbP59IFOLdBs+nydV+YgIjaLS0gUnjeUIMZZPlggBgTnekbQbeO0gzCZH9Q2l+s4S+DPF9N7TyU
TFJhUWMqZ6gS1CfnekOYEZ9rrvz+SieCsheCYduAIsIeOxEKRf7pCYKllveqwyqGeI3FD7/6qPo9
sMGR+DY1bokc7rjOWy4puQJ5NUCxmTKuRpbGy1Eopb1fOrWoS7lC+mVQX3A0LPI3b27F2ZaeUakQ
d7lQZuboZJnojpNIFWW9toTxctJPpCFkykHIGB4YpKkkK359R5h0ZC3HpUig2asg7LO0LmkWG+5H
ijPHLiKv8cQlB1alLi89VWJ4tZS7BS+mWhwIKnsCpz89jGwPJwNbX1UjonGAdgribaPCx+BhiF26
sM4kfeoVSFd/pjxoxXX16VF++nLtHzdVgBkJ61BBnsmypLaOe5FVwBsRGWMU5nhMnWzvveoUe85i
3BhMujWHjdU0ULYX5mU/lxsmCZpc2sE2TaWj5B8gQMqv7WwhGrytGKpU48BvpXGtGQn1U/QBc9Ph
7QjQiIcny+F9Qaqy0nmHQ30u3CjYDZTPLyA/35QMVw7/jLQ4D+v3exVA5R3gzMsQ4KsrN5qEEf0h
gGseLz1ZTj7ogpl8LQJS1Q+F9AZnDWZ1TtQDFyi2jpDd3/F2qyJfR6iGLGa8BSi0w04sqZo6UVI6
h2Xk0Ao0FMsx6fVkaOjy7bMrMOSdKVBIE2SZ6oVGBopXDuX0IAUkdArJep5BrUXxtIKkBcFApNx7
K7WWxLSZiGXj6mow4DGaghd+CRRf3c/70SS5UxNbQpDvdeyKKiYlfmy/nLCMSNvvFEN0NLwdjOYd
BO1c4fPTDq9WWOySfrLetlv3WjSFnr4LkT1gqi5h5OaXiEf4euFns9n+5+7H9+aLtrbiVYj6a0Cg
s7lm9J/ywafmjIFGYQHt2S4YuCeIdD17tdq7ofBYyoSXcJCeP1b5UV/AIC377pEdgQOb2b6uklU/
/pfweBBlNZMi9NtSBp5sHCwtVTIyKiijmqYNFZ6Z6SDKeLrB7qTzk2+aL0gi9b0U5JQwjgNSM5Q5
hbwupT1ueXjQfzVI2KlaLEdQUjyZziTuSSoTAoV34IS7TMgFIMZlCeuNfYKlOv0N7yd08Z6PDd2b
yDR45+XWMrPyMyJHUA9R1C6/9idsRl0Xv3xxIqpq/jJTIAnaZTEKsRlD44FrXqHSOeKEaUJujguu
Fpc+OY4PkiHqdLg5AF1EAlCblTDbYfHkt+wDjHn1PSfVzjZEQCLnk4HfdcukocGhvtKA0hHcFtiP
8n7yMOwEUi3v2z3vCraH2tmToDE5VOUeX3osYvg+S86LjF0aQbDYh36ZHLk/UxNSPAc8eelf+nnq
d7yxB94UGUJftSTB7h4Z9NmCRG6d9g+5htiX2nPdPvhKYF1zUeej6RZwBJKk0j7RvaH6ab21W2ys
QU/FLwXtOA52kMzNIJW0YKK/f+fnh6bvvt4brNK8C2EBI0fZH3KTSOSyvFN75hnAn/Rktnp7PA+x
lF4UI+MgXoL4ceJuzY7hmBuHRp2VUfxFXWHYjyQZcV0TPn8dtk4XpNbswio0UJfneP2TaF6Y/S96
cs+ZlS3wdjuyyXu1LdQNYaukvU1a+SD2cQ73ZwZr6GGfwnbD56gBeROT+CDkDQRlWLAvvzEez6lK
NMXNWeCXD28Nr5O7oUhWNtPqY7B0iBTCrx8mZ1grsj7AgB3zPuQSzXp7ERz+NkwDgedzR1wqmAOC
8Q0yZJ4HS6W2clwSoLI+rzvYpcHDUdFYvl6dFwq54iW0Ad9JeJEuj9KzzZDXnJQF6V9g7Xl62aOW
fDagbeGzk5Fox2qFwCjsX2NKvFMqtc3DEfg4mheex9GXSblMuvc9f9MO/KJHlAOBui8yGvdBMs4D
bXdKNw2+IrlTgjvBKwOvP5xGsiTxWT5itOhfKUGFhKy1UXglrjHOYD62dlyro3R9wGMxrHN45mAE
wjG+9SR01NRCKwxfF2Vy9JTa6ueJtvrf/RTegc6xlsuQ/cEFg6tO133yOzW+lYkp9ayNRaYKkD35
q23BgxTCnABv4nyj3iyTes3KaU2jT0luysT//KQeqXj/CYkTbiuqrE5e31FduoNk2OBDG08utk0R
nigbhp79ePz6r03yYnNp8ZaXSZvawCza1cT7Vuz8OeMUaM17wsuc1U/Drw5OVp+KVH10oAIWYW06
ikhad5yq34peeQDS1MHqETiduYB2+ndHPAcoIrCTjipq7wQ+fuYATE0VtjKwtPGalLnzXeuYFFq0
AcSOMc8v7J50PdIeWtOdMCIsGvwqjf0kOPn7UvtOrD3xarbb3UgcCxhbKlse7srYekV0Anv8xAzU
IyLvsYSc7IwyRD6l9eIOyYE9XHZIcX63Mr4ePdu9XKkITvEFloP+0LOkS7lAEmAKrsoIttAofU0F
vxFFASCW+UVxUq/8XvJNepAXv2z/2Y5UtOmoorPhM6Z7Aa1KaFWK16q2k9l3JI/XHidZswzzvyQk
6RQMSKprHF+QWKIZzifpGKLjoFW4rnHWcb/8n9z4Txj61rPsWuTVFp+JXwr/3kQvV9+5GjicR6d6
zHIk4p+PZw5AzY8FTXm2TmOVlNcLB7cj0uCHcpj7vd0VVgENL+bOU2yGLmiHEkX4MvtiUbVMImAA
HfADkBR3pEj0ORst3C/SLHHEhSlRvHwYZ22EQPygjRmprxnk7Enl4HhiiyDyLCd1iw8csD+4GkwV
3tsuFXJJn7XaYGpSLFe1ro/8ayP+JEINPNZ0c/9D7oA3SEglB5Ed7nny9upY4osWOuLAca5aaGzJ
YgABAotK5+vzs8Gqp+/FYeXnTqRAvr1ExTF7+UuV0SjkB5hlwQ7rqvztaTZMV28ybvyZWVjHIkqS
MGE0mtAvYQKWtcKT7v8DG7y8zlvrdcz7VtR40fI49cLON1QqcReRbaiU7PatZD5tthfBRqDagg0f
ClqbgJxvHYmZ4S6eygocjiJoTSZZEkCsxI6YGwVxpYVPoBO3L0VncwATTRIfK8Q4fziKEaD1XiTi
Uw/H/M3Z4zKOge0G5ZISqWFJ+gFkWOmrsZ12MBy/HRmfi6kLZcCipWEssirXX2pr48fi2LITGjv1
QnRwTJ8osM2Nf/HNXPvD7AbThQuL5bSdHS89HMU/g8GzHgZheHXPtLr7tlQUF3t3xS4nXa6q/FIF
1kmhOEGzUtiQJIx0JhSDBQKMxK0gJhT2tfOqUapsN7z8GlQzz81M1DPsni9Mh7g7bqeKBJhAMNIy
qiyaWpRPH4mmwtrtgiz7iBYk1c2aKR8kYdBdtR08OwWUiMZETrE3qLnulattTNNxgNQz76f4uisV
+DSQ/BuhLEMFERbt8tgqM7cROhZ+stHIdz0EumDCZDYloNt/xD//NG5z3sV3+UXp0G5ssY+njk5+
LjljNv5rud2HvdeiOC8rxPFmQ/e/zPRa8PE+oQxCrjIw1Q0FNG6hLTPN1tVdw/EvwcL034fhwoN/
O7bI0adVC+0Ug+caWnIreDSMPY+ZfvDOmVZlgwmtz7ccWfHhvHyWN6DpbFX6Uh1v+gWzMgVDsiLj
j+8wd+upgvICfyGz2n3dcFd1kJ0VV2w7iPpT5z1fMKtYqzxoUE4bEvFzvqOsk/4gSwXDN6WS3xr+
O+fnKccEhnqzPEyvfW589rlJfzHwU0EdqMyXR5eqRzahLTf49yJBBi+imwyuSDI+y0VxZsMPNY8S
v+We6H5+LiRe54cDBqZpOwYc6vlIJrErRK69O3SV5zDjhFBiMw1BeC9UYFE+yZp+hIqtB7C2KTfJ
HZSmKbJM8Ns27uq8FnCF4UGXOL+Jn4FVI7Cx07mXxIeKHmYZtc1mFsS44Y1DY04bnATqYJfq2zk+
xrs1V9/F6JeLho4Y5Z40RYTBFHbIn73YJFrxzjYjIHbAkonXFlCeRvsW3tJ8rvq+Z2nOzmEcoVXh
if5mPSMNl1SpHOHsyEw9OoIa8NBxPlaDiYrTAd3TP8mFqMRfBc3Jp8KihFmUqNBgNsJMYbvSFlWy
j/0rG7yiULzUv+cHQsdOdJTMEjmyePeTyrg7NO4HZhp+J8q4F0da8pF+baGYDGM9jO+uYth8gEqC
okk/2+S7gPtqwlM6zjfmIBkkD9m7LCQ1mU34IzKMJOdrMrwEqUP/L+r6tklVbLRRVkiHhGd/iw9t
X/RjvuC+gY09THT1/34zMASF84PessFvR3yRmXLEO+HC1AopmYGHTYcY9OuWKatxDGW94kq/Zn+R
7aJlTsTZvGcT66VB/TXTpKg17SuH8Q+zKeYuvLgDyTG7buk7kf/rn1w2YklNjUB6oMKgmwY540Z4
yS3PU1ZedQEEeQ7rOrYwqFHcATODJAtDM+CUkQwKBzKEik0+FdFOffuR0VNpQfSGKXzekcqMulwg
zs/uWGhxMZYU4dQBB87nYWXNW0XgIa89Hvt0QyoULDdR12A3yTa42F1xeXbOAq27cdFoklNhXUDn
tSq7GUYHKtLE73Az/5L5tIOZe8sVHd+bxMUqiXfemlDN4zLs0hY07wB/d67xZ8w90V4cM90KdIKE
ZbuZPGDHNkZMmx+qGoTathONkgTn+/5rUNYLeXrt3Toz8Spm3sYUtUSMnXXqOdSMpuArFy1bjJYY
zR1F97byIGRX1GSpCWNG375BpOs3ZaZ4Fq1bYKiesyqnC1wu2zAp409jgzmOcHCJ1GTOxw8bq40h
mRCUSXAVNqwYlnZDXKBbDJ2R3sfUZOkaGdcwuWXw/2X6cUXEidav/Icz7d3MXk8JaciClLBRviRd
8MXQhBtu9DAkMCAoF7JwHgpkGDAfbb+eR4IANH5jZfqkzCz133/Qn0glC+jz6U9paj23F35OPyIR
gpnW2J7FgTb9gkUAUyRGr1AUpMSpbIygdxIOzmkuDKDJNVNe3uUJ+ojABS8LvJEXvb2h4WhMfWP0
DrRNURiqoLdYiigk5n4pl3xstsumU4eB7f2i71njuewfj2z59K6arF0gYJ+GA2SLWNSAwpRJAktd
+/VEtDoBGmVN7EBiUqo2HlDucUA2raCe1F0RpxvSMS93ru0VWJBeWBb/qRaLzVoMi7ZHnuZqHwxG
njhzMVEiM96LCDE3g3X4RB+vpwvCrlKKp+6LNmsEiViHokLceGZq5PEdhusey+gJTurSEJCNeEYK
bOn5FOjtIMqBgXT+uRFgW0XwvHniYtHFfIPsj/Nm9IuaRf+ZShjKMhI+ezzyJIaQsdiVSwQsjcIu
1YTiRDWQzYY6ip2n6cTZ8uxepw22UiepuRrgP9RzIkPxI2kP9kYTP1r8A8Ng0ttu83myWmFV85Ls
/vfY19jxuH/eEMbSXA3tvFydo00ODeFrq7ABqREAl6HLI+AaUe2MCJewXeq14eAaqFKtZ6ttsDwy
w8NXmbcqHDFG3xWu1np4YFij9+fDEBkHEKIy0bgM2Hrjyl4kwlz93GRgH6dWSeUPQjyzwKBlre3L
d/bWs+1HL0hoxDPO1TuDhl5AdjQDzwWhCjD+ETXsEi47akI5ZKQbfRjLktCJf3EeJBmuEUAVcG8y
5rkcPsKQm8ogEqFSBb/kCZzfI9LE571/c8UbCrjDDWi+dTQVE4d8bdQJalOYlSnvsjZDs0oVXjqd
MdrH3YFUa3oB/uZj/OvhNj0wWw3uEG3b5iN6SByxo+ettHSzlrcYcd8lMlMFyy/NYOctiVp9AG48
w/XYFJrrFmfq7VnDZIcLRcp7pXCx0oi4161nQVMIKosDGT6HKLvj0l3yo+9WGtHiWQ3vDfxJlESp
qsZrlb43HeSL/XMqu1KZ1BSJVEDGQVu+IdkpGWo71kRsJ/WXSBfvRw6u+lARgP/XLDjp2HgfVtlY
XHrhmkqygbOUXXqeV/BJ2Y1Gvjf/MP1XPjAXzKrOpWAGKChkDkThNgtnSQ/ZmJKmQkYGvURQTFDi
2FjER/RwldHRWuTPe4oMSBEDGJ+7NVwymn6eqDljT0t0qCg7ywHA5FeEOAXTm2oChXp7elBTSrYU
X90hTei7eFJM/IoGxhCiH7PcK9hlc+FKEQYkBEqvH+cagrbI2jmjnbPegUgkjHA5jsMVvEjCAARy
ISE71RVHOxN+T7IoIZDIHS4nlGsB6HzGU6Aab+14+iWV7ENXjO/ExiG478tz85JpelXRPGx6Cxxn
qOkP+1RYK8yyykB03jsUcEyQ1gGcO4+zl4kP35UpY++k3RmMmWxp2ilofSX3IYOtrjJ75Ra8buK5
2NBIeLXBT7Nb38lmMSFN5EG5NhY2WxtwmQctrcd9ZxlYPY0LdO7MEofB8ICb++z8lMjuCEKW2vhe
EgvPGAyKjYwwsGiEz1fu1WudJPG0/9HYtdLvjO+T7QB5KOt6sl17QUAA62LK0DVAwH6/qrbQqTZZ
ferNkOJ7XYIvsFiQnhHY1XOZlp+4cKWv0rFpY/9uji1paI8fCsSL2Dcu1oXk0XjSgOHoFlttphBC
UUUBahnXbvSag+QFy0sIKgO/dUzHV8yI1nFDWox6Ortmx2G5Jdq/iFBZKOU6GxapBntSToZWWN8k
CFGvR00TEJF62It61q89Qb3bdp8KimY4UbSRG1Qzo5O/fv0AXb1LlbcQPWpXcLsDHpmnt8PY3+Rg
OFU2DTK5cj4EA7zWQLS1Z72a9CYVdedc26kQcTocSkM4zyRUlqYv/KqPHdDVNnTdpMyahH0SH1GA
zvYNNSDmx2TkfFRMIc+nhcEQhvS7sDHsUwdzig/ZJpnPcw0Qqz/lY5g7fLnpJ5ji9AnDebAOUl8s
RYAiFlN0avXtrytzvNHWLNeRksbCLG7VyFgDXHbjTHDEMGf1B8bwa9ZhXYxAxI+ctXa+jvSskvOl
aZHtkt92XcW7g1jQllnneaZt2F+76IzQW+dY5G/OdHZr85tzUWcjPfYqWA20OzVgnOVqfgV5jEQG
cvruubmfQrIXmxmgim48/3lmgw8YEQY093etsvMPE3Je6FBBqYfbN95j7I17nS6FkFLmZvG8D6fg
inKPmFiNfH3ekw4aNb52yLv+oUNNs5EFBTW5Y9Fx5Tubu1V7DMlw3sz2joEG9DuzyYjC77ufVsfe
mVu34Ax/S6/oa1Ps6GKE49r4i5V5feQDPvu/LcYxLHpfklX7D6JPPf2tJ1f5db4zGp3vVXT8Ye4z
4jerPahgNzYTbbQNZZYaURzdvTS97udX1MdzjiQQvmIogRu1Y8330XrK6x6ulwMNhstn9dqWgaEq
QqVS2OFo3cAiDq5K7PrKkX468RklyxRtajSu9oxp0tr00m8Dr1FK3ZW6DJCmCrF+RH1Y/3l+wNJm
VXodud26gHeWsuC8hfk/brQlKJtYJVYBUuq92uWiqn/ia4Su5dZVW5X3JghugDxTpk15banzGWmu
+ic5MUEGEBm5PLDs37SiHpVTvQMCOn8yofzoEX6nWJ04zfyQW83j+0RvtOyQFym8Xe1/eZIfDcAn
I15iuP2Dhm1bW+/zbhNwx4/4xC6+hnam5npMQOhO+gMg7h3PUCuC1cHvx0V+NiwCMDBia2Ta522f
Uny75nHoblX8Z0lGuwHR4ZgVF4OJJELNNnoj2NBbzm5Q4JcOCLPe7hHMj+i1wjwprrFGhrbx9OyF
5us4P9Dgadx5FRBLuo4OWBPqMilmZW9yv+UDQF+NwL9FFGWu4Nfc7v6NH8wqCrMWAhGmQrwGi5aM
emFgR+/8bNTpXdxJ50bSN5oSuNyuERgBEPMKLfarC6WUrBty6BgiL3E7iqhTQUKyzyuvqi2tVe6l
aSkzTiHAfQ8Z/uywGqS+/U+m+HFyscoAC1M8K//Hic4g+hNP1ywJ/Eu7u+hf1tmIew4Ctb59xpda
Z2BVZkgUaYQ8WTm0JSxCAL3HhWJ4qSlLKrMKXL9tKYxXoFGnW0XX6fSzCKG7q45ui+IZgkmKfGT4
R7sVbHjFTIqmaDRYilV5/0+jL5FJ3AI5PtNlOA53CYUmHjsJK4vghXwWoM8X21PBrjXwsU8FzywF
5O9GCxSxvvmjOFq/1Tz9tfhOayQb6pUIk/93HS/ipNnfmNRTDlgX5UKfqMT4EAoxw+QFHXVoHO9+
0nkQ8FP02aauusDoeC/bxBnqkjTVYWUjqnAhY/F954yz9c6OK1jESAXA9ZwoKF5+1IVZammIj7uT
djzqYtuzXzD0I5scw6LlEYVaTthIRUPFY84uhiyaNX7Qp/beZo/7tVZD23lNEMIZime5y46+OALM
Yi2KHc7+YdLgdn1nYTyhaIVz7/htaSIm4I+HNKYsWsHVO80T9cqmHmQlhsPjkCtabB75xJFpenRO
ioNzuGOebWzh6Kn9WhMnjVxlUP+SDtyBIfeKdCUAvSHmQobqSqDi3ezfJ8ygJUjnn8UN1Lnd0x+/
qM7jSvvdMLoWIgPVysMknPAENqWCksszLFZzbedjBm05YzeUCe/M+MKrnkEE0eeLBxYc064iv4pW
ucgfbddmdDjYxl35mywPd7ia+tgqcodnk6bTg66QMsFgrfoZVHcbROTtqG1B5k141LFvXjCZN2vH
G545DZX5Wo7zQAmxaPK6nNbSLm0XTu/8u3ZnJ/ZUdbcIjGwTp97FzgS1PaWAASj3UFfFFOetS0Uo
DSAZTNV+c12gZXDnI9talNjzmJne5ReQq4pIkVrFCeIUJ/JabwC1L1wNzDN7gIyJuoIu1HrqVJXT
KfuuJ2uS8s6trBQf9ZjblLq+c8MScmTJ/BxYbdZvkkK6Kv+w+71592Y7Nl1I19XbByrtiWNv1tL9
WhxkftucdvB0x7AMD/D52qOadUSYr+B+PCqZBfGQf5LII5v1NwteO6LS4nT3nVf207FjTmZqjqSB
NRsRCBBf3+UqSF0JZyQqYKWvxLMVgN9oS7+cb8kq73NGvfBSd0V9IUSz+weLrxRZxRismHG3+9mb
OqJfdur26sbdFot3YfY+akvCABzXCR9WDifoWzorXu4pcbH3R0yrYTd1mMozMSIIxNveiWzN9qWR
rQwZjSVDYvMF7bYGlWfYKBZbezrVbZ8ElYIn2c+oZmnVtadtPx2W/sW/an5oUitvFj0Y2BfaCapR
+tcoZLF30kyI2o1ovcpP73/FUcrKpN7ByaQjLQzjzzxBQDp1xo6Pxcfa+8gL+/uMwPbG2+gKQsLL
AYiJnoG9KXnE+N9Gdw9+rU+PjtRaW0dPlCmmPCt001KlFCkSUGQiO6rHQZ4Q3DvgxZ1fhI4TEqlW
wA8M58uqeBrid0DJ9OZarndCB6O4P0tHqwZ9uX+b9OvCYQCFpBG/Y35skN0eHfVqSk6etSBRquDp
9hBvK/JwhOitXuTBo1Vj6OMgPc/ySvpVqMpQYHU+r9JRQyotvu4M+acaQipV28QvFKUwKJ6PgNpp
1QAr7536SbTqd4iysPrw6BplbGrBgJpnU2641cVYBNsHg3T/N9AOJmu6G/oFeYDBDANXPkha8PWq
hOXzHZWreoeE9ZUaZOR7Nr3iRozzCSirO8t8J8Lnpvtec+nEY1SkLCQlBLAd+lBTeheDevqZhCIs
8xg4Otb5FEs5MLeqoGpTD4kwNclV9cz346Eq6U7pTDGeSApyLJymrsmerwIK0FHegz0fZciAM00Q
GOBeVPZyxbWzj2OzChts7ww27GB7BuC1cyy81pI+5du9C5EMyM79qgOFwXry3cPnN+3tO3M9CSrq
Pz3WGYMsonX8VILWK8XXGIbaXdSYALyESm0CiStYxKHAi7x13DoQRIJJ869Dj17NeDMWdx8HAPQ7
T68GGRH/hL16jHuwCAfVl9y3qve8rcsp4cxsx1sea3AKHty2aU7QGabE4ndWen4D7WWrov3xAX5c
SHV9cEWZ9nw87LA++bIWm1a7wXatzRwc6aD0seJSfFQaSb4fxLa3q+dMyrvC5ocI+b+ItVPv1BYK
ev93AxJbYr3vcUot+T+OaEHyOFFk+dJsE8IgtCXc61/QXgm42WGCejd1oHKicH+5b5IJQT/d9fZT
PYxnsDIAkOqd7ZKSNpPJ80W0C+77bKB/8ZnMNpjMWrz+9h4mnCNtjXmJRu8lxyCUtF7N3XD7aq9P
KU/o2ujFfOCo7iTH2tHByQnM9K5LRGUPVIJUDe37OktS5KMOejsVITfDi0mq15BlEMPJnsZrFHei
pxU2zYdbFA3T1b/NLCfXbG6Ok73KsXmfmXLOWbtI0TXNbbZaw2YbGxC4D9LA3j/8I1oyxp9RVNpC
mfj+YLC7PasWDYazT7oLHy8LhUStotwK/80mE8KmUK79q+ZV20/DIQ3RjcjpsYZRlL1+rhPA1+Fd
FfzYAV76aEnKLEhcOCIkKeeoBEu45W0O5M9dSA+5VgErfY7e4xatHpEfZ4YQPv5MQaW+jYcgsCUi
I5ephzep4ZGBPQe9aUKgSddmxyaQUA0tMY3Q5MpBqL+VVEPkvba5CXhTjqMel+eviMWs0g/s2c82
P1KSs3Dp7de2tQD/gfe+K6Tlc3fdv7bnpQJXbjBMiXw9PUMeLYrm0dxzI+O0ylEKahItuQ2h5yRY
YnngnGXYRTzFAdhuzCgV/+ntFBY98ea4sejgxOqaMQSrIype3uoAbFEnRUfouL3ao5Gea4Z704ay
0Ol4mOzYxEBOmBhu7NHyZ8tu6nNfpLV9RIFqo+6PbU3m7bhfpcGoAC2rdedJB1YWJ3W9/9aG1UhX
ytMKPP5y19Vhgkql3R+QYGz3yTwJnHt14qviTCPoYGRE1wRifrHJF1Se58cu4OXtI3B8FHANim/M
UbZS2rAOUtNKn0iZlO8N99g+BMK+kM1zj2bvXrti/d4BirLRgwTTzZkCCRCwWKokoUYLIOwKJMzm
p4ya91+d2jN8yjkbWo1Ukd7UkdrG5M5/pT5VWXfi+hoFXnZ7s3z47nQqCzOkZFk/wN4YAX70Ib67
uWCISghIRAF3jXQk3V3MSA9abxB1GshTPbELKaSMm0Bv1nyAA2FAIb5gCAftKFz25cpJIexnX1yi
CZewIHuQ0zA/YS1/yZ71k3aBD5+jDoJgjSK2ah6UnAyPre3dWHdS476M7r8RmOif1WojQMWONUGP
ZWKYKIHIDzCuq8j/wgqveNJEsxZWXcexChjY0RiCGDERiCaaGIsYc5xq5iq8YodHj6k5al0lJyCz
VskkMOubLjydTmBd09PL2rHT58RYpJUUijYjEZyKHAOaWfThJlzfedB4ZjydaxaTUzJPBvNQ6iSu
+87k7le0KHcEutz1TPpk9457J7o0YwJb8Y0agKqg7FY0gsy/XKh/7BDIK34XXmrQvUHUsx4ispbA
mwvT1XQoeF+Xwb+lS1renkuXpYXmhkTHvOBzXaWps1lVogu0deMRPsBTORTDIILUqUrJiTwI0Gim
HXOftBFKklbdDneqByMAU2n/pgkcDY+Vz1KCQpIYJPqRWDW6texLt2rrRRDqK+bSkFosk6oGaDbk
j9X3gEVlhzbmFv1ff70XmgSPIyvziV3sF8Rax9DnLo8LJKL/1dcYwKJLCxQp+NpQgxBBkzfm0DcW
/AMk7HCfMhdDQeGVR6sVfHo11ZPyBA00lvJnAKn/i79xckPlXSpN4jocwn4xIag0+wsE0ZJHNpoN
3GN1a1RwOI8rbRrh5mjoZYwPEGmRPLH/bHxY7aNsBtICHbK+wzaCgLHAtdHenOgdo66JaFlgmsWK
6W4oxqiec5w2HivSqfE7jlNSdV43w9z2lioW7yGVos5N1L0Reek82ilRWEdtHWA1NU7Z29Wt1OGu
ACFWhnytXR2FsbFiao86LQJAlBNZd4wI0+iVPTE7u9lPc9hEWu4+Wp6+k4ffUBFODEUlbR34QO6n
EPCqYTAwo7P2Euz4aewpTWh5X4q2apgrsxjsn5OtBKKAk+jexUiuviU39nqnUtqdRMLMv8S5RYfs
b4Uds825OM1qJXtrcR+A6BFmwt30rQ5IOXhGHD/jHCsEHu1JixWmvvSYir4+eZO08E++Offa6euP
lyKrp1g0lxRYBDTDDO4DbGVWPXhlS27Srh5mw5DtmiBJD0xTFefDZxE2FzLxHk9n+3pAtMq/khCe
lVxEkc+DbAiWUmptnvL8zSo7GLfOqEK+5niDMqzMLFQ8LiGMkj2c4JRpyHzXHzsntKUxHqVtGPEL
+hjwMqmsXTa3vLdcfUhFNtwKGBWjBKeJVdQcZBXQLa/aShMPWdjfqA233VOiApqsR+KUOZIg+AOB
0wiCrNkuA0VYOC89wZZrxZKxk/GvjNPX8SKUblAz3dU9TFlcCMfmvkOvNyz1KgKLpKoO+Prq2sik
dxxwxgJxrWaxR0kobz673SGAnZWPhzhchB5DUGJwyeEdqxnnRn4SX6DdosfGv1zpWtXbXmeE69DS
poSI1nSYRdJP0ZFt52iun7JKnMDsPQhQuzWIHY75i2MgrptL4qMgOGHLir+OrGg+WyUqwcVp3Jhw
Rnt5ytHLTwUuoyLMHZmpCYOJBsWyIOIgAm5qa6fCZgmPBlxqknvBM9icSHcb2eVWxc4nQzi3laq3
4svDQXvFq+Cx6GcPAdXsl2fBUXRktP7PECzcmxv1b0Vp2uqDkuutz5LnpoUJNP80re4/sSt/9She
gwyrYJFhEfBe10sd6mlnzE7dhma/E+PJHKJAlBkCX6VAMfF0tJGynxGuITlRZPeXdE/F8KLLcFI/
g/TbURcxmw4A8EbyJGlJdB3AFrwGlwx+95YE0CslFdSSM3X7y+bBmZceP2869ywYWobbLtLrt7ki
cUBhF6hZj+mhp86hxXdCkkw4vNyayfdPk+OWqmSjaxG1FDm7rPV/z/20J1GEN0uIuyytjTPBkUR0
uwz3yyEfdBDlW0+YmmLtHxTojp0NQJZ57XAeceYaBFpU9SIs1n34Gw7UC5fWUpulJoBNa0bv65c7
9mT6vKNWvMBI0MceemiOHjKvBJZgAWhTPACIhzpeQjVLvRqmczviixVF80dQ5173QAOyFc1hopH+
2pGBw+bKrPDrzehbuo0mYMSjMcIGVYeyWjFKgDMf1i8MOEEcUcJKuvcS7g862XyipM/A2DSbmdIS
pJX3eeYRmsUHiYy1gSz44IPRAXZ4yrzCVlSJUC+asoXqZioi7nfYLsdlE3hIII4osfzUllg66mVW
SRPWXz16rwsLj6qEnyfW0AZnKL3VuzirCQVH8MR2kEv3tbkR4DDSJEjmrTd7065tYWlGoGYGSR+G
kAvVdJsfPEeE9T+31DBX8YJb8flL4/94lju89sfD1AEd2+2owpqy04Wk02+HGieOyf8aVrwFUZg+
xazdmBjuF81ewUGFBh0jW+AxWk0xr/vILIIYtJGK6RJ3uDuc6J5YJlJNi+4h6agErudjyBSCyREp
w2J3hDqnbO1nLqvBjyGTLZOAoJyemNBF8jrivYqj1wEWJpJXlS8Ty8/K3iSr24oRmTnKQYDGOPYq
tEz9idYpcS9eBgSdzYuujlZhvCj5ZnQbU5RVUB5HlvpJM/nH6sDs23Nsd5hIDv9gJA/ds3DiC26F
yvi3Ff0sKnJEEml/Ro8mE3wCjqf+v1u2VKuczovGWnekraqRAOayl0M8OaPycYFfsUJmzVW12WYk
k1g3hT0lEoss1qRdUTzwVYOAXAVVYZUqj+3JuofRKgghtyimJL89NXy032HO6kD0H4fjQ876YrjN
USUeVLgll2hIqQv7NBP0HOYXnd/OEiN94LqZrqO3SVojwAUPCnJWFwzTpOb0IuveYbCo1ZbnhcgX
f519nXJGtpw/OemYcyevZCQhDINmgtxgm+WWgd5Js/Y7gIuB90Gv8O2M2kbJ7g7gcDD2J/DnW50X
mNfUx0UnmGIj5u42JREbftEJ2VC8kDNbRGH/QTOl+OtANCX5Li4mzk80+Pn5WJFgnw3IX6LZl/h4
qB6RHTf0/kwh+/exspLnfCFlw02jBE1OcZ2BIQUTK1HBCTGW4yRe+b9W3cDUiChwru9rQJhB6duG
2vqBfHpiKY5DRWuBqUGlTG5SmONiX8QSbxC1W1cZ+mJHp4KON1lonFDPacVu9+7t21wvUQwzV4z3
g49OxX5/LIs09nSOng6lqs5FKxiGOzsrYOwNGQ/My7Me5SwxwrUsQbAVXKtfTDdIkSuzI0k97cvK
Hq0lUk8JlV+09CY1VwkEnl2Vc55rTSu2JOzJ7mMGkfUy8Ws1G65sAB+8GIF/84eJcPKJFLvszC5Q
uA24eJtcMJ2/kTBOpuZN7pP9tYWBzyvm7uOUZzIEnxewl4EcvfjIlviW9JPAsNegBK6r3cWwgYbQ
kCNNHXdyMgCnyDPVAe7TnnOKCZo44wQTxLkcFIsK/GaFN2vrIc63nXBaXKkP/GgkvGGTaF23Hj17
arU7TBCUQRqlxVgpWy2I6F8J6qFj2w2pPrPSq4KYDwRtGy1uOnQzWv2OZZxh9Vwrnp3XiKe0NSfq
T7inFd+S5qzlCkV3mPmcEp3kT97wZVbsOPsVrh9XpsLfNaygaKXA53UbOIfr8oN5gGM7v4X74wHx
7k0ZHF+CkNsOjLxrGLyInfoOcyB0Dxg/hQTDSeyTSBfkxJod0CBbYLavi9oKr3reAQbRrTZ/zW0t
vIjDhiagdZz1WOLiPnyKFMfUUS4VTWiEHdFFclwNqyvtTR7nUHTZhSug25+86YI5CTK8x2LFd+fq
YoaXZMqVG355J1ipjuORYHucQJyjQDTUJdFiZvd0ndbF2LmOcl/IVt+om5xEVUttOQhe+8U+mxyZ
/mSMBmnBO94zZ2Ir+rmBoazFV6HYKAB3OcvHE5MaqxEjig9YmOv+ZZKAwj3tNlJjZBBksw1LaN8l
gXbASaXnITMm4t7HZw6iMNKdfsMizqTnjrVQ70Twhch75BxvfG4sMmsrIyHhN0aaPcgKaYsz1Ae9
qD4m3MJazkCzupqIYN1Tgabo3AwQQXnBaCnWYI6N5+cc4LnBA0lFjstGCUYc2ip7ZQkG7KeTd4V7
r94nccYOiRF33kbG+pfAYWAaWy4UgPM//ZuLybGifhtD99gcZPoeWjcCYEjTDwWvKvH1gDujRnPV
PPRGA6b3FKQ7woo2cAZYL+hGeTQAGVVjpc0b1W+OpD0yABDQURJMWplph9+fyQyvdnYXCS9tBph1
URn1o9oiKZvdGZXyWACUUu8wK+Ods93k/VY7pLBGfJx6X6htc/CJtGa78cNL4cNMAsChONWq1bqJ
xozCOX/H8sw7AQqOSJ/5BfIboquSplwcAwN5V+kGk99yTRerN5po4hm84Duxi0KfZ6wwICkdyw8I
68kiAl+HjtLMKH0lm/iG7+2kGd1XLRUJSSSQdizkTguikFvbuNamX0PaozpwDcsXb/hGLm1euq+F
N2f+phzfz/IMRs0Sp9EgUVky43mHy18ssx/wHup6D1HguO6ApxJkp6shCkAQu/Pj0rFP70EyFrX5
MuXQYq+n6+N+bb0OCygfjffvuWbnOWMoByX8IGsZtiQ2gX65AF7VB7iy5IXfhdHzwN105aocNN0x
sc2JJje6eav93HKNaBtoEx5z9b/sKFhjdSMJxBiB3DryhvInM4UjJV5L/g8xCaC+3ajsKXM9Iskl
3CuzWsEA+KknlzTgLbSn8HS2S03vf5kfDjZd4+t13slicUdRaWtGe5EfApvqbST2IDRKxPVoiZBh
1uRLrN/CiVb81upPSYaJpFhwkAjO3233uU1vYxdIplGJrUtTIYJOgwFKCAyPrtbz7DhNbaer8xhu
N12keyGmE8+NhTnFP4X5/nZ8cBqg26iwu1Wk2ZInq0N11larLloZ/RH7wr6fyh4TYZOQtLWYOmps
9lkUFy5+/Q9FkAb6ZYxATg71jQLfSUlTe+JfOOi/lRTwT/0Ge3U2xuNTLbegVAjDI8AndPl4b6XQ
gCl9NV05EmRZluq22OdmlQ3PmfRftP02/UTnrOIoV/b+R0WY9cVUBusx+ZFkFvDdKW2s78VjPhjc
+PADhANJy/KLsUDRUXYUcXt/qGJooIqOj0zGWKd3OmWnqwI3SMn8kj4DaxGifOKQlZ1uXJtHRFpU
Uul97/zTNEtMfstrZw0rcy/Z4CCqTN5xAvSw2CBRByal9RqAzvmfn6wdrRy5XXRUcOhpNcjwLAss
q4cnhXsP2VnNC7rnQA4ZXnuMYRaakvRuTagdJWZwuGvrsJWkl6D8q3jvQkSDGmtQ6i6HUUfTLjF3
SIuxYqqPP98mHvIVxXzNjtjD3t1Q1rYOVFz2EEnf3OKrZzqPun9xDgEH5HQPoqLFkbKGJuzhOr93
hki91oujls4Rr6Shix1vJtCXklXS6o+mo/l+OD4dKvQW5NZROk1p8bBworKXb8Lv6t7ltNimayP9
cpQ6/C2BSyvs/dkYxy16j+S4OHkMuNJkXa+9Jdokb6qDxLM2YrZtXt+ogP+f6o7rlbAR7xjZN5Cg
rdxcGzVAAiHqj+PKzMoaHgskDDkNCk3+b34Jj1NGxnUwRk7HzmNXKMI5PFn9zxye13IAMjPftPWO
J2CCT39ykCUI5+WsYYDukJiTcDdrNggH6wLVsI1OBL6EW7q0c+r6mgTrNrY1pys8HdQsrliJcH7g
V+xCyLgc86nUrrCxujFohVtEX5IFdm0jAWW6H3OFjt2Kzm6zMStbJkP8TXGQILBT+PbTZIQkp3I+
ta2WlsrXeh3dV585A8iLnO9yX0TH7macpE9LFv191zV2VB5IM1bFzeGfsIah20L4DolMyZULcUtY
gEIPiOKKMzO7C6s2ST2AtQ+ahJ145IdxkMCI8A+H/Q8nEhhVMBXvRvMkmC2Lly3KfS/6AAvxUzXa
X2NoynuMcdnHsHqNUVSwk+y9cAL9ihLl7OoYO7kM9F3Sz+p60oP/Bp59Sjld10xHrcCLBA/pahDT
Nr0yz5b82YimUPXwED1yairZ9eivF3ZIF7M16LKOaKz2UBfpCL5eDVdVVLEvO7xHk1Kru/CRvX31
TvykgZ371wak9joIq3axhCl16J3QP881BUb0Fqi/Lt3BlPk8Jci2FZyL05k0KQkdEHQrWfQZnCTd
kJkbhpLEUisWm5Nsx2BUld9YJUheV5pSqPKoX9xqLPXsHBbuNMFDUKq9kYYVMyd+e6XuPP8Y9Wtp
cwHgHaaGtsUNiEww5aiq+OBfgnNS2bJdtSeAVKyxTOnfWROOJqibNSPIv78SpjhH65pxBW/MzED+
LqPlP/RPoRwvbYnQARerUPKMeV0BWKvm02zQAe+87t5OWw85ux5U9qtOP2Nhcn2b9t2OM1h5YE6E
Uw2HzjwebOk88PbF1UFXVxsin0e8gJ06iO7mkExuDfMiWQop6efUWe6+YUyf7MmGlkXg5Cab8TVf
UwddifGsZx6Tc7GS98OweLy4PRB/I66xLDgTIhDpBuEsK9hscQy9RT1EfYC8DSsZGf1vWHv9RtyO
b28dI1pr83ya6ElqTi4b4zP2gY6WnmKooghU2ZMIYnODwM7seCxc13DFFxZJ50A//xBUU5xSNwTg
sKaEJo/bodqksdJSOwHnTDXxmGvMAtQq5yNIZbuem4Cb/Tg/KcTk5oKF/4ApgFelKYgvtNNqMLlY
BtVGsE62Kw4aJC5/5tbeRPZ+ELOlQpTyXsQsRtTqnqbsanp9mc6ZpbdRF39Nq0GKcw4EC59IHV6m
7RkkKTMyGBj29xkUm/dXx68lKH4xjr2dhTUjVO3crTtFCXlryWFTUBVDdWjAc7zMOqOserxDvbLU
/NbGcjMw2cB31BVBbopMObC7dDfNVDov5KFwvPBx1iqNQe6o7sXhDtL4jicPy4z8ity9ttQZm00Z
n8lqC7LjZ+VnyGJuXK6Mvy2qODOhMZZOQtr+UBdwxCZDm/3Tdh/WapUCITgHELCSXM86XlrC/Pip
2kA+EesNVYggqaSVuFK5y61CV7tPrZPmLGQfO99tIjRN8rSsCRtLF8CFc4Tkx0sI/wDmQzPwRUr0
DiWdtU4VkokXqkcRceOPOelxn4xcST7QFPkdUnog7nnvCI2sbj7fmp17/vBLRJRYorckeCkc7p70
EI3WJVOFD0zMjq9Bn4SuaFc3Qt1PehtrXj8FpQnsoX8WdQa1z4M3ZLeO+NuVUnsfDFrZuaayIJjf
OY22d2keeJAT1VxSPjvSVc5PJtZCIHL/fcpzgUHtarqmqw6VHdZE20QMTOFaIDuka1gWvNDQAZ9Y
nVRWKa5XafcyA2VnAD3yiSRhBZ9qpqG1AcUvTJwmVSkyYu0k0W6Pa3o7f/TzQkktIQWdMqa3IN1c
olOo4/LAeZFcKNWFU87xEReanU1JKFuZAO02Zt8wl8X/ujX3zkupbPOG0lVId1ND0xEbxb1uIJ1N
s9DfxU80MVqhpTyx2CYtaVC9K6c+XdmsC8PwJSxlTJTc95yH6PVsqkCRTgAWHfnTE5ig+LN75olu
n8Hxy35ap0YboYO/J3ySgVp7ODYZ/qIuU7jBb8aOkVwmm+6RdElcYl/94egOEYtzXNt/+iWgUQE9
iE5f+6x8VOB2wa41L3+VODqdxUYX5JHE4R5US9y3RRhj8IFxz2xfYE7dilt61XYE45J2+T0/X4cd
kXVAn/DD/H7EcI0YyasnGISfXmAQ2N3iv6FFu1H4lj2Fal7wHLj0PPenSj8qAnXOOX6tesG1Njy3
jtZcbTmur3wtTeAjNcBFSRNQEqdZznfoGIdzBGejhCeeJoT7wW/H8RStRGY//Qjl6TMoBFkXEXl/
x7K95VIB6YttD0Y4z1/MB2jfffF9fqvlDjfD7kTFOLIiLD0/pFFDuC/gWq8hQCcv0u9xYWK64RBN
TY076BGeVEbgoDoRBkismtoRg4brfTvzd4BvTnR3I+AUsL4ea16K/jf6F+2RxY4tr5+SHgPdpqjy
oGwhQub7wruvXXUHPNRn5eeoRy1ahU8bKKD3cuJ88DZA/3K5hLtHBA7HIa0y+IvFYEjbpWDRPuny
CKHv/KS00AF/dX87AabPjZdIpbDBi7TG3f67P23hBRrvKYllbPyABQanaR9rk2DXaYiPHYhfJlip
GbdOQmtwKfZj3AuahFF6uM2QoJA2dNt1+tu4nXk5xx+m36satPMbUgCuUYZVeyCZ0wAubQXwKcWo
A+56fJet39d+2inIUAdmpNORerxBOjveZ6LEEP//XKZ5riBSPp+JeRtvuA/1WFdYyfNxgMC0Y1BP
GC6Ki1509wdbQARq13+CUkw2s8y/w3eLg5yHeA/iOrAZx0eoDeG7dR1LC2ePzjmgYx1h0nHbLGdN
JyZBaI1lVbDIUn28DXIl6q50Y6WDZliLL3wUCZUF7axTQpHZEnriTWTY05SaJL6NddzdhRZy1+9l
PEvK7HaPxz/dGvm3YcHIdJit63mLbUVXXPtpg+9LYWHBvWPsACZNLamQCbFUdJ/bolngiwjAPIrn
4QwJdiGuPTK/E3Y9QWrq75HBBPJUeiDaoZYJZ/Plglz1PhEvqdP+bjFKH/3M3PpCtFvq/dqkE7To
ryLCHPETXFKlCrc1RfFFcDwN9rd2zcy53hsqJcacbS0Z37luzJncOI02CiBz5eT6dLTCMTk0b3nB
3yE55Ws4djgaHyYkTWhyR23zETWxUmD5CXDLXD7blJNT9tuAbJLoAiipV+RHNbheWRcDSrtzf9uS
L7SvfwGNzNRjVekMTMt4rWuRDYHBB/FFfAFAAMy5EeJ3w+iZgO4AYfuyv5TDUMO1OqD5PmzdxM4i
niL/wAx4t0CjZM4Zg8LBZPR1yeN4WXioNGcUfyTrxwuxoJmTZFQ4wkYbcQD+4ce2tledgOxFxYGg
V63zrvNbuYry3FpEs9y+C5GOyc6hxVAE8ERKQDQ2wCp98208/3zF2Li+jOnmIuyVeJtkPtxTW0sC
U6upNEeClouSvPqxzw5syWQrxVM0akMfONMSyfpDwhksvOSuhJsoivit3kc/PHEtztznDjhqWn4B
TNfkKssDp+YDE8kRQ9WWYwRJcLDcZkZkoNRfq0G8P/lDOnJspRFw8QwGTgDbJIYrnAC8T4v63f7g
3M2GsR6J0HyVm9ZG8vXT3XKZgFQ6xVCcM9DqVqm+r784lBxmfTBVd6N26S/awtdTAkXEuPeWbT3m
dzI804xB7O4lOi3PqKGGh0IiPQ2zGJjMZ2EUg2QAqHDeX9OX4s2kEOINe68sizs0fIYKGeFi553L
DzoTYOI1L9kQ4rXBX6WR+fTe1c4DodAFo/FQ0eSol4GjGGTbKfGlDLRhjvQthchgEcuLNlhHCJYk
wr6rbRH7SNpf+syYxSVOgmRYHL7t6wE86bDkMLjGnxtNGgf/St3C4exxZ0BeAJZF6o0+Aag9I+hB
U4tPnfrBE7jPMpxY2jsmi5mKTy5o82X9yjWnKr6X8Yp8s+9wpYCSjC/71at+585GxBmmayo8SD5m
Lmxq5JJlHP8nWrPKnlW5mUWep5NxnmQMWRj/V1K4BbtwF2VjMl7MPuC3U8IqyBdKDg8cxBRuifn+
1QZ+xpz+al0skx23s1zbAWSQmNEC1RGDossWWQJEtfUrtyh7CfMq+g2+HLz96W6PqwTbD7O8RvEM
VxTVY5XBPhPsf7N9cDT//5C1o86njQg27xGUXv59mGeEnCPwA4WGnZxcEVxx3CCQ2cqwbjPp+z5p
teC70dRmay4rOv1fl0cpOjzOBbsQv0KrRSBWyOMhBU1ViHGx/c4v+goahU260ZxxtkbiNXE/8Ozr
Mgbbzke02mUgGmsreCvkObw+ILPbWEvDADh4cnjlopOQQTmZSSZeYad1Cbx1CSLqbhuDKT3b13HI
U6eJpdlZgQzDW0EqBidOkPNzmF9uqC8HPh7xwNqe0ptOXtap9wEDYGu9SW1Kf9qjeGk8jC9j81rB
SHoOl/bt4EMc+GpoMlParAtiiew6CJr+nrykJHhUs/9RwGSssJV07UPCSBzvgD9dGvuTpDZL6max
QxMZCEA0IeWNjq7+zV+efVXjf0Aj77tSg/1XiK1raxlUhOYUTMEZnrL5vc1qJpqKEZtFTeF2zOb5
7AcOqVOxkUvU33iCMRcOpEe0nNEs5IjF+zSUKEeqANJ0aEneQLfN0Hv94QoJH5uA7GuNE6J2ZpyV
3ZNBURNG10+/Hb+Q3bWZq1HSXVXbNf2Rxildct7vjpoBO7+/+NsBZ8cns7Fi/jSvKNqM6P71bhVX
y9i9YTAqnMK3+SZWXTyMjiVrL8XfjVb/T2eTKBBpyYlDgPt1RPgp35b2ekgaH6uv34aHPNLJ4iHT
tGirdxYYYahQcd2cVlaE0SLz3RH4fN4h9QFlhIoeke2/yMp0tpY5Nlw88nviXLDmmsmAuaikH66B
JrWesrNTk4AbcJbzwmhocx7dN46aDLpdtj2F4vm8tt9AHIxvtMsdDhbGKyDQ3/XX84HSgeWyOi92
2KU0UjQ+41oD0TFSvUZ2MGsLj7rDLBNEUER0nt/B3qZeM+ixbuoCDPB4x6wNOoXcgkpXlQf8fFtu
3X13/I1KeeumR2DlEy+V5ETX15xMB5KBG4Cg5uD1cHoNb8TZuqHXbMdGQJgB6PAdkGEMlM1cNwpB
TcUKZJPfRoEa02MInXzZnuOkgXXy4gDncMlBS74IBYyV8hcEifLe9Sbnh0rFqHy9n5/5l6cSk/88
Vlgm4udF1V4dZg7JAKDuyZdCMoKKfIMyr54ckTZs9PKFm2CEcS7jUPMOci0GQMuxJS6//m1BPjT2
t+mPPajdFkDfOIYwIXUIrMClqLMztrqzYESw82LGRNZPioMJRU9BJNXonnmykOfuH609ES9rTIb6
enXWEuM7oqkIjmFAr7chSDDrSyZDU2k8Y6SR91fS42O3eJJvPHWG3a2pdXBEPlJuQlcowYk0ZOiX
u1BCl6CAFnXCQdavbRb1OV7E0ACXY6VvnRlgu+4KV1juv9qEKJz/5la98+PRGVeFzNTAIou0w/ud
fB46t/XmEAllpJMqJGJ+zIUI4GHUo2BLfZuqz/MDdu0NV17SchewQ/g3nE4h8M98TPYTbgq9tXtr
dGOdeEEV2DepSBoGdgk2wWvRsjMFS7/loOq6pA6onzieBm+s9rzkUk0x2ldjjla5eIe65ue36sVK
vRRvQSxUQ7U8S0jDvbfzE6qhtUlq/n03NL6Rvw7pIPf96eVFls/Frn6xTH5Ig1DmI52jO9evHWUK
i086KcHI78FFuIL0jAaiOmnCc40B6aiOfSgLs6zaVrrgFgelEVh1Kjo0iETzDVLZA1RW8xnYtgju
nae6ucRptqajPup9ARtoFcjA2tMbOCDRkiUAZDUd1SRDo6VMfR+M2q6tp1b3cwZ9WNr1fRO/2JBF
imuF3fsqkcrAFxJjFfrRmtBUaXOmqdFBGNH65si7uagXP182TC237emsFnXkdESHd+Hwuj6NC0Sy
lGugDThYPtKbd3O7Wz0k/lVmf92QZ7M+NPrh24JkvsvNlTbw9hLq+vkMbTCSjU4ETaL1ZPFgWjJa
P71WLQuhKmXSK8eP40lE39eFG9TIpGFqpXvdTZa6kLQojVRfiXaBOeRlSbfT94K/QrrefWUGwBiM
NeBhqNdMu6Amy53BimtYAAgan9GtMjTYa9Os5vEGeo0CXcWTZDb7FyzbOf9YUXguKc6riMJc6uI8
tLiJ5YQSc/4oUdS/5W9al41Ek+jdnrvJn8sE+Pc03xfdkTvG+Gaw7wLjDyRAosdJXa+LQ3Bmk2n/
V+HRFF7DtFQL/asMwBpGyu794YL5mxrE1/7b9g/IR4BQ3dAoLwivs8qrdLTcpliQQPp1ujgxL0+w
EbhBtOtNJr4ixQOhyEfcaAhuijU7MZ7TOjzuxddo2rlM0uahIpw3tMSeVtmeMo1u84xMLKKyvj4v
7m5bACQh7uzBDbYPXr5vriq+434xip9FFTm20WCBK5owlOHpnSw2gKU/WB0nut/lFXMm9vxuEO12
ROoP7eVAHKcLjc/N3AS1NxNFBHEs+eEz1DEoYouXOZlyfmsAywwFjH5RRdUbM3JoDEqXZrViz42r
dkNrPI+ajs8uqN9G+AytNr4jwkADeXRX5oV2nsRtJriv94VdQeu3MMb5zopfl5UkXmm1N674fY0G
LvrxF3lzokx8WTmt3M8+eevtf3/Jn84FIUgjmJW5HhRA6/Ar4j5tKkPfWvu/yxid143sYOMZsfQF
xlkhcwfmYIlEaSyqUWPRFRc89LxBBcIbxfWtAWHFl0xGMY4NeFo3HIaZJhF+PZDrZfqAriobqoiE
8W5xBprR6kyR0DNu4USAzfA2ie57G1tY7Q05FBa1QDdu4YnNJaYi9/9dCnNSxx9ZU9Ai9Hga3+rp
9NwjP7E0mK8/ssfgv46k9aw6v7WCOJaDKr8BlQ5GzJxLlkgrD463jNyd09BTVv4IGWTNCNSFjj10
3+TvlZ6WvZyuPOfCZFwY6ftBpY7gI+2timYqkvZVXOEFalw0uPIXQUqsgHVgDE15+iEeCWIOLqJw
yzmrOXEo71Te+8E5PGD5+3PDDWKigOmRCtd716aXBManeyvFhGDAMkLSa1R+Cbtk9fLwyPBxO1Px
O4gIKzRTAlkFVzbL17UC9eJfIPUUFMqLHZqpK2uNgNM6J77fz6ohmmeygV1Ujw7AISO6KpTUfUbB
X+p/LveCIibMHyiylxCD8TMwFb6g6J6FFeGEs8+WG5m3WgiLOJc2S+gswNeyPWVC3TGCPi7/tBbT
6jpu3S3r7n+UiB3b6eYX/0U6gZwKsXaXqaiPkcHNbUIe/kMO71QALeZ7vhZlKskz+W3OCsAB8xJr
t72oO5PagvLzR0Qdk/9oIc6ytV5kZdHwTQLWMuVi0exrtzzXrMTVSDWnIhnNItHfzw9nfy//8dAJ
PFL0TfqO6HqTWT5FGTOgPs+qsxqSVlCJONGoHZHZBywKpdiC52xRAc1BnDqv4q0LRAXdtyp3v4PL
Wa5sjSNTF7a4lckkcP7v2H46Q1Rnz/5QF0cfNNfHi8Xh6m2mtlg7EJwuSJ3xG5Ox5Puvnznd0IIe
tUzxjK32P+uqRlu84Qo85k63u2CF3bVqsMUsEJlCCMESqFrAIIUVUZfGw62flZV8MEXOmFe6NGHY
VLoHOikmJ4oU9V3a2MmjOZBiMGqVa2ivDhK/s3SabSL5Q6i3bIEdXmmZkbjODwLRIigA8O73djdX
e3iqmMbpAkvZH8KcUAwUaAUI94qAHv2ag+ozE3nSrkOy6gvfoVPRvLj7r5rZp7BNdk+r/SDKaJdg
5WdYvG3U9GJN2UeNps80OQ23BWjANh+FmOaCsMOKAJyS+6gb96gmAZRLJbp+CWcR8bcetNe2Xix7
xjQosrNp7z7FymCXzAOSt8W5CGnwMmg5LAJFQ+K9pOR6zb91uJuGDm8pQzLoIfPEVgoM14w8RDRt
snmj05hpF6/M9+yMQHjv9jljqmVSi/6Akid+mqso8jGcoA/ozT+1p++MnugcXVtKevBo+jX+xuFd
aqdLRpYGN+MsXf10kCV/GhJyWxUwUcGXMG1oWUsTdnz4XoXm+reBuWBFYqJggfHbHBfTpE0fIqez
XRn8y7V0c7eESuj7RONmAmZGKTabMapwtjPsEb8vidka7dDw32JxTZuMlfiyY5gBxiu5mFsPIGI6
gLCm4teOpbgU7sgOdNsaLWcQj+U9WGW7m9EbHe1Nk3/mJP0ZKL7cdY8VNsk0sUA4cId9BYjHEW22
6OK+Nr9OhY76w4fIpNLtVLnG5+R1jVtGTrkwcVa8uqvAsZ9fKpSVBOkvKm1026nE9BdOj3SqovMX
OusRIuXrwg3ztGfoixOUfmJgpTsg2hwsNiuhWFdV7hz/v1IjDl8HfSZ75xUfxM9yS9vQ4dA3E9Y3
mA83A2I6bwW5SbflzJHP3cpBi4rv6Gjub0Jlhswuie6c/ZHbZvWoQDZ5uHUANusdTNR3sf+IfWog
9KY9gV+lK5I/w5vX4MMdc6cUoInIge4fO/FMEHWm2sV7Aj4XsQ52h98Lpls2HeIXbcjR7ARf6oJz
VJ6w+Y6rQsQL4vSXbjwjmbOjx/SPQu+6StaNu56EAZWHCj82HtjmNPxMc9a3OXxNR4VbO+knVJ/J
YO3Ne8Kjyd078qRGebEo+UwyUQV2gVmdhB+UfMqcEaB+/C/97HZeFdknzKIa8e069RqUG1jFK64Q
wDIJdnHb0OBdZvwEVV9lZb9F2lVbMxhR9r3Lcg8yR9vUxshJ4jUnOtssXIbSI7SqSm0JdmFYsrkZ
ah1PFr6S7DG3bxwocDa3FcVwpwTvZJjGFm4mI8nh8/vwvnODbDcbKpgT21oOwM2NvVSwyOrE2B1i
HrecF2brDLJSxpljCtBpouQgmGNVyfRmmnTLitLc7UFpyIgXm4pcv3SfUfeJ5QA0ZIOfqQMHEZCs
rvJilO4lygG3lYoAFQtMKzcn/kJqOPUyivGTGXq2qXbux29JQRRiCzDOlmNNU1V26cyS2+H5PVgH
ZgJXNx5aGUFbYieaLno4L/rbAdTkS7AesA56ePcVY8MXySUz324gfw/NQ+T+J72kP+rD19IokBEc
X7pH63Ocwj+8BLLdCZKa5EaE8FRMbsI4V8JqRXuWb4WuobJdBwIFmyoxh83OQ0/KrYWSH6DyvfRx
pSwcVAyKF1sIzd4geZtCQb7xoWwDtRFQ2v606ZiNPBNAzW5ws3UVq/hc7ONMW7DHMg9E8Uw6rt8+
Xzlf2nLLKGawyoFwHBdTkmEDnoPRBk3SsOQP6D4pe0yuiCcg4pmsW3iWO6JhtUUx500A1LRT2yW9
n4KZRHCKaUJBFvbF/Y2oGuc3MRoAMsuRnf437GMwY2vrOk/8HyFS4Wsep5rnuQK0Qf6dZjn0EYUr
oxzrt9UiCWstukRf5sZQAw0uZtvaqH5khE+CBQ7HRWN8JWtRoQ7MWH/4iZv1cQugqjPSB2Kz8DXn
hVhDTcRPNWiP3hH6pHaCCBqlcXh4dIoaYb8KsQLrnC5YEh1SddxZtnDvYpdsZyh93Yw1FceBKrpn
ozyh0DDEOA8kSjvbtECs1QQjCjRZDjMYevRM3XfK1OXGWM/s/c36z2YzTtQ8YtjwXj1ZYQEMSdwf
cOaY5NgSe16IHfVjpFolPZsGKW4cUnoizTB/Lql0QCdAtI9FXmbgozja0o+FLdg2/vrlrkNTdfLy
tdDEIa8fJs93ONQxj564Qyk+XTZrJMAgILQl75pXEe2EKTmIirMB7laUPMccDS2n5vCfUlwJ6Wb9
GI5yAixFaeiz91/RL8eXg1f9wBtXfDgdA3RFh3zRLeiy8gvWiLoZQaB9uYXIsuiToYjjq7Krx85G
9F5v30OhJndk+bjzQlo3QpDXmET1wQ4pH0dQOPjlydIuTEwB0rBoxJC+9RNSaXm1ZwBQjDKmxto1
jWoTp0Vd4+HmGO5Mi4U23woVqBhnNUg540KYNFuR8UuGQRxxLszfx7MLcBJaHbqr6rey1nRV8fFv
s50y1YTwavJgQ2O4rcmuo5H7NpdY7GOANXTB6iMkI5/bUJF0H3cZiUBXH+Iz6HN1GIawQ4nCmuO/
gVoAiTWaACQ4dSzHM4T2oEm4fqqlMqJO7UOdDe26H+QFkt6jNnUWt9B0UKc1Z5yIwwnc4ra4EStN
lTh+R6m2QcDUALQagRIUzltuRCnYS4TNubYOKkk/6x7HMAi9LESFFrDicfg/j0sQuODDkH03BNmN
wigDxA1p0hhGlWJ/mfsSJz/V7+ohRuBPIbBErZvH986B/N3r2fnFFb+0i/splrxMgW/FCINdDI0O
ijwcy786sdOGp/It9PUL/T3M8Yl+G0o1STVwyysimMZsF/XNc+cknk8CTkAh/i2HZVtB3kBhND+u
VyiaMw5idr8ZF2gISBOupEX0Fbo/iLy6gjBgNmD0gWLgjy3hl22lFZ0snY3fxhATIYo7wc/Xjzr+
Zk4nSAJDjs5akYtv6PBoPMT5Ws8tj1mtqkCdkaJQ85B89PLcGiWGNx3DehXgmERRZh/CshykDc3K
UtEK7ij0nD0gvYSy5t8jYfS/EtDoGJHod1zyIn6gSSfWcsROriOv67NKhxn18IE18Y78Q0YaARSm
WXAQ5G/a5qZvWmsrcKxyH+RCFvJ89uyaHFGOgrWet89Dvu+YHSDzRYjAijOmdH+IV9rcAvdbLras
5vYDajWFCv6S2LAr+Gp8OO8o2hPa54yzC3Egrc1ytczgDIHdUk95KC1zhL51Xr53uanXpj/u07dn
tayKicmfidTDt51Zg4rYg/W+LZ58qgyZwA9mbtnU2eUdcPsG3ADlgYlN9JSaIx3QcEfnnUxDI4Pe
A6HcWP/sQ8QahorAAaD4YnR7C4WzNShrT4T+LCKfguFye8tez8A12ljteL6rHY6P+op3RYg4Rg74
V56yJjIWr7/ipDl2Z3U9ZZUMQYpOhcUGSyqLTNo6fy3IkWDj+bKhC54auiKZLxhtHfS7yyxU+3K4
1VkIWaavoNLj48+CUXzGIjKjZ7jJGuaShFh6b53o+zCTgUo67O05W99lBK4qOohQBclrHQRuvRkI
rzzQ+FfrdeSqpOD0XFgrDkHOpMN1x6fy9sg7PpjyYL4hNJ+9oOAMo2C3L9Wm1RWjie0gwIavnWyy
5PMLfcWMl8HzES0YdhoTiOL2PsNVABdwM28IrewxPi9sUj0Cuz1AzxbeY+yv9E4coLd3/N/brLDI
0PfXs2WBkfv2Swe8RW7wSPtU+dWS+0YSlITMAl1une8Smjcqs6OEftiSe/Vt5BxIzm7CgwSTshjE
mtwfwApH1hO/T5fqf/+xcksvX1qBNJePu4XsPFRvQfYHTtXhh40Yl0bKU3czbxmbsQ6bTamd7PIZ
3xa6+h8sdaBDBAcPm2J9oBvNY8RuPskqAsKVDWDfaFyZ/YpCondYSrym1EsDWDNFW6WUlESpH/bJ
giU289CazPj7QUyiJXkJ3U2V4vMY95ELQikts49Om3TNr4w2OuCrB2UB/c4dOkNRMiZoz9ZCFrQL
Uurzc7pDlVZiBWytQLj2s+KNn2YCy3H5naahq/XlpFeXSo4Ap4MZzwWZKj/lHsf0KNAaEJx1/FsZ
OIDOO7j7GSQz6p3d/MkdrTgKBMw8TB8y6tO5uQn1jJ6mr9n39Fb45M+tedODKWWl9MisvaoD4gp7
+I7sbFj5VMdmMfV6MKEUh+TSBilqCIxCy8U2FWDz0xdN9q/Fz63ygqPsg5bc8EAo3mwbx7iusBU1
/TWMXj9BjPhU2RnMgl8iK8fPp6OCzV/45K573DeNZ72/FcAOArWnb+q7W1m9HFh4Ja8bEdlnBQOi
ZpGC4GbhJoCZC/xt6HJlS4QOpPgn53GgIplzLCqFfDUvsjp+9h+vuM8Nsg2Eyzh1cw1V80BtfmfS
z+0VXYkNsSIIyYIQbsHeU2QXYSxIZmVhBqc/Q0UPtu4dCJX+yENsfP+P6Bmx5n+9qA6jg6/6HbNf
g+laKfnUaQkRW8TMSFXoFl1XNCUm7jmCIajkwx1QYIu9mYizJRiUUedF2M0pZ1FG41yYijNu1SEz
cOn7H+7253AOeexeUTHKat9n4b9Qf7N5YbzqOEcLLM2N1Vu7yz9YDXWsBXpoFyUhTmEwaBJW80j0
ng1L9Ol6T6k0D6mjtPCa/sBwiERbxZW+aCMb1v3UVsciA064qVotf6JiqAjk6pcH8Th5wmKEzU34
lEhzMkk3Ltbxxw1pQCDoVUKo5S+irWVppcFYFD+m2cHG9pZ5t01L3YqdmY8pecx0TTVG6QMk8wzu
QN0TQlL9Owa/7SOJVCxypMjxCTLSGwPkG2nrQuXtFVISQH7wIX2dQmXc3BSry5Fa1/HIZVENorYw
dQ/IgFp4OWiKuPalHKTXlzOMvDwOuaSmua9LfxenMiaseDaKFlO7WQllW4JAHNgkv/VBL/F77+ut
LsBFPvvawSgJUTLO2dza3NeVhxHxzbUE0P+nDunucUY0WX9rnmIs848yPwZKW0mlnlMblNR2mrj3
Yl837u2+nIJ/lIz7/ELnqhBhiyfaa5WjHWLK4NvLKkqLa/2NULe/FcFcJeNebJWASeRIFmfeT17S
1iW+qoQnNa+u+0ntYt5ZmBjXGRXnYQ8lWvehriolemoCXlPMr8a07yZdz3W24xEV4I2AN0Nfeu/5
UmO+EjHIARnMfqoNIrS6CxtQv/oNSPO9Yd3L+SATYZ0NsTTaiqhMQbAZysKSVUBOFeaSzJPPs3nI
Huw6e9CwcNP8H4Vx7DeCu5ASf16iLJj6scbnRbjm79Z9GHrBlwrje2IALrZre9Mrb8dFTT/Q1UIJ
IuPzO2D0ArLEajVekdCJihOtfKkoz9adEl4MRieKhMpMRrj6YtkPeeOLZVfki4GTCnWzwCCE89PI
cbpmPyfdoioCzhYj/+yJ1jyn/DgCFxKdoOhd7aOkbzcZw7UhmgHmUPOjNJTPAsER4yTCIHQosw3E
WZFxjRTlLHYPJ+A+f6fwrLjg66WYqYY7ainKPaoRPTmVT1W7YYtMVbBrjWxO5gRE3TL/96GEQ7jP
2QIoV/TCmxMI5xIH69HPY0um1Q+wXLfRVBEsA0FqAit2vU+m9tBsi+pKZ8gwFlN8YxAzwAjO1rR2
/JHXO1tHvgCUB8dLGmQO711IGGM6BfVyHkaieBZ6GcGXQyauth8tGvmvfm4n6PWtt3GVDCz7/4iw
fUKCv5wpsKiBu+poV0NClberwEzCNrUwz6W6ThCE/QuR/1Q4XR0p3rGW7Uj6TbdUGWWRBE9y2JLV
U54pe0nN7rLtmykpAeniS6nvvcUff+I/5dgzerpETt7HdwO/4CUlFJL/RyIuiYXXgmFlPFOESlpa
iRE27Y9jJAzbxpWJYdE3LCfCK4fBKPJUwhpPUtsHdGBRJbk/sZuyxiGPcPnH8WwTsZrMhQkB+VNS
H2r/ivpMOt0DZPNQLM00ecHzMIs3nXHHNse8IQrSQr0jVBQis7sREhgTpoeHT3EEmSAr+Koa702S
bWDPM3gzMJNDid8am87GbUaWODCIA7EHIrZVxdwlfXoeUYqYyXllG9z22u5W6DIWG76QhqZJqTWS
iVRbJ/H7cPXIGk8iJHOCnv4gVtOd6V7XVc2CJF4qy0ItbN0CQV7RZRmiK+YluQPdrSNJjdPCwJ92
LGqb77E4iEw0+ND0D8/MNjoiUxgaJXyl7Cb6KNqmILsRfHCxnVjYkVqRr+TdK0rxtw0uPponKZSw
zr8SkDYuO8nAb5OjVK98xlSB+p7PRaVoNtc2R2mjCEGGcrJ5zsk8JyLC/UTo33AYg1z996P7g4RT
tPR2RI5TLcwLRAlOiQfRSXnbKWMOnLbb6K6xeAa5YEYBtv3kD1wibPhnEn+z7UeE1JWqGVCKQCut
K6Q3npQ7WC90Q+pf0NI/+PBEn5xPqDhbiYwCUO2lobCL2iyKM8EqWciMABsUbgvJzLI0zFTEc82T
KnONPowiBeGys1jtSJrurH2Nghu8pXwABX3mXqCnKTCCb17tXsDLexJKUZ/eMmPOebC5BXrWeUea
XCswYzh/gnAcvBafLURmJcpfToBefNceo2TCn0RI8+KVCORgAeY3MOYpysrGlp5M+0aMXrKkdOYK
2LsrZXwepJ7WWzZt58OILrG3cIjazRwJCu+bc25n9Tn/4551Wf9500cUzeb5+umgJSs8SlxnvF96
SSUnUIO4j8Vc1Fzj+PEWGpgLumFvogXgiWLOxr/d0s3UWsDrhjxIi2JvriOIb8EgbIoMn7UFUxgE
1CMQ/mgPb+Ul8dwPXbLUr4sqP7yiGD6wk9rcuOlhOJ0qnHzBMqUG7VEuzv98BROSddlpOw5uLFsA
xh+zIaBXV7knyQxc0mi7ylkOzz8C/+7chPRASJLevfgdmP46rVw8s7kDEl8REeBFe3+QIRYa2XKI
4URkP0xh4embjhKAHJQ+8l7fuyl+qH0rX5YkYvoG7BzRI8H563H5cK/gzpkncrIKBiqPSaHb7dvu
+p7eWV15Rcbn9OZOmveRUrK8KxFC9hkFH9KbdrrZGZoIQpv5349tB8KlIrwg0RmZK+hbStRN/1ke
vGxVKtOc7gXGsrS1z7YeJg4VRe4xobZ3IAsDBt2toX16NrZjUdAE9x7oUUOASRN8POWwFL3KChkM
QHIgY+jzcEWFt8X6DAWwFyG3IFcUhXRpDkNQuGYCpHYzlw0kPG1orx5/SOsdztv7jytqYYtXmiip
7nKgmmyJEpK44Cczon4xGnIbxScdlFJqxu/Ka3O8ZFPM1jVgZZhv7NOZEkQ6IqTLjmB8hLX7r1Rf
sd/esDfv+SXtPTk4BdVq2vSLA0Vi1F/YtW0vdeOU+M9IFnVVMV/tv7A7lxNyQKLj17vspUG9eQb1
n7XPWZqtPjCCTN+BHo4hdqi3lWntmUeveli8e27XIMrKTLDEg1cK5mMdmMIK2dX97hOVrCAoZYdC
ELO7CUdqUzKyLx/OxmtW2DYIccHi9KY6bdxzTf/4vv9AZHAUFILqrS5L9WLlk7C4zlualTeHlEUA
I8LaEIk7TASqOdY0kroGC+4e3Ao19t33okvCAAsXf9DPX6/c7rc/2FmJU/Z73FPlLe3qnENyiWQx
mFp4bB3iuC0YNq1i78NbhxgbYC/BxpmrGsOmJe8WlhJSHAKEN5tlNANcsbwcyZnsB2n68GXd+hzA
lncIq5zBcc+RnsnChsyykiT6o9KvrVR4OYhENJSa4m2vr3fERCwEIvvqRT7cXe8PCEHwaFfoFGHl
to6QDlxNGI3DThLyLOkPxPWfAQ+yluhGGuGK/8Yp1T+SG1q9Lc84yN1Z0vaO+uMmC+2+sD3HrSoF
eUwK75QR6JZ5vjLbaRiIGEGaiMeSPaDveQSlI0zFlUBnIIyQqY1AMxsHbML8pXSdfM5uKWFP1hV9
pOusKx0x7mA+sFOANF1jsLgLjvkdnV7GIM0PToaWyq174rn9vY0Rk1PkPxyEJFN/ALc/wLy5c+YH
Vv0z807CmOOEgVuX2eBD29rrdCwLj9uvZPD4PlWM1npb3DpyC1T8FPItkKz3FvmPpBlBXSNSNhem
ltgFZtSBUu2SOPW+koOkZVfuqj1BTxuKQInK2Vb8wDI10DeIki0QZQC3/OfHZRFTJ09vFYX4w/c8
4wAXb/5qG+cbA6Ev/a5uK38pB6RrL4ANB5UUoqop701lcNaRLNlGTumExgR5rBcnvwvA3rfvd/81
/Sz7y14tFkbF9tNz9dmtkCiaatzQUFAk+mi/K4RqurqueazW1S5nppAPboZcy1JPtnN2l2lysuE5
kqS7x8f0R3t2d8RFksQMMjdSYtV0P51g6+MEt4vkfrf/yQxwx2AEWkiphJPBZvZO89aFXTpLs5E3
L2CwV51mrVDuqlhqGDeoq+lczA0crZ624sH0rOnfTR2LcUPpX72uq9pmVCsDyAvzGqOxkT+X5mZs
0oZ0mJ9+rh5gOPzl1RoKj29h4n2P2zeEMiAqOlQ/rBntfK8JGkh6l90ICY+dXpwswp3ZAEnkBM2S
ykt8HshWr6QzvzKeJg4kzYGO3WPGhMBEWw1ElpOkiwGMI7BwCVX5rZWkYMLBJ8ffWrXIybMPChxP
kJuCB2J/G5Wq89Q0F+qxhtDxJxB2JppsDdOhY/mGRszxuD9yBAYE7VGCdDpz6FsB7FzLlVdL3Iyk
/gCVSvZC/st1nDyj6PfdFHuNtcmhBB5kKHguxPxMw/MFp4EM5AFE4QdLp83TC3ZIsrZkGUTPNXB2
j4T5SGOMAq7DaZehWvl/VAK2ESTKzpwzNA7osUT1TT+F8TWZg+zHLwvMVDa+skoTHtSXy8hUsCNu
2yFFYizj+BzkuVgEFi598cFc+oBcJaP+djFthGl0kbLcui7A4kqXS/ajXvI0wFO6sjk9HPgonKli
Q5tOfgzeXGYo6Gns/dcu7mZJjYWp4F4VDW6SRo8z89eMJImMMNjUIvPnV057UPRlFSrkGihY8N0t
uJaHjZqwo+UES7zPkgNqerh+F7fNnYyL9m3Y0oliRYZgrTWd0AqVQpy7AfP1ju6XeAowYxPmwO7W
t67OCYwlEFhsVOLz0R/XCrwE6edFzTgEgYiiOP/h1Rv86O1sG9mXg4oVOBpNcLwiVJLQhs2kpom0
lnTPEX6OeqaA9o67p3/tQvuxbK4TStQLaDbnFyQcKaDD6ukzyrbUUwjYcks1yU+1MXqwItlAd4B3
yDwPW9YF6i0jA6ubCXglGQx/dWiWeGwVaJXEPAPVMV8WFysy3ScRGBZ2efqY262tHl0dwXT49zzN
sVtD6ekoeNr+AgYZAIT/FQjAN9JPo5ij0rTDgvdn2Icyd7lyXlMIyWEVc99r1rQjS8mgKbxDPeWt
IIT25zV2dVfgA17yaTsZWqSx8ztKg6AFOHNyKpkorCpBFyc24I3RFqcidww8dsEBOhkivEJ7FmEf
7wSLvWczY+lOd1lMrVrJ9DLNghRBsUivNTPJm9qNbdyQJ4YIicIf+CFfg2BTgQJKJLvQLXVytzCy
k9DIrdroGEUMjUmsaa63OJcZUK6zh//ch3DceBZiupTzaJNqEgSxLWQE7B+42mh99lcFmkEzG5J4
1qpm/X/yRhDKdoMaxrg4UMp6eAi+Zw+hQau8ckGuYS6oopcUq+lTRqHgQGfn584tEscEA6tQWVhR
P67ZJKT3yBAq5Edg8UykdDDfEeHdHqcIbbjd13AYkAsqbq7mZLMvqvzQTjivELrwALs+Ehte3lm8
QoFYptvrlInAhPxwgqpHZC4sa1ckcJ2JVtyjPADAaJRG0hvshEbdau2uoHY2vz1VsvqvICMfLEF2
YC1xUlV19ronP3xyHhxj/o2swFxGaSOeSZmp9INj/o/OU6EqmNYhgeazw1S/GyTDFojwunAJs1KK
5IZ6FVUh6DTmG3pnTUEZq4Olei4Hd/MyX05vDGQu9YKodk04siWoA9nOci5v6ElkmjsCF8OmKYCI
7nyWrhlz+7qOERiGJCAKK+67fCIJ7SE9UCbRG3+GmWQlgB/sNJJ304+R2Km1PHehQRykmlDtacD0
QPNFZwwKQf9cCNxae60X1M7Rxw3/b3CSZyDpEyuWjJxGYC8jT8hap363Auh+a1Q5Fc167irHWvU6
HsXwO30Odep0ht35K6xzC99OMccXWeBTRFVcaUf04JYbPnaP8dE/w1tOeV/dXgXgFspxSVBE6Djh
JjBX4lPW29EjWEpcrrCmny3l1UhfpSg7J4oT/nkoqxQ8B3e1QmrAsEsUCWsAeKiqYNtbMdjRAEgv
3tkCsO+vWKcsKUh0/tn/6HM1otzkBRLqVxoqsf4Twrap/ovn5jCScZA+TmgDKDti621jnDrotUJ7
wsCG+1canpib0wKcTDm29hWbLRqjlVe73XzpjxQLMf/crGmrAQWg0Tl+1QLA468hJT+qAeRHk2xt
LnbZa2apI1skdIBfNCzrc8gvW546OlRzlKCS4oZEFZ7ZG9xZi/bFF5sUR9xyzasYbq5PFMEpB7Fj
hYQg2Jlw6A/XGa7y3YVLHK0UGJFV9kdmbLnUbG1G9qyCRx5bl1tQfaz5Z1EzGhZP+xfpbxV8QpJD
EOXq29y3Tezprbcisldo27BVhPCpXT42JajtfCbaXMqWlR+8XwzwbZrHTq6vWnu/kx1Qpab2nBpU
a2V+iGsQREEZburaUA2f4Jxhr5YBxymWOa6UDdCxi7OyJG8aFq+xAZzZ/3N8SXUxem8nbahQYseT
vtgvo24e1Id88pV3cG+hW3BDa0SEFcP4Fa4sr9ZEGMKKlJdC11qxi1liTv5g1kgwXR7Dlh3uTxTy
U8pr6fRCO3UPl1Us+HRZYlREyUEmt3ulJILjMe1HPH5nsaFX54s4/zKZVUCEQE592XiUvdXa2Dk8
rQ0q6sqG+GjmeZNBtfpCyXj6sZlz7McLGaVzZd213aLOb51yMVMHdAfVUTZaB88aXp16pFUXsjqW
P8biKN6TkqLUPNBkDoDlgUa+KO5Ub7kF40MjGG3N/o+u3YV5wMUhVagAwbD9nMKW1QXVmGFawkIl
tlSVR0VL12dG6pDAL/FG9GpC3nkLitNT+2RHoKoot4A0kJx0yGeT8XRjEZkoTDnmtF/pCOc+azAo
HVRxXyx6KAmY6BsVjHQ7Pgw6WoxpN+TkF0gfg/1ojztDIctUSq/pHL0M1nyf4bLP9z2SJAF2MGTX
Rq41uwoz00QKNh5dpI+8Lq9gNCChRjOXPqe96MEhL/bwdb/vU6U1az14jsRRSduMwVyjlT0LowVL
G2C+xAL7j7GUn2omPEddSvvWimW9f/Lm+oxqCLG1U52aVQp8AQm1p5Rp1e6BmN32k/4Prf6uFSia
1x0L/uPYGQvQ0uPLbFDN4UUFXmZqg6UMXP/Jar/3fKVSejA+Q5eIJ2zEsCRa3lKCLz+Ip6UK5b9q
KVmHSuwWdYvg9YbP2ZT2JOC6qwQLyHSneYFTUzGYsZqMB7ayKmgjuLejAE0Ug6dAu4XCWMFu/IsY
xhNZDA4En6EZU4D6X76ddwQrpjcFgpdJ2glvcdWNsgpFrEMOPhagkvhdaRmrAIFyJzjh3COVBmFJ
Aspyb8m4BnJlrDpFFuqtLpGwNXIs2Kta20aVUxxuIX2mk0dhXqjU3FnMyhFzapn2nSfPAPp4pTSP
9faJogwmoOqLyqfb3iWVOPGJeJGcJvjJBaZxclYZoLksaLu6bZrpzucQBmlPmFwuQMRp6n/Czuor
rd8QW4uKWaUr+Oy6zwH2cAVYlumJhwRikPj9UXkgrl0M0qRtytKTnOsj9jBnI4zMvnrSWP7ZYG+J
gktCyb95t9Bv+nPDH/7bYWZ+eMiwOLrWKiZkDT7UyPNH36TmFXanNA2ubEtfqSw5NA1spQM+rxQ/
aTOMfg6iuYj3TUWaPfV1Ggd7cjg5ZExFgNoE30fjIXqsbq19MUKOdcMVJemVTvTWoZP1EbOaNSIC
H3AKUc5/osrFEyV3mRnNV4nGX8Tz3/NH50bkRAgOJbZ6r/QYe8Irp1sKgY8aY/DAulIiXwJlmaED
QnqBMJQaze3BlGVUwBA81TGxf1UfuSoSmZLqLh7gXE8csOhFG8rxXtu8Vi+Q9NttH1l+QAONqbHv
fCKLH1mrOKEMbZHl/UDCd64SnZZ953jjo1uSMUwHVPKevEsWSZd9pQKfkmUAIAsbJYNKt1rf/TgM
x69rT3KOvm1Hu/kASuF82V48pm2D7GuJ3CHvHeahp2f2niZKSVg3YB5Z4QSSeQR164rMsRZgdst6
uXU256N40+aw2Li1AAC+OZv0pxnzcIZn7f5roegnaUlxg6gUqshy+Oyjfi2hqZwsGz5YyZT/uGkh
IB8M0RSFcz3VfWM38iNsWsqTHiFbASJ0peM3lR9UnIaEUPJtwo7Pqe+hBt1XFgkmOz3qp3gu4+5h
G1x0AEh5SmOEjQWp0u2M/s/aVSJWhwSa+yabASV9Mz9TfznRqpebh2EUZnSLTGpHnZaaxFoSPLGv
mIpw5P8R7XtzxBaA73h1rJo6zZ8gGFRpMNygYZmLc9kaOgglHM7x0+Yg1YpxFmd5pSEjSMxCy1yz
B0GrblBa5/uWqyQgfdjBFxNd0mU54SR/t0W6ulPP1yCxJqMNhtSP76t6cTKtl8RQb8JNADvDffka
/0GOW0jTzXXmHzqwXo2OQhQzN4sQvea6Q69+rggqisOcRlJY1pMPWy0XlemVupD+mPAbfKyM9PdW
Tk7qFMDcvACSZcHT2tr6gVUT6TCab/59BnRjmSLA3yI0aZU/rHstzjgwJ33aCz6c3RVJH+wxZPr5
AH5R0A2+jWN57fxmyhzVaMr7FLrc3fqov2TrhSM/NTSpimmYymI6Le3GJmWP3mSZvZQhcOoZYM1n
1+DBU/Cqcf9i7JnTfEPQpMqMzWuASYYA2fWD5xY+Fmkt9BBAWScikvZs/lgwlvCEaK+8DVFpW7JK
/anAF800tmkCgVeeX1yGR1ndds/AmViMeq1pDqL18UuVZlR9WJDCZ61jlxLf589eBCxAGRMXmGoO
tGxkz9O/ioJQakTPzEF4p7mUh69mnRkdmdtoVOI100zqmu1PP/I/mWfcZJKJWyNXaretJPddEsbq
Rtv0YVpBh8E8DMiqvsXiNk4EFTqsRFcv5ghsPGiPPemHBCizJz0+3KosLIn4poSkstbR92UIbLKS
hCWv58vZ7nFuilBKqiL5+MkMOJm0rOR5I6KI1JO2IxA//PuSWvsVwrI4iNr+29VinJrBLbqNUu9+
wM6QaM/0JL+gbC2SK8qofdd8D2czL1g73oPoKtx/+EX29/QVJASRa3Wow7PaH8J4mJ89T2c+9BZj
VCv1lv6j0ZnK0y2LdZ7l4XR43hrTdwcDzgjgl4f2GT9NwtQ/zqYKm2VQatgAHjV6A1Nmng+WuUH4
3Ub5Wgenfs/iq/MJ3cSJ/T0tQvLZp9LUWKusrZZJ6yOyRVa1xX+N4/NvcmnQ8CkDmhYKhGb4vy7M
NB/BIJ5FbL0RcxzvHoswu9TD9N+IDMkYDSqVo5ls0ALYNexGXGartEijjSCmlg9KB3LkMXkS1Es4
p3dESwu87zrA9/d4RWrH/E/fgSwxz6BKu2l99rg/3CpZeIrDSm22jKgo4SuKshBj8XBN1ZXhbaxE
EgQ/vjGStaF3whdX+Z8M0iq3ZixW9MO0cfrNJk+nZGuYHlvWmAbyK+TR6pWkROTLBOX2zUgggdJr
APQ7z/Sv+nVUKPpfw6WIi/rjEgyTZioZ4WvrcJjlfj6YzuD4gpwSIfCQ69/V/kETNGoZkN7/5fuj
KQ0IKvHMjwP9cm0qixHH3AnOYGeOjGG36/19/kd/pBeWsHBC5FD1tGBvDjUqDwGWEiMishYHKWlG
lPkby9cD8WOYvRXpmRaoVm3CgEHm5bM0Mx9bvHKMHsXrBfX7HRJIJ4Im9A3rAe/zabVD5z8hVF/y
k8u27Gwn4gz5z5VpRvtrSQ/K16dwPtzgVGtgNG4j5Y0TtOTH9Inj/n6zb26ItJvWtO6B2SWKkTW7
5leJ85kLRia7vHdpqE7Oitm/jNyhhPi/nJG6/8B8ZvKDxT96MwnoL8BR6UtBQeC/0gL6+5qwwIAb
xVSMKfqCAJX//YgxWd/LsrYGJbA/r9tFyyIemygTSj0dcb4bngjlxpPAfI9UmHKfUs+1nKigHjvY
yhAkSi7Drzi2bgEpNPXgIKuorfJaMAHCE1hBs9kFbrIwJidJo3MFUoAXTZZL4OqOdTvzhvltwsz5
0O+KeHoGMEgJMllpo+lsCwMMcW5wIWKXhow5Ui9hjXBM1IgXjWBzBxWFSGkHsTCDrRm3oPyMjmIY
lhHcBOjrlm7eu4MMAPZHb5TEyo5E+ddwJZsMv9dOMVuAnsRJhKKyFM0WVd52etdTyEOopnE12mft
d9SJbSNIC/HNOSgMKlxTdMh1nOHRl4KZQdHgKTMjRTGou2/09tXBozqDBs1sAFS6JyHM/dXGzYQ3
EavTck5EV042aFU4sKIYpAu00jslo3MTejU/V4PK74XfkNWSni5BQcNB6lhP4GO8mnFDcO46mHOi
d02LlNwHSFB6bPLaq+rxmsjqjFLars3fy0MNuC/B4Wey7urRlPwcrySWWm/hQ29nGpiHmgz1yOGh
/Dgb7v4TMhHds5XtEVo9O0XqHOrWk5Qp0XXOimm9hikYqEVMiHd5jVrd3igzIituyELGiYjrw6i0
+P5VZwvBTTbU9GiKhg4D48gAONua1AOiR2Ber98/hbS7mOy0zF81JQctdKEdOdU4FMSg9WMRuCPF
VbdjFsCvOwebzhOpPjxUcO8NJgqkcenFVPCBdq/5s/wBtkKgfTdgDwpDIK1XAQ8CdOsyobtV9Wt+
LZo99SX6DxPu4Y8JAMFqryzGCsqToJIQ7bslfaQ06tbfKJW4vnwRq9WIH/RBwcZpzfnMbmMh5DA4
7OZgFzOs9Wb8YSBPtzeVuF+gqu3uR7dcN/FqtuIOYYhfPdDPN10E9ofGy/zzXjYrsTcm3d3m3b9q
mWEG6d0/MWZMCqMZayZk+S81sDJwIRr6hJAeVLmeiFUiFz+YIE08ToMkXARv78mclqGz3i0EFhvI
7jg2T8PYF643iplp4JEwC8EBtV7AyuYNvpNXurgAXc/L+vDxeBrfUNl5ZPtBwN3c+w9co6t7+j5s
H+/Wo8WZqUQvUh9r9qJc2neDe0PLm/6eceutHCaKaATNJatZQaqAM5cXWoxJYIaZiNyssgF502rA
f6gXOpFdDgyKjOFi8d5C2zVyVS4O2QvXoAPIurNDV5JQrd9IKjn3GNghTBIuI9FrhmMXq0NQDr5M
VdAdPFQW74+RhKBAktbNG7ItN2qMQoV5CRnQXcec8ZQANcB5S4S/2Fe91iFTmzVCofbSvOOOxR69
QIBcyRGlHE5Q7DL5oiu6rc/e9LRNAmT7AaEDE5s/PW//5mTKA83oV0ksVsXuldOqmoq04VxIXhaj
8TkI27XGe4QGQ7iYxrvr+tG79kn2sPw/HsseNeTHHIZAXQvR0v49w8He23FsPPYi64bUyuKFvyiJ
pbeVxwPZOz8VIwKH4aMTLJ/TDJFKfn6rRK/PjY8Z0e7l7CYn5/7mCebFBXIxJ9orXGFk5Nj+Do+w
q3NBSnXfG9MpP/lp6a5kWJS3n0YzgjP2Bk5HbfzX6qDO+BQ7aaWts5PqQbomPiI5RxFsLesPTsEj
TpjPcPRcUHpN5si9gxvC9aJZfZvyQLX51+kGkWv5n891H3aidSru5kzNZl7+dHI/prLMIGGCW7Ho
/eEz6HxUZCy74qK64/yJJS8lieAe6Y/kfpIYjhT8c+ZQp/hhcLliy6ZsqFxDv235Qvh/xJ2R4E+I
GmwpNikxYDBcET53SJSSU575E/U9UOi82ZgbHActvm8xIVAXnkrDwlI+VrQB3RB6fRYcfQB83k+b
7+Du9WGQIO8IpUuRHobYGQT0m2O7hYrPH9wYmMKRYCYaOAadRQenUnuS23NfnUuHRYAbxMScx/GG
MAf5F0y6u7sEZIqHEBy8Dz41BxBmbMTKW9BXRcZPH2WlmfQo+6Vd8uEsATAE7j/72j8xJ5AAzba1
Svvgxm79v29IGekkpdVdBqshxhv7wJTdC6GNM1k/u/meIXzdZLZsYRiDv+kcNhd/Mkdsf5+lMQdW
2AY2RdXxFqIKb6UdjCMtMt/lGehQ2cEIpyIEJB5OnK/ySmadvqhZWkgF1kKU+spkWqbz7bBFFZ0S
rAfK6dMp9/4ClhZqmR6qJnxmc9S4FX+CPTzQcGgNdyrHDawrvMhw55LJ9SetAeWVKQ9MVrlA/x7c
AYUQets2QTAlUe3m5fh67yRAmzH77+SSL98coIn67WC4YK4al0Bg+JelUFYI7Jjq0HscPLzOIHHS
BDhLFB5+EOBZt9YzLc0rlUPQimao2NEMmzVLpfnhZJ24/ZOYqJzTRGqXUj4d+Eh+FTliuTBYIHSh
km0LcTWU05iolVn6iI0ocVtWIWZe9bevYttDLpifGEUTaxoqvFPeWcjE0Krpxm435j2ScHuopGu2
l3LIVZuIl+0HmbF+cQd7ui7PC8E8kmKYNJABZzsTSKCCl2dWf7P0OAl/F/Illd3LxPqTf76Sq974
EqzQjO4BRRdrv58JKBhYVntK/Y5OuAi98FKaYHVwpsnz07x/9oqNHyGGxnvAEwKb6BSKFpEznaMh
lGZ/TMQvtM4KOasLEtdGxGZnYpv2+QlznxzVuIiMeicD+17Z9o9g9grAMHoDdjy8dbkTZU/Jy2wZ
ThzJu/9X3s8TMg2WWm4EJW70Ju+4ETWrPEu9ZggRLQ51xGendPnljTMrwlHavpXYyvP57lvDUgPb
rquDD9Usg9rFvEyThUcwAGrxSPSfWUQ60Am+ls42qvpdbqWEWmTkLuFKFMUpX7bpCuilYk+dixZl
hrYtXCP2PxqSqAnieKHhFvbdJoWt0NTbXUqJnuJFzwRMEwnKJWgJLsPo76a4VwXlY6mCA8ZMsx53
R99BGYsWAQ+gOOTG4mBrc+8xUL00N+hfn/ulvooSzYG9HmchjS2oJf1/hb3DPwI1zOD43hACYThi
t4iEQ2hzTuru+74KwUdDqr04o5cDbrmo3jUSDCCc79FNnbGqcQnODwHSafOMwAkabBvKtwhhyilf
sWFOaqCBV6lrm3tODYuUOjTWlJnGumC0eKpBqevEEehg7n8OgCWoqJ2DMpBCp/v9h8sNDFKgWZrt
iVpQG4k8xeeQtPFwuhk6vMPnknvXNa1rxaas9/L3JEaiXk6XarcfLdln2WVhbLbZ695q1BxGDOir
HLQMD1OyWVTVSRU52OFiBevIira1iwnyClmHj5T39J6QDrEtWjeuZRjdTdxEl8J1v4IVK0CVCtEx
FmZ6lbLLyZTsDvJuKYeSBcNMWKJ7McwbVk25H5CzvK67kRjEp+ZKuj86MpMXxASShBQSgHw3sdnM
T4BhNA65ovKTHkSzzFr9rtbzqC29B9Y9TcqypGpb67cLDqH3jveljaBItOCqdMjV4DxU4q2K4afw
Tm8zfrTQM/Qul0apy4PhmAMkr7VFZXSFtoPXuaX1zjcmFWmkXvKT6D3bAIe/3kIRvEE978/9pDuU
GGO6GykgCT3bYHKP4bfOH9mn+EMpRT1bkmRWiFd8n6rt5A20ukztUsi40zjEHhlIAVKdJz2cpV4t
h8j1ie5V8PyZSqXWOuP94tSYzDAQ/l8etVjdz+Hp6ALaSUf+gGMDhB0Hm3pdFsOQ4jKKjP88Q9da
hpWkGiHBeB+MyMLoLaNGw0XsbgTR3vHSd8l8qqxbYAUZNNO51kHqINR5nWfOU4AyRtNLZ9XsO/hF
TENIU2Vu9dl0sV8NQzxXlLDf1Wao6GoJdr2GjtT2miiMBcO3wqyGNBx8nYQcolqG+OOVa+fEC+eG
FEuog/8iMXKKFwn9d3m4eUNGAqRDK+inXS0uDODgHnNQEmq//V50DqH599gEUT/fJyD6on3W3hRg
DCzoDYNHwqizzfwb/8/U6e6XyS5YXj7pdGEx4azgnrWsW+3lA9JcxGQvOWmok5rZfbBH5wn0HGht
gAhz/Zy30iuYn7FiLFVWYuB0U1lnML+LMsyEnZf7zrm7odKEMg2RbRMbPB6LFbbFrUc8zO4/SGbZ
uVfsb8Ejs6wq1gtOmTEANuMX1e9yv0t6F6eEg/BUSG7JW16djmv0rlOMVCDaPJ4wv5tSEHJmkG8r
xQpWsYeiap4vrzq9kFg0FXR4Luyy1wKujhj1oOk9ykPr5lFML1ybgQjqTpTV9m4G/dR8ZgjUV8hM
PR95phrgF25Da97LQKNASewShZFBRGw1oL7wgK4zXSZsTwO/pOsWWHjygvL2Dp0ZB7RVntgmBxZB
SCRuMOxN79eAKsHNa5s8O0RY9Zp8ONXAxvBuJ+vJNjSEaoRVsRZ8VJtphJLhUm6gZZHDZ37J6oMX
Sio01/DzIy5btlNr+VdG3LGLAz6Ulu6Ffw1ppu+vJjFQZtiBCEn5NGHWxyc3BHSmgurJosnwe9kb
27BnmLE0Gz0YEnwEhkvlu9JYCKvYLSf+c6WeHrTXspkuEBv71swC43rZVai4SPE4aQz3ZAXe2sCp
vZN2FUZb34kMAWw1zcb9TvCLYc5BM0zRDyqzfWFI1N2sTwUYmJ2CzqQE3Z4HYYDVpyLsgT3GncmP
AOE8wEJ/9tpNoWVhZuCHFf0woXousG0aZt2AUq1OHVFu6DLBShpy5OMAievW/4VCKtcH65suHF5G
4hHeBUa9ARLYtPBZNgpqvWLRFzc/r3s9vlx1XT+cTq2RvnMpCZNnn5aGCik8Js//t31thz7dwUse
r/Lj+iMnBvk4/topvHDwEKpXt+5Nx7ByIz4p4gkMeaoxlRB2tqIsFEVWU3ypN13gAnJpSchktiRF
hIGwAVfe2FUZjnpMBPISqutSmeWV5dGBv7QD7XyATVmvjJD2z9IXUUsa0dyMkDi5ZXMvMl3EN3en
qiStLT+Pd//KRo26iM+qUZ+OdD2PeQC9elEvYMgMmEkglwWcsdrv3+VwUlgafT7UlhN480Y74Ser
/jsGpk79PBrbOgDDsZfhV6kLKREhSfEvmY7p9PAmSK6N+noBbNaApZi/DZ1d+5tXldNkblJX37nb
MeHq6+z5FwbzGbSaLgegdL/SSMJisWTJF+w91pgh+7J+Jg+gcwN2F1hBThwzRVbEPXLF0rbcqg1V
tcrJhz+lbAWzfxmLNLMH8jcnA7/en77XTao5u+NdGhjzG4TbFoTRydTH13EIjE14xNnmoqNW9J5l
Pza6Z2WAOktsFDWF9yovMRkiU197VU8RZuU1NmcFRhyUO9Mz8bv6i8vPSh+NlGUVvIaKayB4MZhU
PPS4amsW1gc5wfYN1l9PWTqApQ6yDfG7FyJhVf+wZ33SBv9Ecg/8ITFtB6Xzj2lBwxzK64DM8RPP
v9Bs5hRy5u/afWj4nLR7u0OMb7R/uoiyKZgZcqoPMJeFh8fbfanExmPMwWrs3b94Z3L3LiIET5Xw
B6N2JHoK8ATmGwq44krUsZl0DbVk6ptdKQrwR0w6Vn9maGA9sE8PJrbyptZGdWUFTIDSqaMTO4CC
KW+QQJ/r70cN5F67t+vDw9nX6Sn/1a8qFhXISscifJVSLEOCK/6uGVdzWGC0Qhqa7ig283JwsfRk
7b43CHILbmW+2+MpcqO3hhtQfH46ytN7GixbJ4qI9doTI/VF6Br32gjdMo8D41c2t3gRc+FgufMJ
zN42PZrJ5TGF8qJre37coT9H9OMqPLAPtj2s9Gh3eYH49Fc1neXjJ09Euu8m4U1l1EVTktxZTeye
iZEDP9IlAnqBC1lZJzgPd31kA1sPM036V06qlogHbI3cDSGtAyxgEmhRJE9/hKzr5DSmo9fIrSiS
1LMxVwkNR748uPNBrTg4o+fwQwgt2lz2cnQSjfTOHM6zGfmrgh/Hps3Nz1qydxpuSqJNwcrFiMSI
HpHRNRYi8e4aAnJgh7MdW6LR4PeEGTlq7FQqUYzZjEqHSUrzdLxdnPT2EtzxLA+22/HtwIv7f6vW
VifE8xgmcrEfk6qqvzsQ+gn4RyntynUhQAiG0CDgeWtRjBV0nyH+ng0iviMeB+B8/yxOl1/hlKYK
Njtxvin8wf88SMt4ZBJ0MYNxkKNGYpROFif2G2N4MlPYUvwWQQdo+AS3uKkrILMSjkwYNcRdnWHs
dkgkcyGPD3cWY09ix7TUthi1dCeFqwZ15v6xXwS4vABasEoCniIZ/qUWHWEYhg09DHe53HIShnA2
Ue1skek6XFeXK+OkBIoYdmllwwWhti7uofSdFbHIJ8dj7cU0BGQGSTg8We07BsfU14Z+Tsn5oKU8
5+9Gc2WmvNfmhCZ6bIb54gb35DZRH9bWU38QGTB26yEarud/bgOj4KaGv2uekEZjxLTv2Nnpy4oB
7OaBRnJb5Ap4dHsCGONjkkjDJEbZ1033cCRWKXa81L31avjTuBnrK7A/0pEveSD7uBOF/X4ZM9UD
IFsYtBmSLMxPtmE/Q9ULT23X//I63e+PMRqhMj99WQioAKdl0TvcIWh9E4HRPXYjzYL4/IAL3arP
lQUa/Z8ONNa8oSzlxU0PJYzH5i/5u6tzQanhlnsuKRnSgzRpi/1GWSl/gn+6G3zhkwJtv80Owhtx
m4zobzgd1wX7JHoVFvtV8UXA/BHAUJDhiqS1h8UC6evsFDDmvX8KVkLfjHbAW20hPZl34uVgsU4V
Z61xmMtuepncBPy/oyJDd9DUXwStqd5WnlwrQWq1zPAQEGvdZ08crwr0D4YYStN7a/Gzg69XcYp7
oghFd/v4w7VSd6vxLe2J81kK3RQJ0+mj6nMf7lsxnYpf51Z20aGaF+nIHbtun4/OFlEZQn6Gqe55
kQMvOgU5kelmfdjX1e766dxWk13+zZOpvxDU/eWP+yRqs/1YNFrV2KvW4YXTkWBACujuwJMpy0Li
WdiVzKy9j7Iu18CRud+/71Y5cZ+LaxSftLPn6kedXj5XRA9fCjDbFyZRgMa/s1cf22qxOE+jACHX
YhcWRMW7yeZLfAsDSKmYBdWTQp6EjOhqjKfQwnzv2fSckJ30cJmZt++o2NRAJdP7f2nnGUaQx3sS
vKgtHGuPpVVz3o9EA+DbzXwzPl38pQs1ypkLDPXyFjtmieZRpEX04N5pGxpWaC7w9OLtExXsOZQn
W5EsclbWL6QyGAOHojl7R9KE4tKi6x2MMqAHaY6VEV21biqrmJbCuPmcXvz1GPwFqjnqpJAolQNg
WSEnKEo4EP9YnDArYEu+CfFzrGsGoe8kqBjX0zfCJ/wj2DPJTq5KXW1e9+mCs/CmtrqyYV20OZto
p76FVPnCSskuu2pSzqe1Ap+VQza9rbIr58Lj3scEySavxumYKZBmEGAgAU3zV3P5QzajWsEWw28L
WcXimpQNpmnxbsEhFlTQi7JXnbcHCff24K2KKBol+7fBTFBwIdmQHtrEe2gbeQQQw82Q3KDKDPQM
uV/ZzJSdPtvWsNNgpmXyB1EhocvPMS9krshUfYL3AxcSbkleW4LTQUtT5t1zerofpbOSl/BMWxbC
B0F1Rzh98p5/RGpiwIanYrvi/aITdwWt3aPyOSKyTnA2Ne7SO6w1ayh+pZ5av1dOG9gMo7c/Q0QZ
XxLQEMt6DX/NlyfKTnqONixyYkaX31IXSv+uG+opNtuGwdwStSSdbHU7U3zchO2hMYzOap9At+p4
0mQSMpKNjzokztjao63t4vNBVnIUnte/uND2V3joBwQT9appEqBVJ929Hy6tJXWvvpZ8sPOUxFEa
ioX0YVtU55963McSYXC/DnatYRq4wBYUq217rgSd02OjrZbZ9y23PgFgxHxY4IuL2PogqZIotnWa
vhweTBPZQhdWif3HfWd4ojoQe7fw4fcWQPmvPTB8JXmsxfSS8TAnHF55WVd3bBH5rCg1H0UZV9FL
2+1M+Dqo5YXp/ezoEW6J0AzGeUQ6KQvNIQ5dHQo/sE5IgaFFeABcFCSCE6px74J14W+yv6HKhg66
W3jyw5i4PCg4DF3ieWYYrg/tXXrD8ZsfB1ybeWddD4Ea38l6FoRvCue6UUMKd16ekkZJIERMMUMj
qtFCUgyuz1VfSyu7Sj5Lg3t1KWw5mLc1X1XFJbTlX3NowS+xbd2H0xHKVAtZizwaumO6nmxvWPlg
NQgP8xgcOzDwwxqRL5kMrDeVw4OvJmVIaVaASMlLUMjL08s0ykZrsSqkfRmA/4EP49stoPyQyz1A
hNVHhySXJ2w6LXXmq3KRF795udB8cohx7SqysQoYz22gzmM54UBdCeXQGDn3LmAt19S7UT3g5rth
StbnuhjT+Jp5QRd+VvrxF03+6m6MN/HATpaZmvcYiAaTNaTo6Bb2JMhr5Y/usz6Z83W+BYmTIUNV
4W7+T1b1ol2T4jGQ2ZVUgOKxBVTCc9NhGH3tHGEc0m2YOFaPTUlVySuft8GaKbQF65mLyZHTOFha
MaY4ftTuxAHU1c+vdrQnBjyLfkdcwxX6iDcSBy8agM4KD07PydJPVH7QFA90kUXOYAQoIBSkZLw2
J3ORVIUzaNSQ5CVhAKDXEe7cNG4bxfjdyo58N2MY5ypgidmeHEME5FQhTIE7waodBU/f1WkPFojC
cCizaiZGkYLvCQ05wwYB7/DNwO/FODhHZjcz5jAFGZdkxMguaTaszGEYe6JpM9/GpVCI+UnRcidd
gUKUULJqz6AtAkxtaMucxL/Zz5pYsp36mP4V+7f/Vvi4w6GYR/1uTdh413Gz4mqbpyod01pQzFGX
RYV1f9R5ecDxDTZ/p5Ko1780o2gtXsKOBZz3qbUrJAozVc9rjviJBEfrgemyIjqTXAzsXWIVhxpL
/hnVo3rXwtXNtf6ZfFyxfU747uAmDetK/ezShlio2f6KacadWSk242fxeMQG3WmgnY3885IVerId
geizuI4WVLfA+9Haww8WjtRsBFJw4pZPBPVbohnNL47/2uMxs9bZHb6rwhyTE/x6R/JXphnLbSgX
/LMuCS5q/t5rCvFVR/wuD+a8HnwBPgYh4atZx9g75EVwx6Ze1B42Bh5FmI1GYEQd4Vk5h6J9zCdi
KogcSMvOiU0A3YqaadndV8Mc9awk60IVvV2F77AnIEw/UW8DhP7u48b8wPNBGFlqOQDLZHJMHnNw
hBfySjGMuHdo1G1+5Qryf76X94xPb2Z0ACuxORUIv2Lx1LMxz5tcS0vaav0aZ8mKpxii6vUQl658
teBpd50LGXLOAnpdJP5I+9dwmmtGeueLxDFLSP0pgUCy8O0ACt0qkNV6EU0djOziiTjAIQZArMYn
w6VQkOFJUMowLC63W/NqZ7TtFeClj3clr1TLC2kQvKOJY6/27D/VN/lDhdjvX40+HNBbWhhXqMbe
pt/7titPd2VAtcynR0boNgP+daql853af2n0Vhb8q2IOLFjxAemLmMZZUgP+zqRACJp1zRhbHaT/
Fmq3qJ+Vn1+FeAPPzFoRtRZJPiB4lfDaFaxZXpdQjcD3y1DLuY6Z7c7lbOnaRk40So6tzC7Yn1FQ
zVtpDGQS0qi+khp5yaAyAqhtuv+sOJT86Nr32n8+gtuSAlCUkTcq86mYSq0fjYsXvXxhHDyTETSD
FEs1libT6+rMZ/Jw5boLvPYG3CSEPgBR6B0uuoNUiFM/cnGATsL3lsKI8KQnEiHwF5iCdez6T3kd
74F4Rlvjb+EZOEeewpUGIo/5T864q6h4mWugEgpM1k1hqojAle8WAharU5QyPTgUH3Fe6Cp3N2Ua
pwiQOM0fRFD8i2TrqLwJpgwx2bZ4WSz+LZafu/ERf0od5hvZbU8asumxBAHdGMeDEsKcW9DwPlUY
uw3RJkGkdQ5om3XeYnoV0EYtQEK6y0zUvmLC3uZ9hr/MZpH12UZiTCN99d30X3etQtz5PEyEVtRH
dUG/kbwupXFZUaO/0AD3JhmWI/d+yk7ZeFkZtG5P9nRZ2H1o7jE8LIsfIp8e3Yz2WzYDAIraWUwH
Iq6cdjdX/aUvh9xUWQPpx3EM0qDR8haJcal3M8gxjqAPUvF1plXzRl8BjYzhaWJkSbveg3YdKAKJ
NCSYOMiEaxD50GFWZji2LNsWi4fJYEpg+9w3jMlwSfjolixJA0tvvRymDGGBXvBGN7DGqoYEsctf
PBwQaUyhMQYiJWqEKru9M3C4B2kd7IHhny+zuhNE8KxoBvVbQE4BFVba+isTG8kDVbRBHfIqhQWt
pRvGheoclliypA5jFPWEoX5wCM7AeEPSvW8KhbtDih6xlzEuFMdn/iZcePkIMI/1OgZBG/VXSF4g
l8svbz6BKRtpw/nRFUDdhgjRoq/t23zzFFvYvb1F9e3tAkybbV+LOGreOPD/ForaVXGruCxg7O1D
N47HLyKJBR05JeJ0EbaTuJH7KUy8TkPaU+zTUceGsMUemGAeftKDf6ZuNI3j0xSiUZBSUlReDdOh
ivDXwpLxPd+irR+stUhIJLCZD1GfmPZRBId5fqzvmwRCQ+J0HLbSLidVK0cVFlmjxkKmdFqaRZBi
Xy8wogaMczbJmumZtl4MN4G0nIbPD1HFVqESU8fL9KbYtRjd7IHIbGSBBgxlVKYBvBjI9ERBP/tM
gVWvU4hVCS+v91FlQEdLjWqkgin5+mp0rcUQuZI7X5PPLZEjzgJU/hKqioeH3/uz00f/3II2L15q
db5+yZVY1dljJnhhB2rPil9xpJdrOdGJMrOImgl/jhu4J/NiIhca4MzMvkNbjYBav3T9WmoNV7ml
XJugcXCrNJnjifoZG6Pv8Kl4vYerBst4iqRgAtNPTLSpda779PRU0r8qVvcv4alfyOj1wRv+NHJd
3oPSJ3z13z5ij6KSvCBUeYrNrRez5Jmf0XzmqqE8tUgKYj5uHZ0w5ddKV16Bxdmf4NpXEAOC9Ajw
PR6IFqUUstVONyXylu55letmSRipnj4Vn4tfg9EjddY2ijgE+3DIIz7OAZcoEFemPD0hbSx2TAgP
dvDt9wr3kRAC8Wh5ToOmEiwuX85AcKfe8yNXAcIGhhf+X2ANtCUi8Dq8iS8mDmkNqZRpBwGTyEH7
aPZv7NHJV7xCV//8IoDTDBUfS5X3vgfs1CcaVrP3EE/VFi17v5TUqc18W7to8cVr4IzM5vgxNpJH
UIzdMW9dM/WuHsN0LRhJvnOm9HbTdcStlZms8ZWROOZKXZoEb7wtD3vTtDOQPFiW8L20fsS1pWRp
a4WQf4FkJKal+zrDcOwt1uaZ2gIsT50n37/X2wNeISlM989oLa99FtlzFyrKvmUGB9GSHiFrzES2
iQdGs3hV2SwBIxqK1QM2JyaFlgoQvh7YcwHmnrFzNlkh8vckswm722og1Wc/bUN/NxHJ55W2Evez
QJrcMeM8eJQCSYkygpBFCnb6dXBSU8bCP8CheD3Mfxj91iqzFeRzWDez5bwCUOE69u2LhO3uwQv7
kCG6ZFfiq7bOKroX77O2wS4LQOP5ZzuRa1O2IWKkgn5WjGtLVZ5Ozss3CzQ3EYVkQRM5XKXP5YhS
JxH+KiBSIG/KapMlIfkQ0CWe6qX0XhJQwJuhs3RCBCO426iY2oDRqVs82+i9RtZGVEk1vU3Xo4XX
5UzvUg4xIq/sEwVnY1yaApxAkO0D3mKXzNDNQgaWJtU3qJe9gyZmC2wcxynlc+Btw3UZVxtk9/G5
laMv8j/MPcul7E/+xi1ptORoduY/uLsQoNHtgCuIq1ofRlQgXBIAUaw3cYb8WIJuMmOXI+OpDj0R
VV2hnRCa/IoQH3l/AzZMFnjkgr4BzrbcG0SKlxUkJxXaC20wZvy344BoYZU/rMDsRVjbn7Ff41us
wcrGzrYS1bYUOWC8XzuGummecfbRIBrE+qouVxdsLgrRJWsRprbc3+pL6xci79+gI4cVZ3/gn4yq
vRuSRmwUQV5dBZZdMXpWHbrps/3VUUnqGbbkcyoR7a38/fNZOBTBCvgWpaR6dWvZFd/P9In2fmmz
z4be8C7ttFvEuXozhJbNObFEdRq3Q5dK/qUfGWXIGQhaM0M6S2E4gcAgzHAyICOWXdjAnTJEFhEC
NJxcfe+twWJ3U8ch0FT7ZeS3qa0zAc3N337O6ji2oO894btgy/JJ44SAgMioDu2atk+a71LbxDdP
I2imDEQFZ5exy/C6Qttld3k7wn/LNk9UnRVn3Lim8T6/UKcDeRzRbvvRoAQ0EPm8tGFI7cHw8jzA
sM5oiP1gBH7RN6ax3f+sqFRfC1/q2tX4u6ho10yDjmuvEvA5D2eoOSDn4AmZ6Hrxp/FMRCLS+v1c
IdCOliuI6vey4JPuLEU6n0HcF12M1hi3Te8qqgwvPOGwjFSi943ko93OxFlyjY7yqW7+2dBRzyg7
JT0rim7Z4wMEiqon3olU2BCbrMDgq2JyvOlkHV2cJRTMKnu6SgYkloQQ6Ehosznp2x0GMHCygrkJ
mYS5YCxsAg6CvTkUd5UCbPbcCLxyWDtSGc3C7mpOgmksho/2zZPxLzT/6i0By3ITsP90xURQ9iMd
BTZFiIZCq/K6Mily1aKewKiBI+nEIjhQkUTW7hfqta22UPk3Fhu38GPypot7ZewiT4odpNuQ2TEk
K0+ytK35e4JaB3ffqZiNxz7MJw3Qbg6INjXJjxTw3E0HS4O+V+ENcAWh2b/bRkLrk1xwZdTMM55O
gz6bydC99HY4GfWaTuQbMKZc7lZ6eFf1TRqd87+ZLJz+hUvpYQDh7QCYISeEPesZxdgFqrGxe3gL
k0bWb0FVgIPkwzjnrtaQ7vmwrh27RQZ8NMTvQOgluDSjKB4TLxtFLYIgQY6MqZOdo8helXs6x/H+
y3A9FAxzwpRZ7vB+hzkYrhF7f1ixdG4FZCzJBQ39E/d5S5B7Yh6XPYOmxXpk0YRUzNAsDkW2C+cm
OC3GyuELDZnnEBce1g7kTyGkFlKkjhB+kGJZ69ANhhFwq8w2AEy4ulZG9mJ7RPw7SD4NV6BaWY0Y
nh6OyS6uRrujhEfm90Eo3iSL1QT8YldDl3ypY8JF2kpkYM/9hwPzIU5YLklNFR/6opdVI+HqykMG
Q4h3emd2QxTln2YO1WzEqfs42Ctx9Gtq0HUq607Oy1INnbWfEA9ceItEjjDG+zDSmAamWtI89EL8
p0TCuxl2m7XCLFc0r316N09w11QkaEBI+cH7287Gh/ZusDqS3p4v0yZqcsofsnYnyqLE4c3Yei47
9ZAJv0xcvv21zbMUO5MPbhJxwgAOkgRDrUodyetns45yxMuC5RSY/ymHSm8hCbx0JKA8fyif/4j5
liJrNaDvfy5UjYPExdQ+larig9tHldj7m1kemrZex8dWQ09APxQFlau+jS3tJa2K+JL5KUwZbcrw
hkQ+f3uFWYfO/3jifaly/ifpMZATA+yHbNTWKQ3VSRrc5XEPrYtFq8wxUsxMuZ206/Fj9O9vemMz
0mFQui/x6Jmz0Z1uUO/t/s97Z2LMYJx2uic0NNuO/wwIGd7yecdqVkEBa9jdF7g5jFP3IcB1SRi0
hG84KhbpMlLLCwG6/0kksXbVzkPFIGJCWSR8tojyDGGs2Crit9V6/tj5W4/6l+3rfJdlzlINoyZv
yjIHTdhyzAo7kZxWEvFWpg76Dr9JkkxOrjNA/0+OfJ3KT8NkJmKZsXY4DADiMEI5Fqr3T+KJXKAh
bx3CjuMrRy1wR/3+cG1rNiETpXWmbZFJf7JtelamQQgBB01LOc6bBmRoTEtipgYnDpe71DbywDnf
5E/WJ8NNhoJMbAK51j1WZYHI6TkC/wbDWpPJHqwSqKABReR/21k3J78Yh5begrL3tDcehB/ilX10
fmd+EmwJmdDA49a6velmgTmyTg2f6WCbMTtDL38vqR7DRtMnx/NsZ3da360X2DpUMOgEr1X+WEVg
wRUuzp+IHm31u9QOzeSflX8QSytNJde0m6TZpJ0mGSZo3ohaDZe+YG2JrvKbDXwsUe8CVbu3xtHQ
7quIiT9ksbIZiObtbLiq9uVQ5kmOyfKdSiZuOLPgchDeym7MvNgZ1gSlFjzkteyxQSIDXWbf4oy2
0cora7SkEdzZg08S9J/Tx3XDI3jqdkq48xEGad4+UsFWfWl/hoZlZQxik5H7fFdu9ai/H6AJTzzu
qJimnoQdk0y4MkcSwAHZCqKd2eMNyJ9iCHe5A2utcdUfwthvLiggRWwxYEvsKZyn7TR6iN3EYrmW
pdFG63rUWbfx70TsgXLrACJ9RZ59K3hvFKpG97jaGtWzdf1btiwxhlMcb7BIVL1v8OKbtZHfLvuV
XKRxJHrVuDmTiaR5Rt6acWnNV3pVhCogh2Po0MOFfN6zPpWF2udpKJcSl/0P8COise/zsaErJ/zC
j4FbKrLrBwZLF7zxJv8m3APyGM8uxE/Yu9/JhPhPllDZsWLHou2GsEm8UgV0qpod1tkydsACXjU+
rQO+wAG8iIO8R2rZvGHG2xNyWAbnaPLUij7f7wULEaejK7CkdhCfS2QzGunyZ8ILaFRslpAfLMiD
tvmFZbp3hprqE3Hns6TlSsLlOaY79P+rs9ZgyJt2SDVWvL0vWpTLix9NMRQu6vRax+cYloev+pnd
edwoGCuSQd1XUjCnSylOMr4AHcg5CLbaGKAgKHn1yWj0W6Ew1orOEqYQ3HCyxV5kNq8pC0YjFot7
uTYE6tOL//ft2wW6uZalZlGmcj2Ulm/2wEtyETJHXruShbktMqprk7QVB5rnqfNnxeDnbPV7RSnE
I6HFpJGrtaKBKqmPOdcebDPzHBDVkKx2aGkDdJ1X1SrfvCzRatUbYMM+LbR49DN2Jp3FD4q3OLHX
3lYj634yi3Ut/NflPSr8wCI7fIa9pp2bEixrYA3jlEkKk/RE7u14ea4MiPkSAStKBV2RvxGPv/kc
CWCN17hxF44ANO4dhhcTVcNCquXWyoO7duhV5UZPHQHUjOa13kfH05Szd3vN3fokmm7zOqH86OE+
lb1M9HM9hKN51HX+/5t4RcPLKvUSj80qO7sqccgLzd8m7BQhE/YZurrRwYEOwnHg+qJjorJscHim
HyAV7whNIUBWv/KeGRTkaRPQB0KlGf2cGJeh1eEWaEJwydnZK5XFAsqnYuJEcX368Ge6fR+Reoka
rQzN/MxCXhze6i/YyriYhu96IjB3r/QXnF0oOROSSHpEBmAkwh7NvzH46A6pxx32VBfYPPQWhC5P
PCnJVsdJXOZiMRo/qQiP4TJVllVI3z8RifwYWjXJBDUC6ISy7lH/u1zH2Aqem129V63ManQTk/QP
5fAyKQEIO6MlVKkB3Giq8WymP3qcwdKzFqpGUVZrJ/Ab9MmOv2D6Qvyj0rinCw93D7HUceM0uBj9
T4SQ4aPdXb8BS3p/P3mPwiyY9TWn9tnBmkc9hvU2Lnfw20YbiFgV/5yDZx2BzJ6PMNyco7ULrTdK
F05L+Sal1dshiF1Vzyd4EWDhibleYjLe9tKIaLr76tgr8WLx0TG/FR42BNU9BuRP58Muvw2EFP1h
+VO9H+KscdiWmi16Z5bD+ti62B2eTpMWNc1bJWfd9g2UgJnSWjXINsegQaeT4j4omromB9xR0p4I
myRjkiwrlaCDp9ZsQgJomWFjUOuUJTGj4K0UY7nYrwBvxh8ZnWtbSb75Y+e9CyyHyPnkyqxO4mOb
0DaW5+KVkI5dGlr4Cq8v/uByNtE9zOk1GI2HCw54Pr6JkFB31r8bZt1SWenuaKtYeMIfNI2rX+nB
BPrCrujxMY2txPmtz7kVz1wVmORSwXFB5gM3W7IovvUqZeVtGNyKBW9u6aK0lCcaq0Me/+2Xb3aO
LQQL0rhw6LGSj2zw0IbEDsWqM7Q9G5DKXFHajzeUwiITe2hklKILSrZG+RApYGKTDjnm3OTjgLYo
lJdKVgb7qjpT8KimFUDmESCxklbKP9U3a36UX4Clk60MApP9lKQtpNUFOKc84vUaaImUKWyqrxhm
PbZy+KFmnus/jr9qChm9LH7Y9FOAV/3cT7ivMcSQEuwNkt/ewb4iHKYYX+j2TWIZBXErqDsS54SH
/9E+gLMnhP+07euNzD1tZ1o5ykTDzCJtVtjUzHHbZbWTOmAXNHo5me9tUfD/2i0orCmQegG/7vo+
mNgg9g4lDx1kdxrPZa1atwTswBGs5ZjQRXbt2t6+mEp/VohjQlnIGbTihPcKMJQK+cCHbxpikzPb
Bax7WAPE6An78Jnk7Q9mFPMhXxKzCWqBku+/R8QA5/EGwA3/MYlQKooz6IHDVCOURL/JbuiaYJUV
zEcN/hbVSWGg6+VHKCcMBxDZQYW9EiUTizRxYz2tseYJLC3GZS46cMdhhXAFAJWK0ODUc9jan12K
/+8ul+n2WzzJbzefuymWxstyD5J7TPFQ2BkRgNm3RV5rQr7DSSmA/aOk1A/haqLUPzz67hPReIPv
3k2+vY3/D4GJPfu720XAmQSVKD2zoEk67/MiRqdlXH+etJUzfAofDlpsw2GtYalbA8pZCbtxVUGC
xwmv0fmT4Gv0G8jVk6YjFsLB1puAANKzKl0cIviipM3TXz+8V/qqQmYA/RixIOo15Msf2tsuFIDZ
CWlIctjhG9/H1HyX/Y/BIOCLyyn2LK2slZnE1r0l+jLv3xZtMeKBpET4OCHm51lbl4zmnQN1iUkZ
SkLIH/F21/dRc5JWIyjCoRxH8njwzwLuO3giIF6cbqq5KCvJP8Uc38dP4ulLsiOwAFJX8nlrZtnF
BHWgjztHQOC3ZdF3efiza8P6Fsh3E+f0qwanFOxv1IjoqvPFXPtol8klXBRiZR7HrwiWJTBCMg9f
ySgMh2FTo4y4qK4M2uadj/zpwnxVEEP1fEnOaCaP06Wfk/nPA23geLzx9OUq6uWtBfQsNJ+IYpiq
aVkm4VultAsVTGDaF5AZH5Bt3WYcPFNRWOumKf8NuTHAXlYdIPE+FfUFxIpJCPMGTbuxlyWuTECT
AvK9iZcKTNVewEe9b2JSxrHRFOzWNn32Z3wpEhIFoscpKGsieIAuwiYydjWgkR9emnm5Pn91gu1P
JCFTnvg2cFZTrn0kUvFABiOl6KD8D6WUj3STP/w21l67aaARo12Jlar59fRGIPIxmnlXVU1lUMWb
kXyLoZwBEAoiAbG877izStsoFcFNRgP8jtbdB3EjjN2yQ5aAt0IVuwKAnnPKs0kKI9X2MUQkIHAd
Quh711pVWT6OsYUOcpT8NqIIago4biqhbRHz2vHv1yF4o43/hYY/BcoD43dVuUcE+pegzGjFmYIY
XOPGVjbp68kIkFk3MgsW9B8bpumuMsP4uhnyLR1JWJforqqvua/9Xjbs5s4unlBxMM79f0k5reRe
RWM4qp/+8vMYpl3FWybY9BSV+9crHi37pqQSOkB7jbiz1PB3KfVbBCVTbkV7BHiH7OqyQ3h3i1L/
v1uTf+5S797thTLV3hOpiXsJ9tfYcn0Jca+9W+uszWrbSOmG4gyyBrBxTE23cyz5ztukOlliqgjg
WgRho0vvM1mrbpSvz0Bi4Z4+JsAAf3+iRABaeDXyPyYe7peRnDzWBtDs7QquHyf3v5wxlNbf2eef
Zi3u5CWDCD4gVvlKtKaI7I9uhr2AV+T6yLuvr4A5NIQc3Aqe/Q/ognTrRu4MxDUlsku76eWZHeAz
RqQ9/u6DyKv4ThLYdnKGMOahURX9MPMGcSD4H8u7G+YT0IEyhUcmWoRkVl9O92qX/2UJPxCkfoFk
6ir4PS0z3by/5rik10UNOol9WS62f8uJDrQc3/K2frJ/zYv0x8E3Chd82Usiq51uBSpkhRAhuB2g
3WXfT8Hakm7k6LooQlHyGs4K+w1DMO4xiTrTQT6dSh7o9Ju4dMplT8MnAwVL6TQ4FFYZdt3N/Z6D
h5l75EGb29KehowBdI7/DRUZjf2wWCv0RU1+LcbJotSH7ZToI+X/lm4cCIAIQZ0mIqhpwLvV/rB+
SQGGv0CLxSok/nFRGYmF6/Ag+Zj/Z9ZmnE3SPPeKM/TgUVrVf1CMpIzsBNw/7FGpKRxmnhTetOxF
gK6nhLD5kI21XJGkpBbp3rrwj+Ukr+yBBRJaxlpA7BY8pjOoqlnw+NCx0M7xsxmARZhoP/aeE0Wc
IuhYKHqt2WnBUjOWmUr2Y3t4c/jyVI09iEKNFKclZQHK/sq2IIi11RFoInfqjtw6LzItjJN8BXdN
HdcGYlfSmElsKxydaT8+cTwHoHcQv8sIk67wJKEzE1pei5xhbgcRQm3N0Al63DaCM1CRE3r9IliQ
szTtBdPh8vsOYS0lbAly0WwNbCM8/9fPkUVKRkNHzr/bTseN+xFWd7L9k/jTzLdIrBbY/u5O0ENd
8cIAP5II0Q9VxRkqMkX2WB2TvJum+NGPG9j+EimUdW9bzAcZshaHAf07uoCYpb3fnBHyr5UdHl8I
NpLiKTL/over9WrGLaBAJNXYnfeN5dB8f8s+rtLvB7WvsHgF0xpil+/W8/4r8zXcybr4CCJb19Tc
QDMjWpY7jrjq9LzEhfYoRc/nG4mfHCgN1yYD/92hropBpqdaLliFTe+NbmdD++e71MEiS77MhMkj
GPP4EgXwmVfzCR7+8EhuHgphUN+gWh4QoDFceNW1XtjzMcoXf4PFoasN0aw6c6Em9LLKl2IU2lRH
Or9pn06gX+kIK7bjsGkeuFELf7ZXOqlbk8v9kSNIf9YOtJHX+ckLgiGKKY+TedfUhzw79C8RHP9f
clriLZzCTt8iAuUduGJXrbVSTN0tV+idAjT4a9u8W8VOjMLKvtlKarGRZNfLfgcEW+rdJM3/vft3
ZnMKsk7uu2K3gWLqY0a7qHEnFeyXLJKevNcfw3P4jrtElb+//dVMqGIBEdURjpMkEiY7hk1x4WQn
2rwbu93v3QWIj9n7TTVjDL2zpaOK5uJc5RR4004hOUazBkL0+PKDQT4p5Hg45ujmaHwq82836P/j
cwpJsVV3CVUUL72OQiExalPUqa2pmLOhdRxzdr7LYbC//6N2slu1ULYO+xVvpDIIaiYM0oyYbqfl
4Y3X0/MLmX2QYnabybFadXnfmKi6F6nV29a/trTmKHqlDq+JhO4tlQaQDgY8kzl50mCxYxke9Wj5
3nHi+ZSwhPabgXVwufrOIlQcPCLWAvF6CNtli9kiQI1BObJfYb1oZ2BusN5ugeHSoLyAueCjzt4f
S7npZFTdLonXiPpcjZy7L/AMph9wAL4PzBc+1sEkH9bohPGMuHXt7kAYfwnWpJsTm9aIagz+LssR
icWdniP5cogse3vPYs1fHTsOpwvpfl/kzxJuOG19pPwMX9++p217PdMIqUY/DpLr3tpr8X2b4tYV
BSwCU0CKXdpNcGLImpseQaeeQcBJxZUOMXKgumd8eprSX5DNVwtAr/FyV1fK16UBkUgS7oDgAsKm
+CJomOH/EANE8ulkiK7EqNkkvy56RwzK/HApaRK5mJ6x0f783lt6q8PZGHeLNm9E/BR8w/OJp3fS
jMf10/Ec5RaPV4cKq09ilkvwHt/9MXcvu1GvlZPn5U/tC12M2zg34U6helut2TTulxVm+pvhLDrz
2BolZIhjkZrWgD2G4FpoEbE/o4kECzYeXCHQamQhXUymJCGnAfGt3accnQY0dsIBkIQS9hm8k2ZL
OxyBVofwtmL9KNkypbWUnLzx9Qfp0tdByWyc6lTwvWi0lE/jFhfteASRpWMryLhusm6aS8tyDEHS
k3bz1FFoZ+RWCfstDTZwpy7nLV5fNN0mFWKl0MbnyDwuMsbZrcj5zJw70tKHrFo/Yc2jqw00uqvb
uEJ+nm6ReZHh8E/UCYGACvsOeaUUvIHK1HXp5K8XbGUndqg3IW9zN4CNmNq569bDku7UfW6n5QxA
Ghv8afTyISm1PB13CJgT1T0pOz7qIJGsjpmwudWoBUmL89TEbmGd4pUOwaIKx5cGDxFXrY+EFO7R
UGErIsD6Wmy0XxnT191iUYPJHPz+pAyipkTM6wsrPkTRft575FQrBnFhjCThghOIiLEufqKTeJBX
I4+OtvviUc/AvWcOrfz26tEyQIBvnN4HN/bW/1wHRJDyas9jo2ifVxfDqDJkOvglK+8NqPLxse1Z
qy13KnoXrtQo171KQqMMVgRdtPlknffukeXLGauHP/3okaHubud8TlIDjFgxEfJc1A7zoiu1F3O2
BPokYhbN0azaH+wc9XmbAxa+aEiGtLxcMu7pbVXhqgNZ7Bpc0f7Q2x4t9qo7ZpMQH3tffh7NU8l9
L6mPWV2SQHBIGZR8+06FukuV4lhr0ypU2TjHv2DxDVrJknYubzSgn2UYQzIIPYpYv1ydpa1l22es
6J70XLvAgZ/vDzxji8WDeWmkc+ufotFGPKo3yqrKzlg0qYpVko27qifcDnL+eGQTjX/qJ6tCl6nM
ogT1iBEvXtFdDV56BeRSmJTCGLXe5+yjMfXRicb//b4m884GzFdlLCtfQ0F9G2ddjxjKUyZKccHe
Cu8z9lbx//KRBY+CDGBAIbO9VA2hLKd0l3Nr0F02aMcNAvFm7Zdg35Dl/LboYAgA1qV15wdTThxU
orsezRq0ZNpmRaNQy0yWZaqAMweS8UJkSRgKT2kU+6o0C/VO2cCatEs92lQhw3GaeX8hj67B+yIZ
LXx5axOUL8z1/j6BZFE+jPo2cfDnUIKgqCurXl0ystJBJUYEt3HPsqjaacQXvECWClN0z+H+yvvd
JYJOyDrmBg+f7hZiXGi5qN+/66O9beAh8mCalm/0UDAS5KOcP4dgAyV7Uq5/XkWWF/a0DLSyRkfd
BZij57oFqSnnebs9rgZpvP1Bf+5iEDfRIZmLSOEprwpzd50tbU61U5dt+it4XxFTa8pmLtfdAkpw
sZaEK+qLMp0q7hqFycJq/sEoVvnwcn3yE1yEzsoOplzlzO/y8EpqA6ZfvzAKLv6UA0IGYVY3w7jE
g2uueJ77vGSDACWqnRPiCqmjSDfk0ub4zY4f3xmwL1unThxeerABSXWDe0pylEmwW5tbdoFIxbdY
lDCSiGfSvzv+SOKsxdoof2Aha7C3/BDGeodmXSyKJ16eZq5o3wTqqUtxzr69oc2OcQnJIEz1oU0j
Fma66495VxUrD5TEyVQyR4jHBebX9MsNGXXCWUBi8yaTuf/n4AvcGGyxOPzAQ0Rj7sEVVxjp7/S0
KvKXAFkfxPzeK+pMge0MtQPG2j2gOdmg4ZzH5d1wOvHgTGhGR4h5wRzVZuMLfUiHc3oxkmm/DoyY
j32c3q6Yddm6pcuPl+fiO3CeGZCa6wm4OcGBhA92VLH4W9mE11AeQ3SqOKDtqdAoBqaXOmODNVqQ
Ul4uY69zpkdK5/RiUC7NokArxCd8sVkcEU+6VlkOiY8cz95HG/3k2m6lPMF+ELQzLHsDY0mZKxkA
kraC0Ya7fda0ZwjRAHcvbpqD7QS0AKi1mFaLYbKntpA9ffBe7MYcGU3p15rRYHvduie6hRFlqAaO
Pus8lCVc2bhRd+qkAl1A7L+QcjueLy/v/CzjejkXjm4e9PRqZrmXys8Qb/pbYP4FFky8kdGRqypR
esgeUThBLACvzEZkCWNkuS/aIDpJqvdhvgvvEzpiHQK/+dlIHAI3tr96uYqQtWtWtcoed9Pskdys
fHxKm8wdrKmoQofmDSzBZEuNoUPOeGFY/JqCx1GxnfBBT4FOxe08crryhBFBep9EB1yIaq3kiyPN
jdLqxcDnBuVjs9+QR4MInbpcegzLHNjwJruta0logy1IQjDg1vrsLdIFpgYXusNl+m/PcsnQ/VKZ
hu7KaO2gZCGIvXGIUM1/7JlUxGWjgF9GOEM7NmB1IyBFUGuRF0g4MLl8VGs3Df8eT37/vnqiXtJP
CEXPW10CJtifx+/r/1vGD+Pj13AHewhSqudElZwb/b7teqOzVWXm/kLxH7kfYB9EdiRAeKrJ73dv
YkEoHPtJy3Mar3NLCV6/vFJBRiK+jr03P8UKUVBYLU7YNSQZZe0FKoD2a5yuNpa7rP67elq7l+vB
WcKvLds1MjL3CsslEmpevyEcsQ7EVYThUdczJRpSzAGGeYmdWJjLsXLljx0Ff3LAMl7XZAS3+xAF
u3QJQZncZleruth1OWtdRSoFHPD2EFiTPW0DE6tgvQmbzFGjGvIRBV/Reh3PcPUuKPRSmIIE0OFh
TgY/7YEGtO94cQ4TLhRXjk7tILUWSHIIcvTvm+sh9hUfZq7wgXrgUaAhfdU/9ucf/X3u+0uC14Su
35drcSItuR4b+l8KCEC04k/kvEAuHZikdqeEemEUUQuVSL2OLEC7U/MVSi4cmDV4E9vitY4pJdx7
/VHEQZ4COs6GRPtR2NE+flsJjF5j6g8gZGXNP5GhC/i54t1wZ1OHAC+Hgdil2l2RXribrL1V1aLw
GW0aUZbuft+g/pI+AnIfzDjWFzP5GjwAx6QrSPosWWHIR4aQRrhYFk+RHjSLZgnbcydL1IaR0kMZ
CyOnJbN75T+6J9hJwKOq/0xSXiF7SL3ZTdsGtv3xGdSqKy3R71JBOWZAua5pevgU72yO8DoLT1ph
VoEH/eO3h5lACI4I1J1YoD3mLtjfYGm3EZHocmyEQUPVLP6Oq714zoVH4ERCEz5lHgcIkgmUW2ef
hop63BiUHGlga6XZLjJYxza6V/dIjqvsk/3j2M4/mazhdkrb7QH+fXPYaVRcPEyc3cxhAfQTWeID
0792SyzYRPmNzbueEZ8eA9bUvNBkGQMNPNHU0gw4+C77Vcb7ljczvFijz4ZDWbYrZW+vx9OOWDwA
Vw+DQD3zrg4Y/ZtfmvngXV0DN6Z2EE3ShWxVZ3cY9V/0o9ImjrQbRig/3im7eP+bL780Zeivl1Ih
KUEvEsVI2qjiVOTGk1mzq9Ja9daXi2DtO7Kn2T59VsN5b1r5Ve3AOdwpV22d+vHLiem+2HbYdo68
5fO86ZIoRuoGaffx+05BleLKyyr0lZGJ+JR7R93ElrhtC8jzYXSF64USAf/yt+2mziJ4K66tkr9N
iH26go0vCf0LaR+quNKkr38d0u9rvXdCaBGNd3dH9e/V3ls/WhaSTKc93kOAT1LenxPOonPWj2eL
h6HjtFaxQXs5EjwDhQArIspzhPXK01SOjk/AcZLgsjd84830ohArNxnTHiZfB7oXCMuWc98T0Zdb
/mbdico8HxQIHDorhgvfG83DjvKeB7ssp1XbYfRl18mDodeD73xa+9+QXu0jhX25n1QMEn99ifyE
OuioP0gG5RBL+LX4zcQAaIQaLvWzNJYOaEBTp7fo6Zww1jINGn1r+Qzs1UJIFBD8GJ+Ftojul8wV
rpNzudZD3yhEqvaiMxIEUK2/pDd9gkfOQr3RkKEuhrQDMmssPu+nQmzzaes26J8j3RnswEZ4Oxrc
BPrkmzftJBm1UouoS/sq5U1SKBTAJ+v9H2xYgn8KFwenRSZI9fLIylONa5il/FuEUzR5if/GUG4G
kJDd7yKaT04Nk/23vvy9PVwNkXvro54ZJiF3uEibkaPbcd+trf+FlIV9dbW5O18Q+ClB7PtmqAtA
3dTJc8ijzqUm4M/Uqmn5uocnc1xCk70kVvkNoyn4sCKIOfoTtaLPGi7SJoUWtnGbLmpEzpp+FpMj
Q3UMaR7BPUYb+UhFyMPWvx0UipFT6N8UydoCMGhMp1BVE8ie+gIwRq+uyiuLyhT/HVHXxKIM3eh0
Tl6J7DrC0wh2NPQh9YLBZFVflGJ5WT7XijTOONfO+UbNcgZmUyuE1qWNCqIlGGO4XODZsfwtjeuV
87yrjjOQaoehJgwWqX9SvTwyv/4dO/dvJUJGvsGHfX+rNHDoV04e6GFsSojh8pZCoLhnypbTUOzz
a4GSqXjd5ksg7WS6Kq8KI+aUQkNMAZbni9aaKcPiHHqZTz1JrfyrfzYjMRYOZK0M3x8Z9yLJ+qml
he6a2Q1/6E5dIoZUMuGTHyhWYGpuUOUVTf026+pA2GDyf79u/GPxAPYX1/8+fGNajIW4r193Lohw
zHkr5VHYetyP67Tn/g2PeEA+j2ATikGpXVMNiekp84Qu/30AF94dhcYsa7TIMAAybd5AjX4ERNim
O82rqPCk6Y4P0wqjupWwGd+hsBYCt8B0/znyflTDar4Bf5GxefPTsyfATasK19hHigMylTWMi6wW
1Vmea2T1k9e79AijPNqfPB/qoZKXdqoN+ddmKyqehCgwvMAd2Eea8yEbrzNTnd7mzqnD9ok/2nVI
DxTjGUMrdt8xZI7N7ttLdPcl5DOasBtTqw04lSHqD4MCbJwUm+p6p+T+Y/iAUhRi9eelJq+3R9Qf
BY72dyLmYEKGAEqabNCvDXAdZ8cwrOAS+nytAyihGdK6zwPk/SO4oUetL6xLRr1OGN5kMDHwN9cz
UGeDI8vD3TSL05ujRMm2viRH/NFf5u49PYiz0AQNhA8bdcY9g2+YMGftkamUJ3C7m2iNd74uQcHo
rfxYq4IcIfOXwDpXYsz+GEoYnQcM4WvmtpcrrU5TuPDUTpJ6jbnCjb6YXOhlNl6ep7NH1H6bpUp5
S36/E+IvzU7MF5iI145A1j7h6DcEm2KScPKX9MAMWhvsihj98w8kPPZlGBXEyMzi3wxdHy/82A2q
qvUTxY6dbl5Dkv1Pi0akw9dlSjnQL3sylS3DtSrdWtqjESQrggucqwGu6JI9yRjb7oYh7P5CIvlK
0Um6/Wd/w3IGkqzAIV08Ms5hKmlv2Kbczkv4o+rNfQ+UzaayjRWxLgIbXcBCpXN65LwyrXOs2JIL
cN6dM5kxV53nEQy763WLQbpvOG/VaNWSBq8HXMTGjGlY5P8Cgs1lUI/xXFXURZkg83eNMox36mwx
2r7gmFsJ8DrJVM/zUmyUDw6zTS1Ff3u8CbBczSQp+K2Z8qKsNMAmwq4Y/vuSsJU/XwqNTX0PySNQ
+uuhWAIDs1wuLW8sux4KOq8GqjH/my0mKFUh0U4nP5zFfCGk3HQubqBk2ZTyDLasVVfBQBlSyRHH
DIAo5Q4YuqPztHKC3pjCZwMLTCtXNzkPhErNtg5EIvvgYXfYOSj9JelcKinijk4gD6h04a/NnwBn
4sy2geSIIlAUvD+O0eXeoT9ajUUPx10gkJX3+obfsRKMoL7IM8LMg/k3H8vxrpBf7+VZwI+5jZN1
CF9WaqzkFZFZjrpi/zCeUDNLlzHZmjhgPYqMY9sOue9DUQWh39lK9bjk+zgNZKXJZFB4/XzLWWkh
wyruoICtri06jKhr3bcwc2r8Ndjng90nw2gOQy2zSj9OjK7xdifnuk6hL0S5/pRfKWusBUCetlXY
aLfw81LJ/J6LIZuZxoilcVmMFl0qwsLsb+teWhUwlOdyEcKLh6LomGrjXUEWuv4bHWLy9XKb7voI
m3o2XNWfcUysNbmGzfy6C6PpB2EAG+65KN5JJ5kFCo2x2fs7NihMO8+bkFEvzQykaUOujO1DnuOl
eMZ1tul1bwJ9QB1t2v9jUcjMW+00TR6FID0R0wh5qCQsLZOYmdiQtP1NKoE8wQoHzdpxxl68wd/l
U6nFzmWuGXyYu5KIV8HYe9qhA7QoiCNuA+U3Ks1TaRY8Ev6nmpPS4o7I3G45PlwGLt2fNjgT/HWu
Oc6+PfkBqjnR0xIONs7bbABhJl3i1fEnRVvYIeOtrkyYQdx7smRU/0du9Z3BoMR/gUwNa32c65HB
2sxJMVIYT7r9Db21jQC66liYY0UM/o/d0n6YBjssktuamXSlK3oHFEZUgpAhrMgugj0hT7KOkkdb
DJjOd7BUUbteazlubimA5hrdXh84w6qFRtIcWlqPEK2sLJrv2pLjbtbFPyPXCYBliqvKNop/FrtT
gjBG8vbcVrWAeGXwtDDLUtN7KMRip2D16E2485Ec0vhq9piGw3DeVAojl54UFveRpgqgvfl939BB
1PHucV+u9qrQWlg0X/sxrhrWzmPhSsKq5VJAfTWj5HiCiDHzv1Shrpd/FRGUogZ6bkT3zUzVWNTU
qlMRbJNIbk1HYEi3kx8xfd++H+/AQraEBhusyUharpVby+7Za7BcOd8kBU7JYFLcL0lwULYM0WGy
8blf4cNjDlZ1tyM7sCKMk4OLCA0NC6q3YPbQ/ZdmCK8xtw8QiWPLiD0Px0cKeIu7RqPXZ5UGeSex
lB/Gd6MKv2GFVudw384G8qDyQh3QCFmO2+DvL6AIzM9ErtN0Y6UGPwtYUpwv5G/6wh1e+VFS3m+q
LhCJBL9QJfgHMcxZFK87pBnU19wERoYZHdgVDVzYXp14X0/ya4hovcKXhfuA2+ZbuOJGXsw1NzI+
+PbYpoX7As5nGOyzrhCqqTPrxnzIJby5PsM/5Ze5lRxH6xRrRRq3cEWibvA7wi96d4GGawHv0gFy
WEdlsV7MCyAsG+UoVcaL/g3dhCUL5D75XObmeVxpyibd2q2664tQlytC4I0lG3VnhzJYIr76D4T1
Y65yJtV3zggr0mJU1wpdRq2wlYRhcN3dMB1TZQvwRIBPNyQrM0gsYNBYydZ6II6KkFmBKF0PHoz7
IHT4Cnm1dgzPIl501NCN2w4VDPW1Lu0IKqrThk1uq8IYRCVgIw3ql5bjRw/T3OpjRSQPPs7LE9fI
pSAmVVJKK00MVV1JVOYzydfEavERdPhB2E8LkWjZLzj2CP9smxAHazcOATSwCNS7SN1RrEqCkun9
qAVppuxdIEO/GCxGaaG2CzNIhbmnIekCB10gzpEmxFPzkoVg8ETAGveN+UXqMTQOc2CNEakGSnjW
Hzsk71NWFHbmn7SqRxygEcgHh0x6O8pjXpn4AkFdjTVmhGeP5JmKoXCscETFzquSjLYhI7IkcA7r
179wdntfZJCN+VGxXVxjAmit82k9rEXsrG8TC7ysmyUMgAAaoBSy51DNN1SpPEDR2axlTJXoy+Si
x+ZJzu2F1aVbH9Lrp9yZYzNqS6QJW4h6wRORM0cifNLRklzbmy3IWzbbMCuWu9sCvKwU793g0PO5
zZnI9YDL0Zh6PdTiDFoDrPfiNB78N0+T5jN3YRb/jMSwRXp1kLsQ6FGacYxtLmtkSJoq9otw71L2
JxTrhh5izM8mj74p1hjB0WRwoJdUsaaEOrOHExcyxaLloxIg+S3FfSQV4GpNbgLImIKcdiX4oZIV
vEpR4Lcn3uR2t7PDjDYKRSW2Wfwd0Fqmi9OOxIV44XQquAM126lINj62Cz3WNNpIqanak8SaIia+
lNuheMyEIx8kCxh008s86Si7KCoVz6aBHWX9KNgmdBHIYeJR0684tSd7BK8VRBL/jhwtDUzppPNr
Uxxd2VnH2SelMX7rvYDxPwoKZfNebPNa+1VwdPkyvLsuZnsigPQRvbt0cuVAfvHcC//rgvXW33Bx
Ft/j1584wtCFONdaHF9LFfbBe1X0rAXEG5pG0yrK44ErkZfSiYpfsx90dJAM/cBAx4PUuQlEFpDM
mDWFYRggMjDOQLBPUE3rltMaFsVy0bIcxqqDSMSl1sDfoO2tRjcPrroKdFCVfwI7r5ldOXe4+6As
FnMaQ9y2ZMoARYb83gBvQRaTtfNnx4f+svVBKQ0T8v2qJV0k7PUfLvv0fwUCLB2b3AvuxsTPyHDs
JdzgrUSC8e/GdyDn+k+7bQA5J4soUchoEOWDWresZ8pEEAbO4FYslJNC2Gu7E9LTVwOhYiX1GGql
kp8yUrXkBtFMb2VI79Y7+mhCrFy8N+pwIDRd3QrAEGLTcrbyBmojUKgsw9pBsZNUOJNftAPfJAAV
+gVlNgbmaHooRgC5KqboSRwWlFFKeGhLX5i29sKyKmtXsqCN9vDSWTwuzqQBVhZSHZ6ILsDQcoNw
X3kbysZUuYGg+mnVwC/6jNi5iYRGvBUdn/+8NWP2tvPWZljwzNLWxBBUkR03a6zKw/dA8vdbXJru
GZ1RM6KlS0zhoibBEr8BJebseO0Y72XbMX5xEN2Fhf/er0oVAZZJUc8iS11/x9uTZ7qdGjnAfL2d
qOQlzJ+yDsyfCJEPWHfYfQcgAgp+EmKkw3sN+tqvQd1JwFlH6vmhFKNSbk8bdxyXiW+x3qSe2y+5
zyIBba2I0Zc2RInxzGXagh1XYlKN/3trmveZLct39Zuqp7jCHTBnoxpPk+hzC34j56cC3rfZOV3B
EFm1DRYWhL0ykEGPrIK+bvEZ8cHSUpm3o7/+e/Fbnm/CJi60stMdp5fpr+lw6XIQAyAeVlsC2fja
ZUaJKE02wyl+hh3UBS3HHw5y7ezmH6hnFgkWKLoowtz0kOrJfqp1OiU3ttrsJhApt3t3ZbmsbRmX
8bMUfvWLXxj3QkiVr/3d+ri4fL8U//P2eNRd9snNhYE6uttJlD8wnJ8s0hNzvEoS5BH8curbzULn
30wXwHLXBcNSvL3eau8e7x7AOMUIEmZK2FSwmPAn1vFJazyeuGwtkJsKMuttqF9QGbFEBXGLdgwN
HaKDjF6UQwgsUqx9FwnyGSHC5bg4F2z5R3RBodiFhcnCiLSBzQkTyk0IKhOEak/6o8vKv4BIy234
jyWi2SyKKHXfTeHLEFoz5L10v5sbOMxHIPeU0b+LhwiaNik+9/CAfr8QEUQUI5TrAOjxicws1BAB
hA4GBtaAcKPLPNqjQLJ8gQR6GuPwYruubVWvF1HY8t88HFYYhYYz8pe1pclPdOGplkk1Q8W8KKyD
lBw8WWVcuCcDw5BbcGq009XT1u9pMJ1BcCghYP8mj8Y1jmOSU/Mn7MTbj3L4AIW6KyQ3ZVu5K9mU
aup4Jwv+ymwdMM9CtIZA8HGqgVXpowhitQH7jLu8AnSd1r2Y2nMNnPib86C4XL96B34J+Zoi4zCd
LhVFy/R7vy50mTgPv34oJ76XCvRjdJfdWt8ETk9nNMOpRz/lw2TWMVAvdw359k1MG0GXBjA9MtF9
fw6ufjaNGbs7vGT0FUnPEh4oN2FSgqFNPhZq6aZjxzi7XihFDE6IoRZOtjMI/V44pHqVq/TXSbx+
QlxSzFU8g74rww5V7ie0yzVdxXJbngaXmDIPrw0KN9xzz1CETOO9P6B02Z8R/duK6b0YXLEdAWKC
x2C/5jn5aeuPS17vZ0q0QVXQ7rEmxWDR/gb0FlURGEdFGcmBY5oRaoKPEEl/UwTY3XumkEY0KbXI
/QXznJSQpsHmHQjzlljgrNr6MHuZm4b7/wkd713yc5KDgGaPxVXpI0sf+39RaTOBAwOWmy1vSJpk
oliSvQEBEXTab3H1KboNnsvlAM2o4gBRg6EXmP+vQrnII3fQXkh5wmzrttBrpn0s9759ZrDlY2J3
8KJvFd66FVQ3lSyy6AjsGtYmuvooHNnqmdJ66aKAzf2RVl3emmJ+wOwwpTAattcE/JCDN572+DgA
1yZUdKWD++iElEs+YZdadjNmGWIid5ugFuw5odktrAAvvpAiJIizvD3DCnWyRx4S+/wZjD4YqVzL
And6f+79jfaHDww326PohrTOfvLcCBZX8z181CZGWuZ4OZmdpXKcNZ4u4t/Lwrv8JlUX1ULueCVB
otizsIp6owdFV5LGoQs++YE47WXHCPnnotvdkMcu2IEZlc4i4jpvqiDh/+pyO/4dSZ62pHbGAMWu
F2+4xoReFJ95heAc2tUSdQ3ag81IY7yGirIOwCsdsIFXQHz2YEbRPRa34sH4E8CngtFIrfproLk9
o+CsayZU+T5Akh6SSwFljGjq/QHTmuCRRVIoT291cB33HTn6oj3KYGfxnL7V+IZbmvsyqfI20DSB
O89DqX9BZ/tvS7qG0/P/y+N575nHPabuwAk2bawft+Iuu+E+dnzzlJl03WjQp9MCHPPVrjjQY+Sy
XJcD/0WXut/tvPG5/y1msWzHzJoWT2tQg/e3cnK2OLt40/LjLPeMrTRDh5x26IVo3B6wT2li56oZ
oDopA1vG1HQdC7PZA15vjTZuj62pSITAKupl2lvjDxcEfvWZRLVa60PY4jQgFq/eHziOGvIJYNfe
1E840YTaKEVHBDnsvaXGs5nAbBaP1V9/CGvUpHPzypi5Y1FQpSkl8tHtwuOIFUVPeEyTFeoeLPjL
0mAjaBGcWM7s+iDjCbfjDPqzV06r/UsafF+OL5tUnK37pJQKFG2sFenNy/dmDMJWselG2yXajjEz
sgIwuJ3Kwb6XKLBRw4/yAOl+UmQI/YKKXAm0dfnYo7GsvO4EsSC9efJ6YwA6O4IuaYer8NfE13gM
KCA+t+ELLfEioVxPxHC+ASeRhOrqS/SndUpraMOTgJzlKyjip+17nO6VWtWoLvfHcLbZ6Z28qURy
KPZ6SQVGPobLRlOe0deiHsqTUIhY90gEJnhA5gxN4PS86YET8Hgamd2UIr28AOQB5uhPUKBVRSmV
wnLVmCT491bcEPGW2OTpDhRsMmMqvo9LOShDtEDQKq6cifF+JAl7hdcIrO4J7GHvS1XxGWwC054G
0S0lp5iEpJS8+RdbkyuE3M70ew/zCw7FbcyTEoZTIVHGnrobKlycymo/4Z4zSkcsubFdgBNyCqGQ
1BwnlYdRJ/uresS8Ju954jDVGhpcqpfMvfpYPIoXRtZXMdaCa3KAF560Shy4K7SF7ayCa4SH8dpN
dR54Ed6gzibZy2xG0aQRwCyr8nfUFJMNdxOGsz8zMXH+NDYptmsZ8ZGoLToa4+dXukh4BpkxiN2w
jZNg0ICaoAIqRegINmJQSyqVWi0x+6RH6AeOCVmP6Fjw8m4XoEGZCUwFhKCP09qSIHPuex/ou1Kn
HRU6+UDEtJgIQSSS7W47Bqoyyd8495Hn9sEqum8ucyfKc7EE3uMEl63sEuoXZCc7TVF/CELIFAYj
5l3/eMV/+ZUjedKK5AWdCtMbftV/98jTMh6D1PZE6zM58ynbSXUpgdDheCH9kALB9ebTxi8UGRnM
25HlLUIBcOKoncFPjXkTr3nGkZtxcoyXUMVLcPQ7eSKv1UUYYkZI357qukIh29Y94/wU/SZYZXuG
8CmKhPS+vykCTtYEymOAl9RIuiHmo2+B3OtewAQ1D8wDw6V9mvOk4cI4lNq5dtdCm0MitR1icvto
jNZ8tcZnVg5GxkXfmxf9+vY0n3X72WHJnDZ4ZEOx+XvNYN678lgxCrpJ0Kamy8tFHr7foKJQuGBO
Z08Ip0S8F8UdOBULi2R1jZHWN+qITLsKZ6TApVM3Oxt7W0UE+trlhPufhmGUKSXmmromkUdZDggS
4keUxPwjKDjUMvRo4Te1tK9LPLRflFECMXVrv7ZXprhz/vhF8Srw2DHW4o4RrX1Jk7MdGoAOJq0F
5A6tBs7U2DzyF/22D3qKzBjzEB8M79DHUOl9lmD5PNrA9IVyQHnMprSk72RystQki2UA9DisbXb9
EAztYjFo0ItnKRsXO6FiFyee0rnFIJSQoPjCFyW20MEO4/9eOpzVWQpaD0gNXt0uRtXucZsw2o6/
8G+A48x1JTPu9QICN7Dp6Md0gCENX1gIJ+j4jci5BRbMtMezHke6FA36lzjCsyyxNs7I1f5J2tfy
1OYHzDmEHv9RBRqDQqLKRp5YpuYwolzhDkxrDNn/4vQUE2AC7HgyHWyd0OOdu1bZl4MAbk8ZVoSU
NLOEENGhT2Q+tGSgWlRYe3tdm6K3r7io3miPeDBsCNtIAuR1zmkNsQjHQyXdA84/vbr14nygFnMR
j+MWsNMbY9MFEpRnLrtXh/VzEdDeYx/ExYHgVPv6bc7/WP/Uhj2yA2pERpR/Sx2OesMc1AQZ2Zc5
HJ9h+90zf4agbIqfi/O+xDeRz2bLdZmF0hG50UPyY8hXyfBnmL1kWmj0MbavKBQ3q5k7pqvOapn1
evj7tPRsxU+ndMAuGq2eXwvgzWJBO/SlfcDsPV68LSQIakNsKS8DzxRqX5alHz9E8fbt9oMNvFF3
BpPm6maHK8ww9KipA9xC4kxLADwEZcY8mFz1ahPZ54tpne61AQVrbU3BGiiAoCzz8mOQJJQie2Bi
p4917YeSTPCXra73BY4UAN23EjtdWCo++srErvvl3zyXulEKOketcvNrCRMV3wxxM/qipKndUbiT
gwbANc3IYH4B8VXSmHoZ87aLwfX9vXdSYt9acTYQzatgxBbqz0nepfoAGzqTlZOpJvg/L9KmqSjl
fFkjmN8/viWnFMo6NxIcondBWpQtDBHuZMDnkJ+mJdkOZHg55Pypa68gi09kT+8VmxrHeuQj5As9
1oZfPg/r/XCKLv7OhDXX5pURrJfobrXoo40OzfS0wrtRW4d13KQUE1mMDbHHQpWvvC8tt9GAOwQ4
CqMz/vl02afZiqg3A+eyw1RMF3WlkHbAGa5e3dAanxrwANbprwMHyjZYyg2xQ06HOAdQNWUjdeLP
wH9kh3cQCfsUqDzPiBFo2Iv6wkorHj+Z4+1dJkuCCKcuHpn4Kt0IFjUYu9dspwycCdQv9Z25dOcl
iSTUSNs6k8ekKIL8nui6U3taelRgmdVt567w9O6nMJMlKOf0sOdMBieKlHAb5ieDVJF4f4sMKBHK
2bMXXy5WFsNUtHTBXZSXXshbWecckJAaSlkc0NhuRE9pAKuFJ7EDO2AR7fMD/EIjf6oaXydEXg/6
rcBrqIHhu2A7oJpq5tZNJEdtBJnGE5wqTgGUDgIa50C27l0hyFfAcjshhislR0ZNdI0Hj+mopOsc
Td7ZJynp30xy9LZVUtvernkGOFRdzQaWj7BCaEmP8FPJRh+LL+Pmi3jNdHaE49jXox3OUH9I6r+u
xwY1WB7d2geZkGvxWY+xVEi4fA92rYTLzBIOZrIcK5/AvGRbbP3e1PloD0YzadDMKxwd1ROa5+h5
r05tagrpxCTRgw5m1DEmPdYeGLrEJPIX9++gq/bpRK0+58wiz8pRp8ZUNhsFGMSLBIp7z7KP4ScD
NP0xvBzAAeY9XjzBFyyoGvJcRCu6AGThv/baGN3QVAj6mUjfLY0Z2M5iGFRM3thIRbv3mzUd+YyE
qRMPcHYpfbd3hYL3l669VD1ohgLQx/JklQv8FfJRREyauUXHED9gaHudlC0h6ZCnwSSCYLaKB1M2
7zBZnwZSs/Pswnc+pQTH1mNxlzZAgG6rFP/lSaSi9r8Xat25zqCNXx8bPfnpqxKp2ADv/n+j4gpJ
27/T7GezpDM8dK/uWFE0tfsGNUkY0ghaJEqxrP4HqqMm7i9BP2OwflV18uYF7jlb8BhhtlcfoSzs
tzX1Uo+Vxxzl+3ICFxjc7YMJ0NwoAOhahp7zFhkmL/A8Q5dDEyJqJdrp8V6nNkFM9yWIr2pD7SFM
Rq1wfmyo8Alsfx60es57xUvTCIaGYS3Uh6CsbpZvSdepgdUxAG+NovLafPb6zRQf3s7zNP06GmWC
rj4Hn2x/3/L+shgpiC3q/yYLF2MF7XOgdyw3J9264wysfI3gE99bHAwglhLSU4zdXHpxmU5/YlAn
C8tytJr4vFmcLovrzkOfA7YwZgl5l1TD7R9dTkQQi+ut6edBmzrqPRzbALQIPCuyWkWj/E9iJsqi
I1uoaSi4myCcQGAhFptReZ39JmQ4O/crLKXPaWmrmvUjYHfWR3UsvMi3sB4rXCg2+EObbqjfvnQM
eCi75WMdpMRjnIi9jxB19TPtmOTYqbqQ1+KTF0TqTYssUxYN9RSRTvQpxls5kZwkT8nSH1DwOKbW
zY+d/IXfTmTpd+WWiLrVgVzlAVtXGjIP/Jk7GBvMYa1hjfC+iYkzJxhOFIrp5h018QYzCJujJ3YI
hG5MIgP1rWjDNws9/UiS+QderN8zZxGinqn7xSEceq0/qp8+QmPvxi4PCcaq4K2uicut70WES22C
16+QjImgskDAUu9PWshwpD3KHLZjotNqOkbLQZmNVpGqI8jSt8WD0uxbSzblsENJcvV/mi7YcUMo
vObgVbarpOIhe0p9PlQgoq4U7Vw2pRq7uCj46OK7xc278nTrnlFSnY/2cImb1vND/6m7Wo/mdpOG
ooJoZnU7LCa3+N3YUE55itPn5jY6F7ovCv1nk3TFI34PdWdG+V2Hys/M/A/xsO5T/rUYL760w3p2
+S5Gyfb8m/GvZ2oXaXmB/iif9gh3SZmnA+O83UjjNSqlfkjQAnVIAhbzMkm4oWgQQTa2fpL/x5PV
3A0UJkJQzYCcHHS7QznVoiH5olYMplyBRQlOsUv78xUvIuUyXPyA9LbBovTCIXwHevz8Hsn3dENo
d6rUWTAVg44ZfLaSiWbXEJx6W3dhgVxzmd8VLr16vZguW1B6WdbB3dUBCPi1vuqIQutxEQEUV/dp
XoBfrh+qcoX0bwe8rGVNmJbZGVVYCeljea6peO7l6F4LPz0uNS3KbXiuO/hge6Ap+EKhqQJWlZpg
rsUJprJBOh3Wx7y5reSQFEd4XxpQ/G1shZQBqLH/WL6a4gqCuRZGsJOriRpicLdiC6t5brI8rg+6
dlT8XTqhoqx6774aGWkUTfL7lt9lSHrpfhLRARJvIr0PEUPzKfqaTBnGUxpAQPiz4IH9UGRSdSCJ
d5mgiy3U73PfbXum/i4NFpCVdKzkb0ZPA2xNC1x8sC2uxL9ElmJg8p9x4v+UtCGj4YFPlJgYU2/Y
x5QP/F7RilihJmGr5zlLfhR3LpgyS5ogMjbfJT58UGI9ATQhual8U4hij3Zm6uT9yqoD89AS7vyS
X3I4TF2MiIiohZWsVr1bpTB6/yCbuh0w9bjWySMLYB6XWktZRMnXVO+GsgI/xpHABGcn5K/w5DhB
NtJS4JzfeGlpAPnU6Feypmq1R55fvLJjcGDG0G2zvC2/55tTNz7IqijxZ18OlgwGJ+NQrMOHbMRu
Sm86csdFb+d3FdhirF7QCYGd7J8t+2FLxX8UUby83ARVt6IFSHebZh9/K4aC4cIht0DN0A5ja2MN
nIsw39CQkJdq1SoPZVJTVxltcOs5K/dHdmyS3DSu5NxNo40VmIBtJlc7E0PUustj6toG2AmU3FU+
MoVF69TR9PiikvOR1ofDF7eSiGPNo8PzRZJbyr8gn740zDxxHyKDml4AgdUcJfXIvXot1fb7z9ey
KonJF329CGp6mHSVK4+qw6YSqjIFjOihAqUoSbR3ujo1V3XrOfHHjWgjndEp0ZUit0h5CWTRnijZ
A8YXThvRYdNqM80T0uUgwEHIt3CFkdgaL8CW3VTQ+E1dV2/sGIoH5SA4XbGQV0DBvc/venxAhcXz
pHbQCLBnOL9AsQIYmjeniRo4wIPA45bEaFlpKzp7Qb3Jd2K6qg9UhCVYoyVdpNIvXLIlLzgvhuLk
w2wO2iV97JNnK8nTC+Gp98uH8ZpKIXi4MGw8W3O0W2rZoJyDozjiC/OfKDPpAQ9eJSQ58kvGlcKP
MTm7+bw/bQcKQIJ4Y/spHxxT89hMl1Q/XHEvvCxr+ykSSQybprADuVrAUPPV/QnmvikyKVp6TMOx
wtkqFxgzVdnf1lGDp4ZWZ0HTD/Ue4G1h7TKei1zKG6OE05M0mtHKpxSPd9/er/79LGwhJBweyvhM
fTueMIq78PtzDjsF6yS8xIQ3+fHg5CcdMsQt6fKdOAQOkR3cuQKYv2+VZViP4rUv8/xv7xMa7iVd
iXNhQLtKDx/ZsV9PAElJSV454eAv9KG9luFVKwBjzsLNTtmIj17XWGDnR/5Ts8/8/5u3mx6tyciT
1WO51n+yqp3qMGULCrM/Z5KmBa1K+NxP/DDEOoYw1xoxJvV0gFgRv2mFN3K4SFt3kUrdny95i/uv
HWLDsWA+pw3XggGKVuVk5vmFZ4IvzoQpeglWdYO9ubA4YN0fjnUURpm+mgPVT7U6v5uJPcHWeJoG
BzU6l4BcH535JbGeGFEh7PqhHriU6nPoOghu7OKmxlQA75orS+vZNHHYbDXmoXR6ima8TQbURRIs
ZX4Hmp1k5LAzhxjeAsKS5SbiHhuamo3kmowhyvNXCbL1KEdhM8gnABZ8ighqujs5P+LkakS9qvOR
K2RpNWW/sYJmVmmVMUzicWc6+S52PS+K6uhF13+6n3EzTPOnfJLa50NmLKD7co/vsyfZic9HXLWb
nPVLBNizB8ZtUmHu0Mves3iDZIuD6Eyw94p9H5Z5K54JfBq4G9JkFvIaElUrht/GD5xqtNDPjGuk
SB8+P3Qu4Q4DlEyUcUmB3CbyOLZxcoAz1+Atf4/W93+xwSY/KBCqvXiV2RwHhHE5HP06UDGyoEqw
9H89QvRp64arE39/XPrEJ0jvRgU/z8+Yt0OX10r/Tn8SGciAnTSIEAUxfymqVIIGkiF+jH0WDPNx
AnUYtKGxoKs8W+GQHswMPERv6K9o7PltegzJYvAbGmSrgwiM4j4ZxZD/gejvuRKJHeUGJ4XIF+oC
jS/JEuiLM2I4P3eN2EWTmFSdIVaSqbPai0AVsDJyZkyMQn7yYT6FMRZxAM1kIcezCs2iQzzl22IB
xTIPHEVd0Mqp+UNSpeJuHyqluHFi6c1kP9AVf9V6tyDmUE+GGwUvxAgVayxu5T02CVaF4kw8N2jw
yjfunvZalNtwLtY7HS0IdhcCWKoMvz1H47ED8MRM4WRwnqpfeghTDkXzvCwJACAe2qn/6JQKDvav
UyGcj7ZkKDZwDwBT5zU7Ig3llLT2Y5F7ZmeWZQrZcfZdKiszVhsRibeh/aYmFrKhISrLO3cynB2q
euKwPuhaUGETbVSVztj8UNjeoqUy1sKOqSpW2h5PtjgaJfMATNeTX60y+b9Qmo/7vrjIiZBowD+R
t1rs+vNLeQXBBoMoE4UQDc4uVD1ZEXbUDrCTlegjAPXghm/OYBdZfV6yhwZzng5s9j97BHvkgDKl
BWh4n0tH/HNt+UCj8+vvStmgVwfTkdKAVh2DCBWpsmYFmpTo33g6vYQKAuD9jdvwCJ/ivIBmWXO/
XPdlpy5iHyIhQof61TqLdEsNK5UtfHJNDV19tuqbsS7pR5NhU86get9C22ddvL1ABwFvy4ZKImf/
XKttVY+kM+Va8dNpyycViK7mdlD0tvBy5xWs/Zrdzu1d2DpnFWCg4ZP8PUtMT/g0QBH41JIwctjg
QEIYuLb4K5moqifh7+j21PpttfJi4PTm88kYav0i2+f48TJrTBG6mN/hH4W5skRtiBVTVZ7jKmdw
CLWQOs05TFc2UeFwkyptPzz6P6z5zmmg9TxtGSwcUPz3RkH3S2vOGztRsPHIEZweru26H1QCRlOy
AtGh6Y/JDgMMfB0rjRuKyxEamLXzpJq5ZXKHqF5yPNtJ0d2YRAqOcq39uTDfu+hmUPqvL3MxUcBn
r6cgweFON3ovyqI0hw2kqn2uPFIqww3NWtxuWuBDe8vTTnh7wzi7Y8W8pPYtxCpOmC2s8AiB3dqH
P8iDtx6xrADaGAMNjWwcZ2GyOnD4w/wFrpmeFlvr1q0lCaTIYSNTgFeV/Pql5kdOIaZCsp2Ji2wX
b+FfNP4Fzw1m13D+L5xXlAZ7PLxq4aAAEMjv6w2ToDWBuz/1LKfzvSvvfnBjSBOav/b1FSDSWBMB
0LLJ3oHgZOsiZ4h/FBqnBJzpUt/RllPcla/9Xc8L2bnz4Ig3Wycvtoa+7GfAos6oPtDMxYGaTWsI
3EXJMzTTQ7H4zyK0Ly9ojjU6QMo1CX8uzUTv10GulxizTqcimVP6IjKx9p7BfZtpLP0KiDMgoft2
0rHcyUySUStplyvqRBlXlrda/jvWuW6458pAZu/yz+S3Wia3+fHlGgJCqaC6v6aOHxz3s6Su/00w
TTPPNl2LDPbcOyyW3QC9qrqJbcbXNBHGFn0tq5JdlTUBudEWkfBdYu0RbeQeYnoF4bNeq/5iqYm2
19SvXCxu9LmvaCMnpy+uaI8xL9rLCQ2Wk0nzYSLBPvC72d0vbBV+ex5DkXoaXeKAAVctdQI4jdan
mG5IDJHftKe0dkxs0Sc/HbG7TEQyu5vr+IiW7yPw/e9Y9/G6hovdMoM9rKkvXPWEOjrRUqQybmVJ
KXnJ/Ci+rT4ZGmWSgcw4g9Cg8Podug7VqeEwcl19jOwr26qYAJK27WU4doWmmpHPVBHd6Beltced
Bi3ESwL7Fuf3zi4HEiCxYrkLj19+/7yJzFmMZbWsCCs3NvdlaVJHf1lrydSDCDM4oD48jLQUZPf+
F2bOJQBSIRUJTBeNR4c0ICiaxMJ4DacU7iUFte2Ixp22KrMJ7ZiBYj1Y7qbC7cz1+VZQDVQWUOLw
6NI09SXDcgCJxCCl9ach9pbTx5iioMINq5mYmRNRqeW39H2q9RYDoB3RTFV64/4cu+o1fcBPRICw
6lItdyLfSzaWATpS63j8OUq7J71IbEg0R7oOdq9JGu5ym1UQba5YrsXFkr3zTlX6kUskEW1aJPqg
DUvSrJ+jbbmU8+ffjvvNcYrKVcoIzxY0AjBszVB+SkwBi/nzMp5g46CxFRGpfc+QDX9+UcAPteT6
SUmPcVz7P8W5uW0XZ6bmpFHrffv1EsuEU/zav4ywmNBlXVBzY0sE/cIQqv9gFkI4/Y2yfI7PBoxH
b9k9gAjWS1hN46Q6wsqLR6rv/EB4NLx2rQ24ZpCgfK1MyfhKRDervr0ApTGXrDoB2gut0YMt1CtH
aBtlse8mvrY69pmSIUEgq68VxU+s1PcEOrKuk0V8Jp/yVC20dvdmuNzbBRD2gsekflcW90Ldp16R
TG2/P4x6Xt2/HiGpjd+xTMBdbd/8zl7iH796oox/O45Z18RO9HATZkSTd0tqMnZP0dPVQPKAxkyP
St+7dT6gtARViWwNmAlkLbX3ua4oajPFkEG4YjC659UnMcWo0xIxxT+zFQVa25sjcdGIQahZF8Fh
i04V6d4w3mWySul0k8AR+YTqFHPtMkFPXqZGi4ZlM1SXJgZchWPUc1Ph9Cz028NeHM8Xba6RzbgD
XSc6dvLaeAd1hW0SprSUGvnSeod8glx0ebomZUrslO3GxFnv9Z3qm5dhGrBPYPh0Rx8wdO5NURzy
MVTgJrKoIOKyRCSQUJZHRnCP0gvWn0M04prvNQXjFc8yCKlq2aAlC0iZiG5beHAVbRZDhYFREkth
YfEFAgQMdrTfPlZ0HU6qDEhXuT89msMZbvWYNDtVJVph5QkyOo1pCVX4AMOCz2fGYIQ9puXZJ7Sg
vFxS7RxaiXk6iS4kKg8yz65Cpr/BS5T6WOSTEfL6zqPv6UccoQIP3TAw73Y1UelXYy37tKCb//1C
HauxC8UHTp2hW07MCKXKPhpB8nmD3zK6z8d46qWO7C4ARjcFkHRce7QN72V7dPJML89YR7+ihEBz
oQDv0o2Mirx5HnB1hIxcUzDy0WPK/14DHdFvwgbIzps0Lxga1ft0rWMYvV/GjK0p6Jlkv2zfcYWq
BpFaPyKKvFuu3N58hlQKL0GRyJ3BYRxlpwi+FaqGlqhJUv352Pu1IWe6S1+bnJVQs0G5iUIgc76D
xT5Uw+g605PNfjgeNujh2AH5MiHlzGYqaNocU3fEUuI8jCRK1xfW7FoGSaq+9NrWOdHWFDmGYHmP
RQbawNvkV0KB/uqFxFw3ZFl0L3XwwfhsGc34HlmAhtvHnf/p7XVAF7bfbLpVoNXB8FD2lfmG8NRw
c6Jmllp3gVzXqLzpHlMjflLMHZrU4XOjsB7m4NIiGZX/Ape2vIslvyb+IjNbFuIFnZPN3XQwfw8T
wkUeSPYbPJajs8i6X81ywqRukj9vkdHSTybvcskUNq9SKyAEZRAidn9O8PSIE9qiqlOg1iOBvfS0
lDcRCD+9yuVjtmJhohlMbonDhwP0XiBC3O57qMZbB4KEtTXn8iYpepABNuJ9WeStSodBdg40qCQG
7HFgrOO0ksW3UALKi4ezRGq8gIiA9nupYBjg880jFhl1xCIiFxxIGAj75Y/Wu+q19w/A1mTptxx3
vP2SuC9WppqjhajnHDsETbPZTmdXrtGisNHnhxHoHVDvN5goBdvMBbQvkYtCpFAeCQP+VFMj+SaJ
00mvKYWbH148Pl40AX4pknQvDrCCrGkdGXS0xg5kJmhc8omvgdvHT1VzDIAh6eatU1wUqU5ibUn+
27cXRUSY1HZ8hEExgxBT2Dp/upzwd0rsYoTvgt9CbScgjgG2VV7XWDtsfweCCCilT6UJhlCmoIru
pcg5nFGAdf0vM2gpntGESIxrgqZdt7YuiGuWE/TUkqe816LV6Ts0N4GE9Ek8anmmtbmDyDygYgYa
c5K0OfKqnxSWlVVeybsEa0YF3baGncN74qjIV3lsd5eR5te6UvNKzPKtfGPzvEPnC+c06maDeRsj
hrDmVSrSBAZm3LEQfV9SEA7XUFQHJ4ic1H3SSo+cKIVSEihPewH7wX905QoZ6G/7W4bTXWQ192ez
7DPjfoh4cWvFYms6JhNGTugDpE4vUPnkLHsMKme/MaudLnTSh7HQrutWwFoE/gsPJxll+H06o04O
xkalV1fYsmd+UQveFQ/jxN+Kvl4PCK7svGQwYAHAgG1R+bEQQ8vpGupdwber9PmaN9LmcaV2K5+u
io6yBkb8NUenrWBHQzzKTOcFljtqswmPi09qCLzU4IIX8PWfXvl6LmMnwQPKzlvhZoMcXiFF+ohm
c5z2fwc5lph2ykcbilwGoPUU4tf3JQPWUO3YC7YZvco57dKKIFGSzpRi3HuHp7AAcI8jDdZlvTfM
CV0SQr26clsPuK4SHFNC+eZMh8kvzGS+fXkniRuZr5NLvj1qMOxytcYMKPJ75lxKWrKqzIllBikM
Dyg/eOWk1pImCvlv5ubtTMc7VKKn/V7SSXyZ6Smth7fMbbViUY2pI9PXZiwM0+jLadk8kmKz2sbC
h7M/PJaZLgsOWYnYYejm4yjPlYUZyXO6QgM15kq0CbsD0PQ8dwCK11AGEWpH4dazcWpT6e9W0RcQ
MHltA8KZg7nppvNNDuxZ63HrPJQMITfMPIZdEXsxgU97M71flzOGVYXSFiyLwBB73aFshaeDrMlO
cSZin1Cp2YybbjGmi/n6I/6e+CMFhH+6rrwKGBTNH/I0ze43N3mGBSctAiAvJMnwH45jKYxubLDu
vd0iI9Ru1qLpiurTw3tMkZgwgbBHW07XvsKMsbmt22sSiipnhSNSAFXPbPINjCwvxsp0VD1vBBpK
x62IN39fuv5uyrOcb/Fsbav1GgGvm2saepbOvKptBK/zVhRhar7oXmaJk/qK11ZiJIXfHChplK5k
DoPFUCLoPa9hYdtykd3oOgooN7229v+cF7+3iZJxcCd89xaikIyTa8GGIfjCS1meVYOUBEEzJ+6M
TGSsm0rjt3izxT/KcwMd7u8A2stpwjG7T3JpS0R8I8ccnNiz86l+42nXfa/5s5nVPKC1RN2RHIpl
ekqHg6MTuX931xJUEcnahp1GMoikE4nnOtLPydXZNZ/CcAaCP64MUkVaSryMU1PPoVzj1HMX+s5W
2DbeEwosElbLYv3u7TuFTsoDH/zbJuGPwubZsOMdIxROxxW+b7s7ET8dxrl4yOhUVxZyq8sZ5QVl
fdDgcKgZq60MHfFITUPVPf+h8Y123CFNxWhb87EN0zlkuftsBzBBvwHc3garGTAbm/IqYr6dqlsL
8Lz9JRUN9MftgaRMAq0uQ9qfH94CwvXkgO+AFK7VmwlBSUYrrIEQEfqGeY9v67JwAL2bFwVsTrdy
mohMKdw6MjunAE8YnLTeNpM60zSjwF9ztFglaN57DL3lcPNhyx/5KOYNP7k3FEI1xyBpShCWAkx+
awrXPmN3gF6zQ6EO6yopcAbAa3T9cZ+AKyCAq2DiUanAEWyITnoRdYSOigjJqSvrMPpy8Z4lwR/7
ObWwIvdDqHWRMI9Yd3xsSyOslu2Jww5Gf4/e2DtbF1r+eUXMb6vFqwthWS+LyXEOKDOFSte2Yibg
xVfuBxesPRqRJxZVNUZ3FSJCvkyPyRfmt5SF+/K/5h6IDej48kuT+zSE4NntgVgmAbJ6oJfdX9oN
+h8C911QZTrKmHjVde/jXkSmkmtAekwrX0jtd2ugI9EX2ZBqzKXpXlG9YiOq7EVFiHifIDfrasYZ
qLH2js5I4f6xmnIeBQI3VUF9agmwd0CqrEtVAOj6ANvi1Ycoc8OePK36/KY923Fvqkw1GG+xe8oy
FsZRoQhMQNbSVTqQVLt1Ab5zeJl1xXP/c6JThxCs/ReGikXOVoRM6N9Zgg4Uu82grmKQRrSzE0XS
lhe1AWRfoOBjJHqzpua+Dy2USAtjIA3Irw4Ob5pcm5Llg5EPBLhOGtm+c6yBxY50J/nt21JPC7m+
92mH5Q01OYh4I3QiFAmDTVsOISRaVH2uO3eb5iY3beQ9NN0bnScaHWfYS8iREfoe+6n6FPzxYFpm
yE4mFcTi6MGodEsxWmjPWaoel8RyMXZaCbSSA3GusprRj5fIq3OCrawYBqn5YCK8JhYDwYsYla4M
9tNFlgXGIsqHzgZMPa/i7Fs6Iz8yVGmYBGYmLVPQMFzXRSYNzJyCZR4wRo34fFSbW45cHD1iVQo9
vmjcACQwFrPZyXhkw2Bp0yDPI9a6/d1u20SRgGe4+eyxX6Cg9EhIRVyIb8QIMDW3yW+N07t6H8dO
NBe+QKIQQdyc1/697+xlZnhg3pMhuoIQ/aWBlHZX1jNKbfew4gKWuvgCZ+uSVQ3R0HmXBdex10X4
AmuWTItcYUiIcUiJ5oF5i/ta5cLix9QjlSXqYPJei2wv2uxTo3qEwLCHyDmN/sFtEYFw3DfJ5cYp
YLlF9TD/z5DCfD/bZe5OyA3JYTbDLCMxwLwW3lSEVqdQzkGLCl5vv+oPDK6QU0gasAAXguyEgqsg
IqGF721Oy27l9GyE+BChQWxlmwfy9epNoCuNBPHPm+JTTvTFdl+vjQRNB1Ig+k/OGUJhEr1UNxQp
GbikyiALYeed45un7/qTOOJlJ78f+Gg/Lz2VI1zfruBTCdxSEVz2/rKCBDFHZX/KrkMcvvETvGm5
T1XeuSymGlmRvf5G1/eFINWSc596XB94Ddga7/R6cFqzxwLmGT0/yfaVASSzw/HHG3SnaQNwrroA
pTFOvdXYfiVec240spUYNHqvl+NDVdYmm+WCI938f5wSTklYOeEURU3dn3KQ0GmvbPj3SQpCsXOA
Yim64D+mG8gGOkYmqEtNqyvAdHIv+MIwPO/XD9NEd/SiZeNmHzpuwaBtDGgKtkoF8w4MzyzeNnQJ
f8t/J0lXcx0dAqELDyN2ESxCoaevE/josX/OiZODTRTTg4u3O1PYXPEQK2cBm6oVlv+jXGD82QY5
KjP0k/R4fzx0mWfxzFFbJcvTHhoteZGeinGQzgfXlIm+bsmgChcwmudhsP9UWTk+a5z5fU9i6AsH
IyfuYuA4yqdW6HdD3RB5sSM45O4I56r2vRsw8eE8Kz0uU19gklTkzRXtUdupopv2pnBHttUpv07B
yqr0t5gAHwdFEB7IrzIWRELcW8cBmOovIAxTkU8+Iu4+Ml3ekxGaPdSZwHj182YLx/Oh0xfE8ig4
2epHHXO46+k5aABP9SpjVTNLTs3sj2AahCGi4YZWY+/Wr2Y/a4dRtGNF7EmJ7G0ltXdDlsJ2yRVm
Mn/9718e9s/PTQdUkRAKxMgUaZDCc2fJwNpmU3P+W/M8kcpEMdvfHwFA+zV+Xl2WjWwzBMYQDpte
ESN+ChfvYYwzYonImgUUzHUrnlRViwlz3ul5/bADlpUA5SQwj6Mddhdo9ruN2ZLxMK8oS6+HnLrS
WYutlb7Ka0ATFpxeqhXytIY+W5ITGwg2IDHldJFbMabPEW9x4lVx4J1jp1u/PePxw9NOR1us5BEl
bC8hHlbNaVQIlr1GVwa0ILehWKcFccC+orgpctFxD8M+pXpEJLgk6ZGLM6a2QqXKqEzhLRZEs0pO
iKqBbGcOUob32B8CrQweJPe3qQOXyBdBe/FAgpCPxMDf3iuTfk+vM+Vj7uCKDy7jVqT72abtBgH1
FT+RTzh+gBXYyX4s93XIa9Nq/mHRieL1aEk51Gh/8GW3fQOp9Oe7MdEdjQs6ZWPJX9jJeeRn3xc2
QXUsKiakchWCMpm2Y+jIH+U3DtxJkcffzFk3hDz62YO9xMu8JSku+p0zvSs54y48cyc1r0xzOtyQ
y+r3uLB13I9VR5FensHudQcnFHuZSvSsIkt2WAN6mIHu0pefOm85SxQN2+TFAoOGQlVvIP0Z4BuN
Z0dsS0pQtXX1NEHkTqmS+kDN+f4PEGFD0KveP7VrP9NXUFv/rC7X6d4CFgN0X5rlTm+p9Du8zyDW
/VhEtsMKWJq5X85AOllcFyndSWbrnVtNkSjET0Lro8dz5CnCF1+CoX64deXotDAQF5c/uq96NxWZ
annQtXz+viUb9ag4gFE1XcbClYZ5Bqsh1oK08CQEXNfbBsMC69S7DeIVNmdworBdGLuNurarp7cn
AzFPv38CqA5+LCiQ/iwmPlFyOHcFWVwQ6WjbjntKBgMQEYce4N41ho38k0IOP9A58y15EBMavPsG
W5HVKUik4o9W73LVo/uozL1eqhA7OcpIUbHEThuXvfS7O1RPIfAuLmwP/2C9sN146cn6Z5bsRs5T
tYVZalsl/qtZKKdLqC1OmEdPxnBBayymkuIUbjg7WA1wP65zEmHlNmvkUkKsPot4akRYFqb3HhYL
zuLPzkfGKk15acIcpBSh3oNacxotZwgnYVMSoZWqvlj4jQcvwFcVQug1I91uV048cwb9n0/05Imy
XBvY9BBaaahlxprl+lPDhjwU2NBGGN+bcBq8TcO9swhDa0Cx5xNHqyFfkjGpsszqrHPIl25ieI3G
XiMp5J/lCApKyiMf3VNIU3oRQnxhXKxyCTn3uuVRz73QsY53VzwYC2Unz5Q3j76TduTcR7TwgdD0
lF44NBCvsjMoZKnrabZYffV9qMIKhlwNqVIeWW5kC6CoKfHg37H+UoDmecWP4qKyVkcox5lfNYIT
eYUQrs2czsH0LOLLu6hNqEZwr10WuNbFNFH0i7DaHdiLhegMtAUOPlQlj/7w7pgHZP3g7vpK0yWt
X4z9x1+uQfdxgVjQv7yrT7Wlz5cujLxJ7RkOx0aEV4HG8kHGNa3p2GKUvLIIs/DOvDBs6FByBKO8
Q9VgsIm2mEQVRp+8zyQ1LbWnNkT703QK0iICarXdqyWJWk3vvwNP62SuXPsPqIqbBXC0VMzv0yL4
RdxMW+diXddUZKpW8adG93kEz/pvwTf7Fqoikbx7YOIz1P5mZze+9Ad84rem43P5TmcT1ERl9STS
8ksWYgDgiCu8uE5xHIOLffz9zT+I3J9ZZfFqrgltTiScIEq3CEEwaZQRE4zoyul22xOniuwD6xIB
BdUEBpTo+DIRpsZiiXjecfZqEDWiWQET4xUR6pGYOw1UHLp9Tk+ByYcEjdRDgRb7RrEISukXsga5
CpIADy9+Hs/LpOsA7fKrL/6qQ79cNU96vzNVTsWbqK+wIlzlqENZj77BkFLruQorBUvvi7wEGSlh
rENMrvsdzoHSjmg2QYY9NanO773kRSlACqwh3uq8XCQzWdN2EUNOVfBXSe+nzlhyAvlywc2tPVBn
mFTVhbn/glPo/LoyRvks5Pd+Szf73Twvw/muHg0Y5pL2QLWzvLMYSisWOng4l7CJYJxij56dnsRO
v77CMmzaUnJehdkTb+J+F0iNKNOPFfL+yikRwJr+4YmZLjDr8pfWnRjePlVDUuBxJcTzJxQSTfuj
Veh97X0T9BWIPbCl7lspZUTFWhYvDpAt5kvTAwb7FaL5PSjkPQPmrVOtbCKPU5xotmFaGsaCHPKQ
AJdLhFnmN9TvWLO0LjLFj+zAUrk57XP7uPKUiXd3QRW+c/zuO/sh3kz5OzagkqP3HTRKXI8n4Dn9
iZzT1dZSHglzn0iR/agqQwSn7FFfTJ6JkpVU0VyT3lk0OF+s9epi51TN9UWfVKZqKuFSTp5ckr7X
fQdOyBK956kAwBws9Muiz8hvFgmUcEKC7zFbtymSk8WgLxX7jcGfiT00YJwHiw1fsHg6SEf99gmu
JIq3fAVUhsG7g/4Ozywoy2fwysV+ipOj/atxpkXKkPqOFLWKDGq3gGgrLqk3WU2awYzl6DZN8RoM
yaEOd5dtmfPeUipjqihdaDnAAZpO64gWhCDa46gCur00RAXx6ufN//le70iMAeFU2MRpgtHWUiyL
jILRff3w71F8TtNoHAcFlSRj3RzqjxrkHwFw/4prVyAMlYh62uozqMw6n6iEJJB80qTTBYJ0zkRx
yskVtpAnHB71MrqpJ05rMWx9MGtcBnzPJh9T6ei709Jdqhlnzr0B8OrKICJs0CK3mYpYz/Vd0Q1P
bfjHw3hO5Fmxln9lFwBxXkmI44M8wSEPLg4TYGmgApUt4w+BPWLH/8aEAazD1ESE/xERBcnn5ZtD
c3JZhhDizXcPKXF7lhuIvAeMf8mRvHigMwmK78OWVWfAWBKCxcHkCHfTvS4etjK+GQ/9uvAgu1RI
EBDZgnhXhzzUBNNkG/3O22KG8YcN7OrV+bSUWMMDmS8WP1Zy432E0lDwL8swQhSsSL9ENpdmqh+P
3zRImSv0J5A1RiovBinh8hVCVcABlnjmc2eD2qIXhILKJj3jFyGibrEU4vaQFY00iI379xjztwen
/ve6ho2cVEqN5SmUTDCosAsVF2y5xmqDoLL4Uof4a4XfSbrsGl58czBEdCfxuR1Ng97EhSu6iC4H
H2kcpIvz/cum1UZ+3YorVpOCduLJ429uzpreWiFEykzdUfLb+xVmqHvo5i4l7oNHs0ZScSTdA+Bn
MzXUjws8DplzqdRXGylQC/fXUY9fZt/rJjB24r4iONHrjmv5WZNpD0H2tuJXWDRqTCr+NRTFzz58
Ro4Q7wEWqTB8lA7Cz7w64U9398ZQLHWvKVG53KI3KQGZEflu9UTHh91PixpcE/Q3Id0S+B4dKKP8
c7DrTFkusnQ9JcXsTqcMvIj6qEXOeg15zkCA3w6CJxvoHn6w7GuoG0THTmii5+zNfVSiTDJy7nHO
U6NwUi34RDqIfFLaCRM/KQXzb144eh/+1KqqAoNArhF1UOfk8iE7+V7kJzOZrhA1HmCkTVWF835S
hbHWP8vuUpCnTb6Y0umehyTybH5uS4T/SJI99ADq45auPS3WljMDiukUO2CaQbwh7W9o2eyYtltl
hb1z8yLRHSRyOuwNmnx1IVELSjloNKXJ2gRSBNpRxBsAMDQyePF4+BALRER/ymyccrZl2MeLB5xn
LjL+SeecvZYKu8wK0kxdCVm85wtbqtyjh1gNv4KdIS28xAl56lVUb/gPv93+ZEItUgGzdpd7NrJ0
w988Klk7zQSelNTcG9jbg/DF3HtzkyzsobZivE8Mvjg8hxWz0pg023BCjBWPOGU1EBdLsVNPCV4y
fT7RAM8aOkQidD/f74oaYh+ix1g9Z+AXbnWzuXARwToU+XV23TUH7qefhdFSwLHiJXKthtgvJaNr
V1a/45JAMusbefMy31sLyrYkDyVJRwK0ch0E1/O8FwzcGhEAwLGfZ9XmzXQjPqJxNSQzYSct2zsZ
gJj5D4jBPtsxLgCzpbGUbEmPO9ddAmdpjkIDjm7sdS/cGUgHe2oTzwM9LegXRjBhKBo+6yUnjx5t
YMmN/mO8lSihXSSQvWgEwbb/GQ51f9Mx4AV1c6HQbtz7XZmm8JmWpn+CesEgGmGyOV58i5jt8SGc
zV4wNPVx0SLACnN0MGOiz3YC1mD/t3wPTLExFKBVPqw7An6U6wHK0SytzRZpFotG7eRHA/EdBVUn
ZDkpP+DAF1+mTJJC628SArB/fqDOj+mlv13o+GcHqyXGEtzuci7fEsqRNOeR+Qd91aichtQpdtW6
1PyL8Tt8j8gsxn9vqPEOceYM+mjbpqXBFRD0oxe/sMmFAwpcdnXk2JnukESTE+LimzntUlKpJH2q
e+3Y+4xi7rhVcuieGOQz5P9iVysT7H27xnKteLm0oKRXjWT82wDwetZs+PZlNRYvUyBxbkArtn/f
jhmoBl01rLDW8u2wgPe/FaQDtPOQ4w2jrbtxybEQGshgNJwxMqAiJUcgo4zgfYeSv1d/H49kAd7s
//Y2bDeDFytup2yE6zyg6u8RaOTshNVIJxMd8fSoOwAk57oxxdrCTWUrZlMXA0amoYroRmfqAJlf
7slzc7bE1HhRjlpDJPQm+/GBo9WJF+wieFdfUpf+kj3QDmVZc3sabyUcjE8sc+s6GzvSSTsQ9DN0
C1vK4KBKT7RGVNb/h5huEmhPXYvRFRjmPg5fk6uzYawf8H9p/uf8n6ytsG/DtSsXLzS+KduNGiB/
8rrGVCHNP9hj6ofAL/76XzbY8SPerkfmcBLaPVJee0HQVk5HoLtfqh+m0M8OwVVOYEy4u1yi2yNI
SEMR97znjWzFpkqlV9Y3FSCoC4QjN7OFZ9Zx0zAO0fyDvIJ+TOqIi/gs5IIikcgzSdQjQegiJlig
2clU00GZbAbAlRQrymJwu3YOT3Ehoe9YBlN95X0SlBCBlpPQezCGsRZc26SVaBgjK1a97nqeT0r1
gijh3caFYUumIjPniB7ZMNofZE7i3qEvvX8iCicSE09TirrKnGrJjWXzI4JmXWrQu5xMpcuuXnCp
rJIDz9aNffncltFflNFD8P0zF6D/8246Dr7eGwc73E4iH2JeIJXobZsdTgXnkbrWUY5UqSQln3O6
2l0bdc50ZVAXpRNwJm7j4AFwjhwQT+BrutaLi7ig70cfcggEnHXbxHtyoNyWstv2p7gYJ94MVSl6
qcEVFw42X+IVgmo92CcfHZksII1tk00U7E0IruALgC12NfrGC6yYflEBld9o1tuFRABtM97psbKZ
8l23XvM5/OQ0FhngfqolDBWgNda9v9ps/+eXAmgnegVXc/HPYNljDqPkF0wf26rJ90wWR5bxHxiI
d8mAX/zYnHVVoX0k8VEq1nnuhs0IqfGvr2JfBHogD7O4ItEHYumHd/Gqpoit+oQGq1AlkqkljORM
MaZBxDxV2OjB5J/C9EFBZPpWvC73R936b7exloWKVbFJhexk/k8NSGeCJqZrRTpVkGoZl4SYBlO0
XUD5cXxciI2XVi+WVSAdPkPf2Edds+EKXp7aYdcw6N11LT66aXjUd0NOung9iQxXjdgjoSV3LJdm
GutZhzVVWSjksFYGYxhvnn/qMxHMCW1mxoFFZxHBXejVd520BPllHW4qX0KpwhsUM4y8JTiQVWeu
oSCeY7C9tuARhZe0GPEscaWHeawFqW4bd4qbQKrqgF9q5Lo+aDcEt5mPotnGtzhYhYTwa1UJQ1GB
nsUBsLFJQAg9pUKY4HptDuv606PgI9FUsMxgZAYaXnLTVGAPMzc0L8+B6ZYDnql9RaJfOTX9gtYT
eHJ8ChL7bndQ9Dc7zBIL9n1ZOGDAs8uWzfOnNjK7sot1yOZHMl7t2Mhp98UlHNqWk9VF7Vhur97p
t9EChTb+KA5TLQjcsgbo3j1vS7FpW9dhrxKE7DuTIHZ+rWgua3/lf5bK7UojU8EqZBYU/Z6N89ua
WqWPRCNp7muq9e/JarYqa2MyH+F0iCpBYjoUe3lAtHDQ1GPaMeB9L5R+1Oy6fyeybJNTh2fCe23v
bGqy31mCfUkvsL+lCgmlP0S6HLqf8FSquBhDNn7mmrzjEjE73v/5t19DZ81BuEO6j9UcA04MwYMJ
rmHmRGqpugAOAaFAYHiZ/E+ALbetvdr+BzxO73Oct1uJfXqf3NOMa3o+ThohpM4+wrKJ1jU+JXtc
VLjs/1XqB3TvyMNTJiE0431LsX0qajHjfjMKXKt6UUAE99hiWZHDqre3uynGoX1+GxE+natIqSPj
nKYFwK5LLIdt+LnVplZ+xxMYvEpuY1BJXu3b1WWahLrLhTFhy8ppuz2khmshBDlawLppqPQiYpxv
N839YKc5DHcixX7To2PHTk0ObDtfsFIXzuih1CQyR/JBPYgxNQpgzYmx08gwP5821nr7mizBmhq1
RJ2cd1aPV3VxaScUxLzVkEDRPsWt6nPB5WQvQ8M8wy2thvUJxgJgXeOEib563bJgFPCnoJJ+jAmm
jlaEakIGWXho26iboCwcw4TlvnzLpSUpcr61VKuMct+5vmaqtkY/Y/92+iANlFcZNfrhUkSjScTb
xY5nKCKnu08aWNM7U7ykW5HhgtHXr0Lfanfulq0sjGnurRX2mZLebLo0QydAIEYf4Ku1VWxnbvP6
tQVa8hOdVamaz6sDUJ6EYpyv835BWgaJLhkiGXlL621JDGkrY6om/k3yAxOfPAEqkxWeLALl+3r1
brS4SGrmdklLP76qLFdscxqKFpmxFz62++eXD4Q1jP/cvu2EE32jGh8vmDkxSlIi5FttuLjsmU+R
vlzHBjlykV3Dk2ecxW4Sc0c8d0lOZ0PfdBPWs6J5bPJCXI/mkmNzlWo+VLXLRB/qCLhSNMKez5IH
NEmnSRXdjD44ua4McdC87iLmPfWinYq5vXjFg3/fAkuzmwRUeE7cMpLeb1Ip2eFWUo+BnwGTsa+D
u7fuRA5DE4J0grycJVsChhMTzJXCPCgGjGrkOr7Zb5pB+ACwNTeoS2x6BgoM5SbRpe87J0Vifs9a
AEPxy/ZkCxDLXrka5GF5JT3lqlnU5WkIjL7P1QEHDLAuh11xgyDEwjn8ixgh217t/2qyiquNWU9w
8HHiKGobJjgRLt6A5SzBEX9cDZjmCzABae94nLW8V3LlAqEi63bRnW5e91AkrayBTmNmRoqlqzKg
8HDxw+pDBn3s2Pr3GG8xRn1I+wKqsGF+dbY9ghzSFjXAFdVPr3mOtnEjYvWelj96Bh6GqV0Md6y8
3PlJkeezYK39qgP/EPv/DR1w5hQWtViEzb83Cu0pEpdAGAfeoAtJR3Sy5IIrXlaM+owztyf6IK6x
IaBNlcLPrJ4mxg1dTPL8OM9JaGsii3o7q+4NtPYARjWQFKfVRc6lgpuJgaUcer7znSYh8I48O9jC
kqjvrHmHHzasMxtZoQxHQ/r5hzQSjGOjWbxEpyky901GM+3mmmlA7xfToZ8y6YeNRA8kKd6E7jxe
9sdOxb0GafrTIzznUgtC8EB2ks00FO+rstHIZ+PQ92itERklqdSuEpWzk6SPteiqg8rjJT7CJ8v2
jsXaxeZny15Wg7f+0/g5jZdfieJY5jNuQhxkf0srcqKXCtZ3tWNxQFh5i7pXtXlbva9pDMtGAbEP
erf5E+EGs7TgJDxDObXX/zwhm9y/gXt7rEYxKyXqEcRsC4+uHiA3fvavIbOvI10A5z932eBawIJZ
Sp+c/rrc51AMzNVrFOQ+Vda9hgig4yFvYXR1gMjKbrIZgj40kryhea3tRvbnyyIzzED4pCU1RdtV
ijszpCM0mhdVMl91vbx3zM0F5yKnr1W2z7mLTj3OXxW5eDMrD9vrQUELIPG1c5fDPUIHkCNJtX9E
/31EHbznf/GnsA7Kzh0NK0g6V+vXvMw5ak9lInQy9wZn4g6zNa+4RkqQN/hAuS1WdESoz57X+Dqk
4iuMKR/RwsMpl69YEpxcgKzI2rKLVxz4tRVlBcNNn2CsfzwWP5TLfVQUj9pbKCjAKzQk+aPXXppE
H4J1TCsJwZH9OaOoISUCXRzte+IfYiayk4ZMaUBOfwxEzyxI8ivy+Sfjwe1NogZmC6pczVzHCe8W
8vtDm2aCRbwZ8w+uQHaLq2Fz0SM7TiHdhCagGCBZF0RvnsjlRBQPP6XSgY4p9vx6O6+56KJolF6v
QAKrQTBKfwtD3kpkHIWapaSUhepWjTi1VxsjfaAlPEA0l1+1qbrrCTl0JLxaJwPPc6eIEeVWkVgN
ZCqAyht9Nj8kre/VrGTDobPabrZCa9PD8W6jiTe1LUJS8jx35PnguTohlki8/qHgCK8Ql6itPlQ+
GN8uGF3DWxUSWHy8js9cbrdgmgTi6j20YQtUI8QcwDo6j7xPRpOgGs9pQLWocgeqSxNlL0GAMueT
0y3a2/aNUoVusFpBtA0K6dr73Q8UJg9C1RuGdnKMvXmV+QpRTy49CJ4XVk0Ul6e2SpNsy9fsszFe
+s/7ytLcw8grmVs3b449LE6w0XjrLoAd9VbBUkPUhK7BDsV4ZDO4u9D+7ZyC2xcSHOTKw1esOOQl
MIr8edoqAiXY/PJEdr7v3vvfQu2xVkjTlGzQPHlmJblwEoimieaXSvxcOyZZeDWZj2bJsp3nv51u
DM+X86UcNUJBsfX2PcmTPt5rMM46+SxLkU/yBqRH9Uv0WLIBrd/i+LFk2eWhFPtZfAN1rcDIkeem
AvanncdHLLOx5bpyoOkwqa/BPdEnpOveminM6GA5vhH91ASYrr0FrQjQ3SL2IY3QTPGmQdzrK2Ql
ZIJG2ntrBdUmmHGPRGR08ell91E1oFN1eMNlMR2ZZIpLEcP+jfUD5dn6rev9j7NN0qctRxChI3XV
mJWVGFTVoEtg4GMwaKtQfrs3FWUsfsGqWfw5BlwLHGgV0qyqbGPb+1dUz3ozrwLFTZCgKIp0eLu6
CMepkSETh0WD/hQeEs/qz0JG+k/MmPq5+0HjoWHInZm+1NYXvY0Eid8nNOaimQCTus7EuZpot4HN
FKfU/6Gt4gnPgwDG+IttQGkjHrpkEOrpzZMUhDU5cKr9acEBRJYdFklxqkoClC9bcNP3HKFWi4QU
EHjwBKKdIvhw7fAF3KUxrkGkiJyvO82ADS2qh6osg3fPSqoyZCbckG8A4rAuEXP6fM6/UNBWyGir
9pQX0yN+SFzT2X7sKGslvKQcqxC//RtaB8dWk/1t3M+vqbAReIHsPdYHLZ0szYjeYKc+JeNFMWCi
HnhqjoPGa+QNgxhxoFg8/2YoH9lcZ/SOIRZrjT1DWd1HUOg5MbDV7eacFz3R8uqIvSljqJiyex1G
zMxSCDTLimpnIFxFqz3eGdSy4/YacdcodqtF/LOOn0BXrTev0PREh/+qLNFfPgvhJjOgnv0i8M5r
3ikoAryQrTN7aUfxrkTA6VXajH3jV7SAhP/wwRwRzqXuND5+bkcSmTooLrWKicqaA6SJZu39tb9B
zxUAv9EyvZ+uDcLr+kTVLaAHZ3NjkhqRO8t8HicFJiFZG6PU+R2/MnlhjoxpkP/cRa/5P9daArWj
dKzEMkXg6HGM1VanIMU/ah+NgtMctE1FWsE7feklZAfEcDY+rHLgOv/Mp1fNbpYU16gtEjuTETDD
YdmIFcsls77jxVGwaebRo/0X8x4ARKatd3+POROQblnAecwH6qmQ2thZVGhgSqUXvQPU/nRKJiFM
sAarjSIrL5XoTYCa+8xp1+AOjc4btdes0HoqnM7WN5TrRdvMXI9klzUbmO8YvraWffAOs6yu3RsL
FxvxWN/8jFabTcODEEdd/dNbrr4R3WI54Cb6uqq6hR36GvrS3jbmAx2ezrQUqBy0dexNOsKdzABW
ECJoZ+lX8gknTFielVSlgByytBl7ZH3dCrW0XFAHqDcqcAACNdC73MfeLfQ6MVR8nY0R2hta2oJ6
CqcvZKdH92xhBRcdnayXluO+WLwQswoWABVviQqRATAJyBqOZ4gMu+YKgcltfHtDX1oNEUE5akDa
L87QX1nENnOwD84CBErSiyiTBc98s6+ZvmP9px+Nm9Poz63st4bL0IvFd71soRUlCZyK/CSFBBNb
iwOJmxaYppSXdYcLogd7EiEP6UKkv7FgjHwgCwXfAdMqoXhRTopQtXBipHE2U8KQoc640F88T6gU
9oTCJ7J9aGwUELpktSVO7SY33cZxmCivYHo57UY2soSyQ/nIYeZV0DX5qntb+s4aS7YPJB2NRNU4
6+W0IcU66KFaab4fhMkncMsD5U3C9H8L5alNZGTOtqN6s5Pvq+Yr8XOgMP4k4kI8ohax7GvqyC0y
wfwl5t4/wOrI0CPx7ykwJxKDeaG8Ucmm5dfnQkOnjXl6tRXKixHP4nzfS7w/SZvsQ0LmRJhPnuRp
S6HMWe8IoMOsUs0xDqqmSyxbAka9TgA0rKR93TkIx4BrBJhwVpRjPbmIBffEf+I+v6xSB5/krPuj
4jlayp2bVxmt7wfYUJccjw/+N4RuC3i33HzZzHZupN+KsdVZ6QhDBVWXFXIb3eGZPeXlSo2OG4Fw
ICIx8t51uWpLpwKlCS2ZKL8T5sdY/iNlKIXfUrNdYbI3w6ckru8OeFu7WVy+R9/GkAvN7YkyOSSU
2GH3Gd1o/e88FrLwFGpnjPJ9SOuro6nBlqwqpA4o4WoeKtgKTFpp9JRgrb9tVBry8rw8V2gBQibN
96Qzwhu87M2K47sssdeeU6ONqXHJ0FSTBTWFK7v37aXMrxJ32xCXTp91C74LNa0+K5WOtpJrYGwg
JxCmoCy0u4ZJ2up/jWIMoFwkXJvk2W6ot/iwb81oZkdgTkaYGi5OPyFHGiwD0pFL18ObhY7xeQnZ
mUESB0o3WYbA/GIq1QLbR2ESBV5IG+znwIp64H3YUrO6B8MEp4G2QfyFwH9s7vu8Z84j0ZKseZ2i
BWylkIjwWGP28Pyx7frVb2Ss/mE17nEk8dZBS2xo97Rj0nSUt+YnIasfhlco0fcKIhh5j9ykA3R6
Dqgy9TFYm8AlgKHePT7eKJDnqoYMB4XhzKlTCdqfw36XnnACLrtlroO2gwGpbS+vDU69pOceO5po
eaUiXREllY1YZLCKs+mYefnYPr8LArC3cTKyt1+v0eahvOJB+KPbkvAsQ+0MDK6lx4fslyZN4c8M
HqOMga5zfpXcJ9AMU4PaXD86QutT5fFIP2+RGsHuVquiMjsyDBVCh9vAnPL6eGNTiHYKBYNsBSaX
CtaYxj6fwRzG59KmnXakB/4TXsHn3dz35M1g050LCBhNsqRjeepDx7OPfN/z6dH+U+rkdg1yK23q
dtr1UKLb5rhMnlasDm/SRUazPC3j6KU+ediYd1DOFpRpZJ5dZrvuT70Iq1gSDO6nwdQFZy9z3aDS
Up2J2kLtYSpO8LRvwUJETdGPOdyM0xNUVE/9Wf9vxUL1gOuC35HCWuJ0vl4BOzZggots7mhqBH/q
AEi1rlb9hbGQo3srVX7lBdNi5JbV69ik9+sTyDlfVqlJ7o57XgUtzAVLaC5EZNDBWuqsCgWDuPCk
MC66SuLL3tm47O5WtsxouZJgK67Gj0pyMmfSBx77mXOBZ1IxfqQnq/mi/tqAUT8alExDnZeU4AZd
Ibbr0rhyMan0dLJPZ50GtZbc5BMeGBsJJ0LOQKncenfmscgAUpW6B5dSbyzPgiPAQ7jREQ0rlj13
n++PNpEAcgdsxeKLgWvEIoe7WC+iv4DZVAFtF1fqqcJ/TxMVZtjKsSDs+7mtnAf+pbFKg0EO1Irj
oOAoyfzcln9VkUnBFC7+TsiRBWQfVR9sdNGgnFawf5KfwqCIgW7QGPkmvaCLjMLwqFvRfLDk3c3D
GD/ipU32ymGu/eGrWBePXwcucTykKbsJLDDhmkbbDXwJh13Pc1vLB+a+SxT/oAKEAe+GHoU93wzd
XfHu5hT8DvAGd4C3JRPRjltPxt1dkAIOORRyjYYk2DljgU+Yu1qKl6cNsQRTQfldwUYm1si+okoB
8FgC4igTi7O0GKbPDiS1bC7Dkfr4JZJtVZqmLiZrG5v91vaK49nLTzpETumZAD+g5qjAxacHqy49
shOlbLT6AWPMoUKf1PqIZ/CMbVpjdMf/lKUXPml3T5FGXY9p4dDDYHoRIIE5BswUSxLb2HTXtMiC
d6yPYLbWsJBtz0cuQrmRk8X7sFh+NvjPmMqOWSvdHW4alxuOy0kdr70u2WvdnnFMdJiY1PgGTP0D
GgFctrIJpysMtoQaP/rXdRkti4ysAGdsvXBy/nyURrKhoB813LeJEWhw8mYXaoh6Q88J0ok0bGnS
rFQPNex2EHfRDIi3G4S71uCmzefIKGBzv4EyMM0xZlX3vnUYnaxUBbxBfLU36Gs32Hq8p60Hcy0p
0kvTFHqaU8kcQeDxwVkEd2szx3Fsv43G7k4RadXV6NgTupjFPI46UQiBYMcyw8l+W5vGD+d6anTG
NlQ5tApmjgivz3B6nnG95+Q+bsUZwawf5u48LCEuCpkbIR1+Djgqjd40kM1D1FXQzH2Ahf4zlavr
STCI6wujTgcztcnRupdl7CCyOcx8EyARqjjVl3aqSl5EflkzTIB41IuKG/x1FVeXCdI3GCdNPgTW
eztemBlfefqBfCQTBZy4H41g+0ZMlP2Qa4mRqvcwvfjWfynjSyp7JvTGH0AGCm/jPPvQHA0gcg9o
xKYBM5m4bP/2EzSevLe3SsO4kE1NsaHiYoX03pnSUmd88Qu1Qx+lzFb9RjD/MxhgjQGm5usQ42D8
6YxhICp+Q3vKz5KI+DGPGUOBSLGPlymcAAh6TuGjNSAwdO6raAvdGPM8+iBi2j/PAMfzKAm6PGPF
So9y866Dp+EDS6EYqQkd1qszjUWpwaOU70vuoJpjA7LjiNTLo15SiJtyOYsgAX8Laf3FTss/MXig
Sghu01E1JgVda1DmT6acQaP/g/UH0HNBMiFEPjTpoZq7vJm/10AI0FDJWzIw9ld7juWWfLmB6HdJ
3TM9I6+pu+BYtLGhwvyo7ezeSSco6AwNJ6VwmdpwRrkyuLLRgS82QNzIkKc6Kygyo1UuSwYa8Jh2
WF15nT5906A8egIX9qx4OBgprnccC/iokv1n738ESivyLxwCrrr47e1Oso1ZMF4RFkXO+kI4yw+R
kBnttC2O8X495rhYBd+R8jCa3W9KjIYNB+ha9aF+0YAEfD4nESQG62J6vTgp68qOzkn2Z3LjwHMS
cyvx/gzcI/76KgBCWLLrhJQovkMnyoimr3RgEGyGfy7Zhagy6u+0VUkcjJm/Pur5Oy+h/EGtvyNN
wp//3b1jXDas+gLYeWBgQoxaFUZmBZs01ApkF2NgzxGW1QOjCAR6PNKTTWjuUKg95JntaVpG8V3t
8835gCs+8Z9MX8zNQfD1xEYqyF04kZ9Y/ua1H3AKxdZS8T+/O0wD+kv1krVwNGlj3zPRy1jq9OaY
OQ2uuMx60v0KRr48YAY7TZwqfus5pBK/yi9PpiWsffSWx6oW5YUcgWJxcL9I1pd9YW1JHKL4u/Ki
v33KoI5zlZu1RgwhU3A6ZakpvZ0CrVaL2rtAxzlbIgOEbScFuREWt14cMLv9m2Pnfc1sQqpC95Kr
aU7NMp8IWoTWzYhC7woTcOGj3q21E2OIAVZ0HQs7poqwipCdYxNc3z4n8qxRdYBmZoKtXHIW7FZm
jNlgLlCY8e6tmbdV8uT+8Bw3Whn3snoS8Q3XqgdBBHQ/yZL9aQTwh++fOgv9OGDoCtFwyDnjhxUX
eUIbeIdtKMv5crOpMrsMrvM7wPC2sedmIpmYuiGNxEszkPd9JDaP6fiqL2wiYWQjBNnWBsY7EUxp
urXUH95MWjMZrg7ay+pDU3Z/AM+yRoU6GT3r/Zrn4blBhgp02ptwdk5Q2A1jmvWy1oR1tF5Fy3YH
bCb82XbbgFP1/XRfzZP+b1NknQ0JXKIIHTeRSGHNT9pXRpVkOVO8UPxd6UscukNYj9suOGfmM9za
Ebf7ePltA7PBjs5zgNxNbFdDlQZlL+SqLVf3gg7ZENWucsMsrQniBxR25ofzUfh/ESHCAB7Zxvo/
TCOKWxq4zpv06dMExzOqQidLjFA0aLrr292aOyVa1TRnlUeBBmT83Hwi+7l/lKpCeVapFH+vgWPF
omJ2tCF/oqmCbTKKHHX7SLYUJ0ainawWcB+dnacutHcgPdc1qzkPdrh0oB6GmPtWxkHKXdykXY56
5oI3y5zu/XWxShvVAo7ftqfmJBwwrmdCS5tSb79GY11w+6NWLk/JNFlymZL18VuJw6/Ihm6xVE0Y
eY1nj9PDD7q+lsx2KmkMTR0YKKB9OjVYJGiUfWjR+KTLMYix/cMu/A0VmxzLJN0ZAEYDbyAi0TFG
Bh+XVsOTJiyuhvokCq7Q3FmEDM69Qne2TUwGe+wpwfSGqZ4Dv5d9Txm8LL/yGJ37E9wjtmkcMMOG
K6kIwqGJyGziTSsQZ+NT8AL83JnmycXqlWr2QwUGyZq0e6c4Di3E43CeqwiZRtTOoKLDcGrZ0FAW
NcjBSyepZSb//5ssECorBuA9j6/E4G6sROcvIQbRiOm8HiFnySNnZseoDp53nb1UrCtwGMzLhGSc
33VPaZUpKJN6eLgpOYZcIJIdWasyAiP/rog7Q+ABZWLAoPNw9Sd+ZL2tD2T3AfIOQh6tbKRvO7VB
m0C6orRO6NZNMbvxYuDXSQfjybuI0EfWvIwjYRbSz/ZHYny5HqfZebKNBStVH5UNn/yCNzSGrro1
a/kaUQadsk/UqPZpZ8dXBaEYS/Kd7GA+YoeyJxZ/98MY1YAcQ8YnRpesw+gDBx7OyfbiCU0GOlh8
UJXLVTGiIN05GpVmTaNZ4Iz0DGl1jcVrI2ccpuQiOcIPwNurC+c18peFYiXBf5rfiekI4djg6/bb
kqGK9Ds4dbHv4ZnT14+rstAnFHA+LUrMdB3fA9nF9zztqxWDXrjOY944Gna+LZKPSlTaOB4Ehbq4
QJwTSIxCA7M3TkbiR8GUI+UWwLJ6ncziYUOR4nOnYn26hGp9TtjIN/ZLYcEmmqEAmf8MUSkzb+AG
ipEj6Di/m9Pb3zkM98JDgVdRekWbM3venRvHjkj8jEMkkETRsuK2wKlRunid9ESQrwQ32NLDCna/
Qpl+ZMbs9ydeQ6L1uC512/MBSmSEoIff66yLNP6ZqMfL/upJ7M7Lmem4n1ocM8IeP3gHy++lJhyT
8yr8LvjKPHd7ZHORZAUHR7elFViLs60DHbQ0N3Tp8UFuaDYfIYXW1dngmsfuhIEuteylggwIlCya
bylqEutVKbhtXSOMV5RtCUrnkPFw7Hw6uC5umxfT23/Ne1kJe20OVVZ8Byhh2stOI0xjWjS7KjYG
65+2jAmFGkvx8cV6ly+JVMEFu6vyX1hmvES8DsCFFj5WQZhx5qChuusR4JFTpBdQpOH5CE4sROkB
C3RrMVtXElYK17zpCtJzYGgWEwo9AP1Qra0zJgvcJnEMI4BsayeJE3anmoN841GRAq+mLcqMMgti
/5b47wKo7Hak4+ksRg9Oi25zl6RE3WBJeJL5v8LdLqI43s7L+cqkwvdMsVVx6GpOw/CKAHlvU+iD
gmU6+tUbQu6Pn3Vzg8MHKA07H+uLEprknzmV742q0ULQ5+5LIuoRbyuRGllbVsgelRQIf5K1xur9
Ffr197id6vExdT0e4w3V2MopmiQGs41NpPSgxTfCtv4fgWe/mZLF+Ab1wEYRQKdKqzvOhMs65NyB
ItOa0qWetMdfbw07DGPhWVSlc2ZE20y5hNn5zVs9mnTY6Xwvwz1LeLzPrd0ng/eyCO7uOIfd/4kY
hgk0dAk4dXLRi2wnQdnABgpD7oVRrC7s0qCZBzSec9SvtwCRiCHitUHVws+4aC5vw+rDO5GNYVlM
azrUc8segJNDwX3LEt2cXOMlbpwDkS4jApmBfxRlimRrtbpW8pHeMSkCFseRe7d0TM/tU73TLTUS
4iaDfvTkH8jhNVY6qW4APCKSMurj0/ypiggtMmC8cOk9IKy1Bd2u4pYNU+FsrHtzBmp5zbpjisXM
ez7Ef3lOU5TiN6mN9ie94B+l9r2B7L/+Vc9Z4ifQML86gBPQSQtvp+n/bxTkNsf2nQdq2UJD11NA
UgpVV4ot/2Mmvj4lAbvj5/S6It1AQ3zh7FoJH5ngAzyssc+j4ITK3EpOGsHT5zB5aj4jUtsgpY+W
dmpL67/KiBCxtiiv6Dq1BqrJLKNVG7DE50dwV4l0a0rrKvJwM7UDzZBfPnditOkr55c0p7EKkuw1
DLMKuzVEJRRu9TKc4TOxYXT5DX8s/9vTlaD/Hca361+7GAAIUDeYRPutR8uv9rNrciGKECWSYQ1g
WcJqdx3jMuGkv9rnklW3oQC2kTV+l/Rak6/JRbwONLY5v9k+someGni9bUA/pK0tcZP2Gi7g89MS
mmHCPvkHLGBx53QTveFp/Xr9AmmrQdSmc/MYrmIlEE4SEZzAzHwKLD11ZWWZQz8PHcFs/JcP/baQ
S/ECsigKXdnoKI73UjF+O4nvZHvTuMndBjW61MzqixreONXRTmBtDscUHzn539dZp0aThkUiDVCP
rEw3M3AWEr+QaG2JkI7/JVuOUuUpf/bPfN1TzFGIH0mEdgb1EJJTzXlNdXCjTk2HaUPeagQJKlQR
DeVA1J0QVUkA7sJfdi+zxz4U36B2DZbHZ4NEK9/zN+FkaglvaMZv08CVX4lOCfsBAJaoePTscTTa
2K60BClzfVhEgSQTsj5ebemmUalWwFtmiPRZUB6L8QEiZbzCd+5XM6TTx40P8pEZVJDe7mRXppxw
M3QmqQXM9eCRGMG6cBXmlC/fZ1XQBZCEVe9xtApudTNRGzANkYzUw5/avYCyl/VF2zloKSacdS9J
bWh5nIueajapJkRPvJB1Nas887qulUsB8mWbEm6LMv56dMT1N11kQsJACtNZgikYYfA5cDBJH+Tf
U91qjVuWWjokf58C4DRehJBjjMpGNcTuVc8KP7ZgS7d2srD1tPL0d2E179ioPd5IWLbVxegToTxD
nSOMbYZaYj7+e0qnyt+iTzxT8fKz5pOO4c6cKS12EG3rhzfaSjMVO00WkkszATgd1kWs1+GH/lr4
ptz4o5yLFNiSJcvBmJDz8trw96BVc40N62gEDbxwRkxj/0GQK92qxjOLSFjGppmMn2g97Pd1ln8q
IV1PWMzJDbN5otWaVzHHNUhNv6J1/A3dAzh5jfUx32gNs65RAWsv8Ra5X+JinsBN2Z3yN5cXcJ53
PbZLXynyqr6Snd6zmd0FpJzqWJcwtT1nxDevupqHiI2luGdXnPKVWN8TPvNlPeDPjweUHOGFrD2a
Vqo73SOtwqSXz4NOWU4BEFet6+yeYIAfZrP3LbZ3I7SBXWRNB5rOxlBi2B6IXMEnZLINMlzJTJI5
9kLovzgrX39vMNhRclt8twH3sns35xXKWz9wyz4WyjhBrDioPR4aIHMP7qA8oOL5Xzlo83vLGYu2
cH1ufSEnZGdK2kQ1WcjH1KDM4FSEP4Aqew8x3NsIg+wPJQaEbShcWrTXvAlUBZv+s57fv3gI/RzL
9sl/jJm6IZEtNlaToB69NY2R9r21ntfPA2+bDnp8OVh24QLPyr5ZwhGi/AVJd4d8GKbpKYf9HVg7
fc+EiRRbzKKDYQZNaheDKaxSmkkEs/0NlYMEZsucadgr6SCpFKIARGRhCwK+titNdcZU4Qseesz5
CTndKxK+kGCZmXkoqSs6WQtCLc7iJ39wgx6MX85mlTDDUwaLuZtf0+qgRogM6mYOxiqhmIUC5fyF
FMtoX6IaiiD4MQ6c+GltQzPFuhH+0UWLZZQtggqV4KUpuPIc+W6QAuhN9iW3161LM6C5rOgXWknm
k5j56jVbO/nakJmsJAuLftbpYJM6uWrM8IuQ2cdkSRrewwOleLmlwyHIbVaGKQAiTOvKchkPUAQn
nf+yglSF68GOXMfF7GSdQ6n3Jd0e640hZ2u6tG2E/ky9wA/gh7zdwnIW8nURRKmy7X8y8EJc5Xxh
jyDgxjeO3cMqz1A0qj3S/glCQUdyCBDd5Xg7KIAKuWj2v1RPqfLAtWfw8kWbMhQMJZBgJb/kOb8W
FkLe4HP/NKau+Je29kPGzGNFFjMfZdsWrRhPQNEnT9MidiyyIxuqL/O4mRJKEEpe8z4dMQqNKHuL
XS7xgM1/7+HwQGP2iu0f0PwuODl77EdmVywtrTvg4qG0i/h8hsJPL2W+UtJE+PYSethTPwAqNZlt
8BUzEBn3TXGFES0p/p84juiuu2olkhbXmqCkosyC26oQxXbxI26IGJ6Q7UhPcz1dMJccnY2oMrOU
ZzXkk87HsWbMATgFAdE9iCZn0/40I4fin0eifTlNBjvWwaFjsTf7bdqcvUTp12TPc8IwJLBzNcbK
gy14VxgWKPaE8aXCtiHns9TadHqg2VH64cH1aeOJ7vT+FnLy6HRfIiYWdg1Neou68I7BjSCTDB8k
qF3xjCJ5XdyzeWbwCh5Kb2LfY3fBiUlnLWiOt7eZTry8JTz0Lv3aU4UfHqAdaJWnnmueqp3cbCfG
whVcnBIetdVwyuPNIWRp0Go41uc4DMnzBrZHh9M1G2qyHlaP0I1IbJNQr+XZUUGe6dvKBHgFLQUO
IovBQlM5TgmkvpNf/fsnmH/1HITA2HxbN2zNbnIMZt0rIiTEskPwnn8KV2VlTB2jUqI9w03mfV1b
o+u7Sfc1BiMTL6Lq7goVGr2OyU98KgWJZtOdSVk60zgUWogTKeVNJ/NRxeiKbDtiVqInryGVSsDp
inH+W1uQt3487KXjjf6Mp6MK5jgL55Ht2yVBFNmwcpfwFVi8CIHU6wEI5yxkcKKMesgY9bePKnCH
X+AaptJIflNeg7P8WgrT9XnYYbfagn9OCzy1oGciFNJDBj6ZgJ39GOJPgoHaFJ2Xs2vxSEydrkLc
qf6eS1wqdGh1itqNIoOiSgPSfNIe/5Y8J2/cghGLwbs0RzvfRGHxKwR0n/nZdXo7EQ1cjp00q+Qi
BFGH1E3yvSNGUYKh1QMcGiZTbJSH52Mp0i5o4N8wR6hlwlLdPDx/4maCTDQZXRhVL2wz4tCu5+6M
d0X0hvNugpeYS6vYeUc6X38273ydri7W2kpgmIrPstq6Jxe1baQ5N7jaMPXtSAbM+5YG2lE2s1eg
L+0+IdOfsDd6w+KK27rDBnjbcqEkhoBsHsnkwG/vkh8DIWK4aRNjJPOW4tDfPlQesDkVH0PYLipr
FxJDpki62HVMpO7y5FSU9o2fllmelqAjOTv9/SiXJLyv1iew2x54SJ1w61vh8M2mX/tZIoeiGc2W
6Hqn5yOk157E7qHQW9Sic20s5xvlhC5Iq/kJ+nf6xHUUgrVohP7bm0F0nNjEtrQkz3svDVAxUTcG
QrTv4cPT4aWoLYwMXpq+zbhncCxh+q7yEI9lOGUAloNH1dKOOYRqOgZuHa95GxPrnAxYQO0PP7AW
YLpk1jTLIRGqrUiY1/iT4w3SJmyudvGqDeLdDtnXs+XKkspv/0mnda1n/yQ+1qHycKP3QR42TT5c
CY4Jd2EvrNoLK3L3ydcrJghTxdwsFcjMRTqENI9WdU6kpjwZBLv3OLjWXKK/mxd2kHpfAeoflKVz
YFLthSbJnbB5+vHRYEiupv2IXaM7gC62u5HZl8BulILza4kqKl7V6xbJd4sF26Gkn6Y+4vsukdST
/S0nnSWYT0Gp7rKEo7cNJElRMZt0p0AewI4bfVf/0ogeBco/3geVsWzgEtspOPtnyjPviMa5+Nhy
q5bL9WlLM9/hdSdqepXfqKzTAFfr/bHP0PqEVt6vIieoxsUCNCtD6piKYyMYSBfxUgowhfWy6lbQ
qs+3HjTGyBpcrGkcY1isdULjKRNNhsrhdTpppX9LsEGerLgXnPD92diP+GZCGHbIwhu3EpTV0u+x
r/ucawBhWMpTD5K1bV82f/Sf4Va4/118Q/XFH1IUAFJWNv6wulaF7keCu72xjz6mE0/mA6zH5pYO
8Y8MBJZFanUm+dfVE5PoiVNBuG1UJm+2Y19NolMlC4O8vFDP+uCibKG08FUTO/xI8MR7FYZyiLiC
iRs0ULxt6XqbiKRl4VkstjD68itW5CkqCaF+nHxFo3tRBIH9SxWtAmz5Z0L0MFmWD0IXnq3UKEcC
7lOwdID1P97Oum2Fjhfqd+sGldBoe9D5e1MtuNWBn4+D4+QnjVjsL3C7aZhLsjPNPIPipeiP38W5
mD5IlLXA3bQqiGm2rFPQ7aJdhYAO62KX3zuj9uZ5g9EB10wnVKIzWdsOhiC78zab598KO2N338KV
8ez5F1+hi7CVLgRwi5d79gbe2fo/Z1KNQJgOTGr1jjU9QX0hGFWtxZtK3MFRFEdP0xFw2h/ZHvG7
5AvKsNMskWUIfb+gpodhW05wPnLeH6R0k0tUlCtkQli5oGHeyqJDDlIGOtASvrqcqx0ueljuqWsr
wEgJY25ZFUU4qLKZjPG3z3VWk/HzZf33+dcM/8qEzxivmcLwp3G55PBYvE+YEDEJO+Qp8uioDvhg
gpCo+qsIZDbn7RU1ZOXl096CMqX4/ajjXqcbvy+toGzzwzCdWROrVPrNx8GPFVIUvcxqJxOg8dzw
9OSAy7f01mng7njgAUS7b3XIcizoI9pLu+MkKiXjHJK0lEc/znRNiWcmyRWLYvRDHJqdOI6bBJF1
ZHeshTlYISL/iLmqg5I3oVM4fAcuv6dkjjP5mGsIzy/9B00EUTHjSYyFj0eN2fsOgM+6548dNDLj
LEH+j3yqMk+2m3/umWTlRr5t5gQNq5JX3zZWPk88UYhbtLcgyHtdszswKEZyw0LvHW1HPL9kjw5f
fWoVngusU2zIg9ety7n+WeqllXuL61WJL33QPtaK5uUwAmnAdLK41myMgb6gukVwqu+ikidfmx4a
9lf9/N90Gm+toEPyD73lkbZP+YdpElUlfYIEUorrlA14o80ezxabZNFA+tk2Z1qDTpVqAf7t42E3
UjU+1f+L/lTKl0zIVtkoK6kZ+y54lxQQkTiViMaj4NmHlkfhDM08N4x/Mv4ywMU9NEJ7239v5pJz
1RpoS873Pam5y7AO3ct1pewyFBs3pvupIwUYbI5W3KjwN4U67VaiPy101/WVH8qFW9ItLIrTfAtL
IUKmYr3vuH3FtIlYRMdlSvxZDppmpLfEZ/OoYC2DfoZF8atjXRnkvRsuBN1PkOWZilE3qN2Z0Xok
vpEu5YBAglsiFvygqkEKHPVSKggDUJo0nLvaLNx+MGIg0VoqP4+Ri1Zo51UcuKhDvkblLG2v6tua
WJZtYKVf2wW5YwMVhV7up/aTbKWrOn+6rLzrNqT7CMliJOYs3BT3AZkaf6LYzEgGbD+2ggA+HjGQ
7ZWnBpIRRrURgKU3oCQtznomRCg9w/qBcbP66QAABqruysuCRib5vqLbugnj20I/m02mz+aYDQbP
QeK6o9tv6aX/RFeWr6MWOM89Z56q1Mqpi3v3L2TqcOcIallNQa85hARwhD0T2o4cZHWJZvvbTc+K
S/EIwxikPRXkcxyCFq0fo45DFTwWBqu27aBJMwf68o5kj4SVaQBvNsC/rxZEcwxyp5/eq/Q/Ho/5
EhXGx2YXQ2KWEf0l80TPnBDwQ9HDGZC9TNTS5cO0G/EjwUj96G3SvDGHBD2lZ4ecoefXaX9fAYxQ
/SBlBoL/8I0DfLd5yS4JJqOUknq9jPzvTcMD1yCoYhcLl4hipKlpfbdk6LAAPAuU4QGC0oyfHqtn
H7WpsYwK+yg1/YfQ2fSv/lXuVfp1S8nqsrz+z59b1Lx+qNsokFleQvyHjeSLwTgBuYi++kWmfx1n
ObgF+VcIYzC7Gr1lCrelI/iqZLqT3a4eo/2G8ZvX1Uk5gIsNelndF4yShpFf4v/g7bJh5mMduOUo
hs42KdIXmRfyv/UWN8KGRXI/Rzngch4UMgHShaypaUMZK6HFyiYLt1x5mVwJhggs9ZSq/5vzHDcN
g3U0gcoqnQJpkJXioC31I+Djqa+yNUJhQATssNWPYQNU7V0tYCPe+ALmJ8aMfwdGEp8gug+wtPJM
gdL9YwtpfEpWOXnOaPm0EbX8S1B3FNBnXHGf6T9QqbcDxVUhSOhPPSsMXHlmZTqcttgjEFiTXbI9
uMBukuTl3h5wW4obsjyAxoiBc8UuJcUpCVuvsZ9DATowO6OHWBrmCfHM5G4rxXKPFh4QvIOpkPtj
7ZUjCM4zA7h3LKP4r0h1S64v0eh4J4ENOH6V7h+fDVzcrkjDRAKbV5Nmtl2fSKz7uqKAHVuqomeZ
s+6rA2ghdn3QF9zFIRNu52hFqJAy1KP4KKn/yFX1KFcc+YevTuaBt2BXwjDVkHGArE9ZCU3ENwxD
L+2LpeqNksfeYex+mYbBrbOmAul/Htczr8Myl8T9QOmY6An+qEY7S7eyO/rdmVVyCcTvJ7U5u2ZX
uUHHZq+ShHdtMsQh/7er1Y6OPRmF7GkMBWbju3K8gdgfDG2SkBYkzLGwPIN3iZD8Q9A2oVmLOoU2
yVfylLeA2+3odb72xXTFSIg3W2ZgqD7f5t20aUEMwFRUKIwkKmwhsK7DUbwu3D8ekmLEUvioUSLv
95KwmKI/WRC4srVeKyXE9MPe8gas/JkyTsgPF+GGT5jR1OihUjfArwFcLoeCVi4TYfXK6erlx33g
64uCh3NSLrtHnitQ0HsuSmgM8AIGsVBnuMF4Cfi0b/8o9Ku3v5d5y+/4v7c2UZSLZ1Y1ArstJAZy
eqG4imuiaQlKSSXN4BGZar4U+Yi6gB19hNsC8keBt+3oA+IpMFrVVGesM6szK+zci6SYdIXeSDAo
kOPI384S5lqiBL4VmSRAhlj7Vgg2Oq3BSlBnO8EXBCCEy4vEodM7HUQq0Q7//GNUFt6LRmEUeY7W
yMZBiT/cGLvboqryNfgY3xmrZTN6/akPp1DFenge18/18ElnjU7+uhB2nIRnU+JkfcIznqeB6cIB
Q0JHWx2yY62EB+VRLoKIeFLvuwep/ik33K6kt6oV2caaU8GaBPQUOD7FokAbJwP/zjDYHgrb6DGq
9PapHpjiAlrcx0wPvmGeYN1wQs12EKD6rB8QMxjx1UgIKFoWnCHgDtSZ6R3Fj8+ncYcMTPwZe2LA
wwU2QhwfJt6lMT0kH7ArJwe6v911hQWL61qZZNZ6582Fxu5n95BE4CKm/+pKGfUk0EVoZcvMOvz+
IT5kNZEk7nfI9JHD6dTWWiL7UIWMRdubnjXor2D4yL43D96MUE1SxIsiBM8Y16l9IME+n1iTEqjW
UXhF89PEJcUTImKp4vEThyM4bIkEGSwMcU/adp92Qioz+3jn6kUI4+76AAf4jv0aSS/wawZDXbY9
i+ofidfccUgRGzmGI1UI74f7rcCq1CnhwzsDPxzN6b+Mc0k/Ros6e1bfmn2y+fVodlLtZ+6T2nXF
XxzEA8T4pf6S5gdxTajGI/by6d4PSixL4wtBXdTBRvsdSk91Q/PmI+6ImmkylasG8pf61/byz8Xd
41HisM7Iy2XToExvHqmcsI056UD3wLBVXMzrk90a0LLS/G7wwx7lo9qti5PNQCZ4GTs/MUyQWSYn
P9d6tU4UBYUe5Ow6EmFM0Tus5/znzTtMmpFGfUhN54c83RArOETeAXfebhsjdYrDSMhyCYWBC9LJ
Bi6mOZeHqIf17kMDmabu636qM9yUtGgZKeVZBrUeGaj1/ufPsZAoFfCzcpJ2tuXbwGSx6kKKWVmK
0BnhooGNbXyWvsbCtK/ZwslatTaafEAmXDlGjSspGAlbi2v4wK1rtdclBECWRik/6s7ZknOKif4R
RCnltAr9+5qXD63PSDbN5OqvkZ65vXTUYDmETJYxcsxxGz+2AQ/IRCSP7V9DbD+HOvZhvd8HchDf
YX9EbE4DajHkzm7PEj3D3aaxVEE9NzNlu7aBuUFLQXq1UZC51cjC+ipEP1qKAGIzFsgdbl0aLqSE
bvYlZFQ+qeXxUj4q9J3WMqJc0XbAwlqmir262wRauTfpCo2Asw8MUvsC3fPbx44lz7HXUkMfZ6X/
9YJQB1JvCGYDD8RQ9p1HET5Iygherj2TwPna4hrF7BWXi6J/O86PLkDIv5txSCqlbwvO9pgHCJcV
q5H77jRTT5y9hZoixiqazK0mH9wsN6LBe+cvtyuyFpOOk0oun27X+Lji9ti4z59baNGVsGaMRkRr
pFZnlwgdHMQrGcm1OgmCr+uwgc/Hl41hBS/HYiQYXiEbQ4Ca3IshN5VtfpbqO5rf7W7mwYTWHsQC
iQG5Q6ovsWdc/c3eoxGAgOtaqEzeGA6Nud0OJmquY0VBlnPLzdNsm27fiwXsrNjE6fXzMwcksKtf
ad6KYempUGaRUugIOhMjkGij+74OIjld7s4f67AIabQqJPuMx+ljwhnUJqtuo2WjnM9IDkFDBKN0
opgNLZaUzq9drNwofZVy+9EAG/99S4r2R+xqHMBw575coZ2VMONmPhC2CLvy1ntXf0JXEo3x28D6
MhSgmTX1LMaxVBPHfoMru9C1WXE6MUhqqBXgjAn/Ue2ettp8pQgb/8N2x7paqSlZ1NeFO7X2MFBr
QH4yfdE4skH5XamKeNqO/ngPZu8w07v8SUcbERcnaloF7pEx/SZD0sGZ1lYq/LxY+FF0u8OW96rP
RaRfjZyZtpD0uIEuxVrlqsb1beVPQWWW6gnEWMfBXte1wwa+7+RlTcmU3Qenjbl7av4MtjhLvBYl
tltFC78l52Geth8oaFAahYRxZlTs0TFn9CN4n5YD0Ak9patG3jRyWSVlqHGE37lysNgvVR31VvRm
DXCX8HHu4j1pfgsV2OoFQFCcoyAVNIqGbC8vafXhleJNkkRIEZJCCfa89xg6QqH5p0vVwwp2kt4b
lb1ym3gF4d6duF6CDm7ljgm/+f2jEbOn9i/E8uksoTE0gYbqr0k0T12upA4Ik5GDgGxJRdLK7a1k
9sz1x0aaWgK1OuhSP2ob6cpq2CJY+1b7zlCEyBmEyKG/HDGkILozU1gfS6icfOequlrb10rvEtox
UxD15/To3HbmxJ6clBJVgeQl4YJftZ/E59IVqnTD9smiUXE3db41ZkYNOlNzUz3Hb5UhTUuAgEX0
HsZ6TEY03RWdR0FsuZ9/bRhU6sNM06/1GPhVv7YFPLYkKbaY3lUE2iLYQoqkdj1cWMhUYwjsTQgO
eyvv+lGKpTU/BiXhQVwzwt7RcOWIt4GmveJKE5CInZI2Vm8xzIVQDuVXDY4LlIQOdlqXT6tn8nR/
2tf5zXOW5ZPtt2GO1TkLf8aRYfCuTsMm1nui0Z5G90c/V1JzRd9ATxUTex1UzS+9lOGEGwWNufZ8
oo0Ey8YobbXjB3/RFkDwbf8UA5EcCbRhA3w5p3IEu0ilD4jrEqQ/kLKc56hXOTn29inKu9YZXboB
Mb/8vhUnDvEBu62roy0bZDtJE03tJ7/5HPOrPX8mN00ta1jdh5qBJzu5NDGK5zuDRrDB3YDoY6HH
0b5LRbAb+03bhXPqbvKTgfkhUC4V6MzuUZG737F6wlaWCJ+tDlytCD+gJkeIN1Cdy9+sMhaLuAgy
6oy9lEhbAHKbsbkUZffQVxHEYunqNj/XSsU9vRyi5BNQoehyhfbx58TuYHsT3fo9Ghw/dEL8HV6k
DPSegLQy+sSSJd3NyNuny+8n1dfoPceP2eUpngxuNBS1sV+nEI/LEazMX1Ek3U+JKmyy0OOl2Ydz
ad3AkXqp1Pweip8nMYFStejUbHLJnWtZ+EVltoDbr+4FzWdhPcuOnZfBc7II1fvrJkS5SRRvoDIU
sGjRMQqpWf+IUkfL8I3Zi4teDIhaEKE9gG1Khp2FKwMnVVcc3C01zN9YSEqHhLiK/vDWOpbGYvg0
D4aO03ZMp3mO6oKZO4jKftMhdANhIESr404GzCrIEr/D/q+AI4buQbTAQvdamsLLHRuGggTNIYTk
7DRrEv/Tks6qfwGv7WC/RnM+GfAHTBWK+LEOiD+JhIz1NCgndgGwTCz5BS8RW6jWYIbGA0n1+JwH
Nik8GcyinjA07PzosUG5snR4jgfGFemDp6N/8nRiWo6AYYfQd2wYl75+YK7aKpnXe/HEUjHJ4zyg
d2CNwBGbba9BMKZqd5jFXc/sM42oMiraRyR9/hRwIa5nT0dsr140+K9t4N6oSumAD47BfUPojNv5
9QYc/CJJWhNm1kuHfLcZCEVHGJMYb2BNvdwxoDFH1wKcW9oDFHy5ogEvgvNEpj/JxfqDKC2g7Y4d
8+1U9LGlf4RxbAtqEs81K56Ct/8Mc6B4NtzJXm32wp01l5T/gYOq6UxrajaUSEiQcGmYWGpxEwIk
bKx9nCrk2fZmPKZVgMZm4+Aprtyp0p60LR4o78i8xK71CxQ+PuaJ4EGrusH+FfVnQO92OQsQgj16
La5P/RvDJqGN+7ibDnbF13J8Tbe/GNa+5EQoQRdLXPn+vdyDx39gZ2nbaPDlF7zWLlRfHZRPWBkz
FhM5wC8lrOMv1XFuEfS6XZEWeoD+7Mpuf9H/KWtgKnv3wWoGfYPee6/KnzmxnHRO/dpqUKRqMYjW
53q8xqv+rQzi2BP5bsC0E0aZd6170v/ry37DRykOAtxScYFlH1jetr0vkWTTrlt988F5Zyk8oe5k
nkheYITNvS9eTxrhDdXNemhfM9NDE5Gl5T1RSGgltdFuP6MUl0NBo7Yjg76Iu7nf5e4sVS8yrwGI
bO4VJT3eMaKEsNoEQ6WwMXw16t7LoQPCDTxRePZmAH98X7yC+iJKlQj1znhPyWdQ60b6ipVt9n2T
pFzZy4Hj9C9Qy3oppixXLUKyDCkikR6hHqt5Ct37ql/VZ/QhhH/hDIYzLpuoPJuUkJrnhYu44OIZ
FuvPCW8WSSLRPPq8vcOYouGconildBhavw+aPm1/U0fhtmqDu1h3/KmjnpC5OBlQxcQP2z1OiD7T
ikRl3bmDpSOv19LOP/Cyi1MMWYTjTvdw4ffFbelu3qwOAfVrOIu7GhpkNFhFzZpgvUz8yLchjySZ
gwqTDZuGGMov2RKNJuB1KSJvbYjs4HcAJvk9aQy2SR+d0GrGGVyuZMBQuLwp2fgOI65z5IRmQSGv
qSFfXc8hjd69W4jhkgGM0JiDIv7jh6s4652kE5yuj+NyvUbiWkgF9KzX2MB5L5/htXu2QTMSTxVe
tYrLrMUKdEEJuUEt1UqqMf6Mgf2GOBaNYy96glpOwcG1VCcNl/YLTtOV7+T27zv0nF2dF+h4+lTo
+eiy244W8QByP45sx1QcJJpn+ZGZsHqfchIYNQOUsd6RoCbgYJ/N6t7nwf8KZiVbfoaQFMUseKZb
v7Avi8W+HYQwuXAv3/gYTzx7dpPD2ayqX90tjw0oHEDUb2nr7ZiS+N5HWC1SaqZjLHZwHhdyMmyG
+cbsxGErS2Gr/1F0WXmn8D2WdMddwtn3LxrDoSig7swqOhYZlfY5JCOtQwfvYZmKZ4FXX3sQc9MP
wO7WWFngsr4yaTFa7clQz5WpL2oKquJhw0unlfD0mISkRgCCzHt4QCUCenmO4914MQSPbyhKfpN+
HS/LJX3jpkDHNOE5g/ZeqJdUla+MFG6f90ltuCxIqYv0sXL39NpppIfz/qg5THC73uaCIcte77if
xrObcVtF+eEpNaAuk7gDWy8Lzp8RsMquIUCwefCF+8Z+c36Z0mjShPec4yHFv3OFji5JkFBHmrPk
XweJNsKkrbPIMxEtctUU0YO24duF1jPp9wm0lnS7p9LAF9icyFDQ0ZDoV9uu+fvVIRtO7YW4ciIu
4C7Gs5FFBvULcDbfNZ5KbSg0/SgbJX9P8VQpBe/ERihA4MIKJ/XXV/P74D+9ehYl/lLW5XKAtfas
HkBdMH8Bn52GyxICx5nsnYQuw1p16T1YeBnR/UEdabHBVSAf2gMhC/vH8Y00+8vSBW1WQY16qx5E
rUympUSZnVGMKKbNCse/S4E8MrFZwVVh6Xt9CwsGXohMcA3ovjENjm8yOG5hSWAeDoEvkU3aMUI7
XMrwqdAAKEoXn+oV2viaAovLR34pSlGmxLaOQTWffx/YHskvNtQNmYwMJHK6EBfwxzZsTjppMTqY
Fb9CMJf+jOfIdXolNgboTzvfD4ns0JY80Z/xUSOpBmt+3DO8gmoFCPuo1F3NFC12QpqvhLO6hqRp
CtxRBHODqXCLHYHxRA2lOGxAgVovGah4diZ9i3iEcQKE2I8jcXliLsZtKnb7MPS/iDv97PhiomWG
VUvjT6E4oOWr1yJcxXNTRmBP8C+ed4PYJwQIMQSDhV+Fv/naubYNj772ohywa1bOvkfkM/yORkzH
LAW2CeCF22vnqMcM6zFIrSlllBXm0LKJIZQ3fSNOGOhoUdEyR6gqyG23h6D/0Q/AKZj8LXV3JdDb
XHycWO1DdITwz7mqNSxF1UB3UGlImvo2uxie777Lg/tvj6jjtLfaZz9w+n4nES7vGrKy2125mU5n
Mf4/jNfi85vKlIN2hQz7YvsR5oXW/QCkeOogKdPGEAWQHK+BDVaLq9h9gXEFcYGNNHBiAX7yjTGu
XSGlOtyZbXuBiieTE4lWAU8HXwXCplxqH0hOxAm2HZhywlT9NH6P6BuFRmlkNP4uqTDMjupaj8eS
+MoXabHr3OzhQAGMWORp2sXg70fwffpA7AQbwnVmjUy/OJKjzZs0jhPqlDQkHnRoYyxSxDPhpa25
CTsF4cRLNAnhqJd8RksTwAPbIenS9MlVjveDB2IPvQNVEEczZD5dm7/UJ7Zi6hQ/N4WM0ZKwsLM2
3Ylcmo7npKTV71AzIPYIWnIASsepWropUP/K5kwNO1ia2Cj94KMLMXgmzziemkV6QIOb8F1HLHOJ
7QdlAJagY83lvQeIUox/rehcXdOZQRBW6jWQbyzfzsLX2c5Zdms5yaE5T/tGI97cdWh4b5KxGNJ/
a80dY7t0dM1y6p0pK7rq8QqKHZ+Mlf04mvJZYkAFwRe5JAvcQwuXUX4TtrolhP21OPZw9T2P+p/k
GXzid4dwijcedCnADNEf84XvfM8k3T8CC20DYceVWl+E2gupDX5pPa4FuHda+dXLfI8sNgi+AWcE
VZu4Qxx7C3kWVQE8jPIH/pS7q9eIfTjOwhDWwWQuBIF/46I8XJfuxIxRuXxVl+IjgkA+aTnLKTCP
Rw6FBmFnnWDUVbObwt0J6RzcyOpw2s8Vtm0ya6pESvYdfQ0TkKkhsm7gViNfdNrSeBgtp8co+jfb
NRmAeh4e0ZxDrYQfc1DO3KhtjisS/+OY6jHuUFQyexkrvRJrcycGPUUQzKZXJgHs+dllsrgAZjrs
3ICGZjN+nRakK3fymptrFdxpuJKamb8bi9ZxdcLnOFxAs/DVWgsypIiV93FomG4yXJe1quxtF0xE
ClrhgjKdVLxLgKlS3aGWu2OP06QEjDuYKiwz4cF6VEQgEZhyUMq++M21N8MTsgtYZfRGZgELRppo
Nw60VMKD44KH9rYjq9w7d5pwfBkXSArupomiQQcd0p7EqZ/9/5U+krmbo+nnfIA3XXcLNXPfbuX3
C44jbqWpwt5G+sBxS6hLW6wOyaT7ihn36jYK28PzijHdzQlB8PDCmyOI0CWL9AatnjxLIhR5UvL7
JGMuMI0vDrwDAJ+JluvePPHPS8HY+dBB0ScKSVbIsLKASsM2wMjFfIFKgk1R8y7PjEiSs46uWT7P
R7i295Gylg+CxlHFvX/WbnC3sA4vSk2IZfAByLx63pQO1uBlLPL/iYIQD/UuSDuhWLgluYN3qHlR
9CpFO1Dj/wmVcsi4BV4u7xq+HyKZuDxh5tbAE3+PugZz03IxyjfdxsZ9oTAMBrkf+4nY0x3FLMId
wzK6WzKsFLLT1u9zIeUz/bQGMmXxvcQdbauLJMAeqUT7OMnlN5FQW8cagrDo2mGxx+oS2TqIsG8T
US2MNKJeoS3+7Ln+Ph0oHFWFS6VQ3tmWmpQCj/qnTIsNyA5BCHc5F901kU6bfayVcA2NC/IeAD8u
tDXGtk+Cqnya6F1EBlLPfvnYaH5W+TfprBOZOI44GQD4v74VfPoI0VKeqoRb+xg7XAAMl9IHoWqi
zvq3G2xO2IU/IXKPGA6SVB0sfux7XUdvHWq3lmBpuDTBslt5My0swuzQSHckq/29s3twDaCyOriM
voMsGyPIVaY70j3DVArisd2Gx/vi6FBhzRCJgAEhNMx+ZqbgKagA0DMzT1wyN8WY+pQytpM1HZH1
1iDquElRCNgKbNNyW95OL4zUhq7+c83oIX4sI1grAgPdN6gKenY1mwJLEa3dP/C+6ePtg4KZIDYG
1XvtSFE0Gem24PRtDn4X5Mo9iEoNzZ1OlQj/KOZXRJ9uopPC66cXtmBy9Hni1rjja9sniRvSRWiO
pGbMQ4R4CsGPD7eywz0j/gVUblsv1o5I25AO6U3H2ihxxf1p2kUjEnW79oTyeseWS/Q7E7yvQi2X
VSJpZh+Gh1+Z+LOAdAdVrHMIQTLjuuM1zjGSRXzgmdvNSrBtuIkgPHcwFaGWuPCIFGk34hZ0g4nJ
ET9H0QqWgtbxABgBXRVbLxme9hE49Lg8MG7idXO+LLbfRZdl3di1m8jAq3r5BNaqJXZrwtJdzW8s
xO5acApnbM++0F94U2upRkbdMH2cpVzVUQxg7S/4SMyM/iwdnHW7gkx5bcN5/UZaAIfvLFnAbSTF
lP8e10aSXLokwgxcvMxePy7SHpsSzlcX4LsYImnqsCQAl51Cwggu0j59Sz5ePAYhGF3QgGqpu5LQ
4wMHYudKufORWZ8R4cpG1BNlqpw8qIPJt7W7BOabKbabEH4n8HhDgnYvqCWJQPT/+vhf4vCvzwl0
fIN/zzzpjoeaXZv7E92ynFvm87nx4Ro3EOZktvT890BHHUUXoqXBTauwz0E0Yd/xuaja/xr8TJuQ
dI3ny/aAgqfsHqTmmD9IbCVDJUvl9/JxpP4tDgS2tR3SVe+t9ktlO4e5gGUg7el0t6Q24S9HRkab
aRrSjNhYL3nOxTH8p1PuHklx3XftLirdgUvTzNB8sjihwOYrqAJZEfCNQv4S+QqTyX8SFNeZNhEn
0YCfqrW5XozTwqRJTsjWchr8V5vR6zRt2cO344Z3R96w81ijpNuaRNNM+mLkYQRTLKC0W+LFWsZX
/PRen+trI7RpD7zVdfdkr5QoWqNe31A6gWkTmIpXjoKC+hBdh+YCqlSf5I3RnXeNhsHwo71v++ad
XoFr4HJ68Zv0YZLHETSVb8ThmlYDLD/5zGtBj9CM8W22DQVP+j7R9AWB8ygNFRSEBwYMKoppqhfx
4tUqs2mJyFLYrCdGrdS5nwqKvwx2yg//wdKnBSglAO45dDTqJLBhOdJQRc6WFuLacq5Ahn/zGjC2
/sG2VRjCVeARDzHcC2k+9F7iEqEYPjhcFaoEjxKvT9YjbHms+kA6XRvW8Fn9+4n6Z/xQ7FQz/ZNa
Q47xOStUvkuqucrrK30bIJBKswSQ4bXg21gHpQWJuJTpq3S/+k5w7e90gY/7xPc8AP0fps2kOKDF
Tas0We2vTPLk/KLg6hrtKXlbM98ZWceN72ZemT17SIJYCCR/+GuE3lWjmTpa4d9oZ0fB+lomSr4J
2F66wr3xQLYVwzO0t4vFL7XPuSh0Q/Em941Eh2jDG6uHpnCVbCB/1Snpo/d8BtAaWJkNAbAN1Pbs
Rqjnl4QUuoG15gGXryROHXVNtjOTW+DrNz4mBc5W4DkBXho05oR2efwdhIzHToRz20Yuttph2/JV
WS6KjfzXQa5WwT5HbSJv1lFehRlkJpK10EvnqxInNyi8iNArCiM+q/amN2P7fLZvVYiavK0u8ZDa
6hv8BA5LSYM40DLn5M3WDOnC/+28b9Aw6ggLKYuPi8zDvKaa/YRRQkBtvafufCJJEdSvu09/LRYU
jEJ09FNpQN/gGmnX3qChtsPREghHB/3cQhrL4iWcleTyc7r0eEEBaA+M77iLxymneObq1i2ULRgg
m+1kSkC1hmMGz5uag+0APxJXl+wCNjYq6F61d1g20QPXQj9ocI/s5cev5dj6IwqvlCFC8y6aPOjm
l7bY8wIxlAKckAbCM4WwWF0vPGcNE5WUnVDEwttX1kfT3ETWDseq6b2g7i7WJvlxlI5YVVOfPF4H
XWVlFh2r0sznanmC49HJ085qa+yq4Xnck2gMoIDj0V+2pKdi2zfcQEl/ibFYRt2KzWQKGVDzAT7k
ikOX8N1nttsWgE+DMfrufE/EoEEgqKqd5+BadSr12F2BFl+M+VZzGpfFeIe64DtTJBrHXgqWpUVX
+ovIirw+7YDQAs/cZ/7cSZXvdBVweJ2dx9J8ihY3XjJxckees1ofRzdk9hIbMrrWjYjCfCkdzbvX
+vgfoZ+vuuH/B1KBP8wMTtCRN/CU8yRJrEyRHd1fj56IUIWlQn1q1lbm3nHgvY6SqVaTB0LPhRl0
wWV5awpx/rG2r2rnEzfHIzVymflp9/XIDNnkU285HgK5VKlrdK9/XWsiX2Z3dVuHuikYfg3sEl3I
MK7W3Sqjqb1edL/yRdtuM8y+Am7Kx1i3QiIIpI023E0q77ke96cKPR3yNo7gwfFnlm5S+w6WGROD
TSE2389S59LuG2VadtbxCMgwQ9F21J8AYkOeuU+gXk/OwtN/jCL/4LVdAcqgztRmx1iv1AR3RBH/
4JxAzr716sFlyepV6T4yEkke2aqKPGTdoPPdMxX9BbjjbZD/5nZ9QktJSvGdElE0wwmsPyHnntYk
AF00oKpwAy2kLb9XU3LRVg9JXTIvtEtgjaFXX5nM90tJbZK+7cZogRkZXuIyv7rcSfLx3fdcClI6
MW4DkY/3nWkZ4dPlbiRia3qVJi1Z572NUhAkbHvtcCwrWVnTdkHUsdxTAKfqa/EkJhDhnCDo9+nZ
NK6CpAScCcO1HM+zqXPpQoIdTsMgN+BG8BJAD67zOkNOaC/P2o/EfVCItmMEBkOMtr7pONJFDT2p
ux3SYG09Z7QRRvL/N0aS6d+N+J3H8WIirzeCLQ4zzsyFfxn2hqC77R5VWArVG2HqCYm8s3dWvADc
V1H/QNcNaerpq/Vxy7uiDGFwtk5YTAVtxm/dH0WKt4PMraMJ/xUA8D3JE4MjtWNaopPdpBm+G0MQ
FzK2d6CbjVAaPnjEmx7KzGn5RdR1BtVQQ3VIjhtb3i1C/hEvwFCLcrWZMyzDdMK2ahQgoklAgfdw
qT0edpeNAq3nGJQRKBJIHlfFoT4LHeeDWWvttbrXZBQjn3HYGFouozAzuz0MFpxC30nihu30iZ1r
zeVslARutw/jO/ZdznOa7EmiPSkFXaKyngPIxiv7cxzW4x2yj00StriKhQ9Uy16EVqdpdwvLLIDC
CkVNR1fc9wpkpiagUjHzVXPci8e7CfWXYARrM3uKSOcxvZDLWIKroPHkAaKPRJqdxor5YJ8Xoy73
EannWi8SAvkyjKVIxHSzHid20EACkaCBS47/XB3jt63t6cIa0qKdNULgEetYkW/0FN4OMEUgtG4n
0lCwniLS4Y83AzV6xnHfoMYHI74mi0X0bgxDOdfDh6H0PIcjunDxVDBfS6YJJfOnrAvrBWxJooSM
mZfiTAISRaE0L11CVJWcUG2hJruy7tPxhi1l0X1v6+O2HdAxK3KPSos5ld3dq20+Lwnz4htKu6ji
aZh9sFVgQ251M+BLTg3QzGqx/IRvS6J4Jz2G73Khop4FJMG/MkvdHG+WYFuV6R7KcfKaPbh72UTY
fACEjQEMn28vW7gR321eKxyTfMzzyYqONbYJiGzgBmQ2xkLmTFJe0sS+MnOWJSDV76Toy2HcZWeC
WHvM7TH3WafkI56NtcKlGKd5pzUm57Qk/qlvVuZpEJKJjMBsPOZMLWnOqqaSWxjIT6pRotJssR/j
vL+jKdVAEM91beF2+7/bq8SF1rlxBOeWQjZ0u2rwnHJoe9hPHntwVv5Vb2cZBTkLe5FUbCaNbfVC
Okpl0USBdQ7P34d2icc6RAfUZu1+6ANpIDhRiOtGF+tIeDEaDeVs2OBEb5yuxxGBb6Gco2yLxx+h
5GwPd8TagPe5emorZM9hR37mwSQ+fhiwTpmZ+FJvBWRQHlYizD4vFe34on9WU4vrTDCenT3qYfzp
eXTzldeT8CPFLX/Dyhr/FJj52p736CyXxpDEJcCHYNetmcFpAtegFDu/hrc6/bmGViG+t2riRQub
GPvRUHAcUQqftPdpi4oZ1o6uXLO4piPK4on0XUK3rwmkjzzfyPb5uPRL+8fAc/fegQfGvW5lndvp
47G2UiSLhhM4Fkz7h+cJg/EbCNZIbFhwQbGcqstzAJ6CjDSYjYpzWUj3M/7LuNGXirZtyD3oPIR+
M4dOplLh3VuiSyF2+fpxI3bxgXct4a7wZgKZYePCAMnLV0KbTmvwh9Ro54nfVlS49Ac+JxMYEJJV
IQ4ZCtvpg5sDO4n1zD7vdCA1k58DWUH06+m/+drKH/7kS0g+2v3ZEMcCGXej5z5optmeiUahQTqS
zgGcJWbKd/QJOeck283UIhA7mILiXfPcfQIdsex1tKL0tmtoMkLqKZrGlp1jfiFJaryc3mKzxiAK
MdykSZH4rz0mw5RM2SS/4Z2Z3yRyO4+YU/JD7D2wbWoUFnRoL1hZQKCC6Fhhqz/tFNdk8L7szXkf
MWARRaU8HXKf+A7NrMyI0oYPaWQ1NPOQxXx7UuG4iyOEN19zw7n2o7p3mr3o7/vuJw1Vx3XC4o81
iNYLH0mP45XmIQoNee7O3ljuDG15/dySJi8NRUc8k3ighS7rZCDZe1dq4bZCyI1qNMZg9JITthrW
NUoueQON8QkTN8iVyRpqVw1A4TjW6vIX0jcIo5WCcbmXTnfydmmMuztkhIGFg0EOlBwT8Aj4Euxz
Bl12qm+sSeVlgHiFIGtEtM2OyHKjOrIwZA8zHSTUTLcQxT8dMw+LzoYOJAmTXaJ7pHb2sY83bi6Q
Gs7shY0NP+zPL14JoNDwVhykcq5wXeSGdszbJmM0oXkU/QF9eZuOHoUalcRvjRsI9kNFVYauemR3
7hrkHv5qTlak9s32nYxgiueTIuje1KVRTXTIol3Jt8LBEE7CYzDG3aSVeQ3nLzWwXQC2HDUXQaEZ
WeOGd0r6Km3PNhurOt9oQmPEmWxnHvMbyV4A+bIrwYSFeZ+G+9r8QmNyaTLvcvhINE631qLQlNhW
gVUjXJr/sgm2D0YJajiFSpp+NmL3OSAJQTND25D6XH1Y1rkIPODmsO93aKWHB/QSYI2Ayp0bWIwQ
mntk+7DGs2tABUVnjmruEQ/bKv3BNnHntG2fMWskLmI7XsfjvPhSPFmBKQ+02TWlMhXIM/czQKCf
ndg6hm3eanm91m8M/EETbrbi0utotS+k8hIfViLrwIoy1X4CU5CpoCB87V/BiJFgMamK8aeNvrh1
i1ytFnnjPaaA/ocemTkPoe4UdJgA/mK6Y2kKxM0CYf0J4gvKn5Zi4YWEXTkWeTcbtY0RxJ14MA3W
BiFrYelBH5Wl1DBjPmNGGF5FMcBRJqu/3R7DVPz2rM96M1xh7sv3W5DZhLRo89BRDH7XkXPFSCRa
4sJooQpxfmykO/pIHGecgvnw13avcGuvS0Sbn/Eas0kuy+rSe7spIN3O1UkKPtPeXjKYjmhyqFng
VOHEliBmt3e6H/9N8ujWb7xOQvqAsSLONMBmmidjwVi0BsTTrY/E5v9t6Xq9+zBZrImLXcSIZKMH
kcoqsbFtXscNV+jEeKVC+UTuReJvKntRxomvH0jVCFpW7o36oO4B6V1XzO04BZv2/mTAeo5f93Dg
OhYZkvOzSEOk7kkoP50tgBQcs9qmQ3nSm5Pxi9q9VkxTcc/la9PItLBW3RpOlfcBN9HdGgOi7wSG
/gT2O099ZC99yqnTUmawBrWLQCMZQvpuyPwwFbAGKGiimR+Vq9O7aZOL3E/H0OeiwUEzlAMrN7jj
7X9iDAbWlyMSWEAWZ2iZdNIEYkjOSaRNqYhEhAO3CpCDuvv/hMyxwTSthLjZY8pjbkqmsvLsIJJM
m5bT8yx8nEpvK8GAnr8P4KohZOkEmH5Q4uaoeppopEYK8ylDQ0ioZHXw4DONtmEu9Ki7yv+Os5R4
sigBRSbwv26+/MH3nz4sgMSiuYX4ZfR6TaDBeHM744x2fx66iIiYSX4MZCzLsHGX2rhV4Ke0LHxo
31ENssrTbqaMPP+3UKaGOQ4yV767osBeClE7HnuOjqD5iTkGp4DRYbWNCQDdgxcKTmZ0HI3Vdnoy
ss7ev+c/LIybbtG/SfAIJ9fmXe6GjKqNbTaCqHWMHMQ7H3cfLlL4Z5szhiekEw+9Ox81VgECAPzw
FA2EPul00/Z9pAWr6z7Rw8gTUtWmdsexeNwfOtRw9EuEbSw6P2WK35wDZfxGXKjTHGXB4Jr32J79
GlutHxJMrnm2yhIYJDdJMZEj11s5c3tl70X3+yPE58jvuI+Dsk/ySwvrEd7JFZDZgu10jqUmA5uS
6RRWZFA1okZQHm+PVFm661jyq6r42pa5RE11dDFXN4ck0BKuJ+qImeuj/gbo+JDiDItkeAn3Erhy
T7wc+XasyINlk6ALgt1wsFruR0ZjZbYe7jO7Z2WMMyiJL7M0SEgrDMWq8dNtji9nvXzJ31E5WD2C
whjOi4RY7hT9Q4zZHR2aTtfn4ITA3S2T5/Y+Ws4d2iHm2JJoll1gii03VsaCOTlGOLsbM9vrqsQB
Tlc7ltYlIDl1YfoSwv72hf90UaEnyzumQFcl9Yuiz++yZmvcr+UFzutKqSFmD/YnRf1Ib5daROwA
CLZ+ZAM4f/mYaFCKVwRXnwZndvxg+jD8ZiyGlBqdkTmEJ0eeHBfNI1kKLWXfvOmF0Wpu/+iZg3Qu
38rQxKA1+8I8bm9Hymn2ObF04k2IG9eyzQ8kfyLE7ZDx+I3EwiwJSumf6eSn8e42P07Ns9yOI4IM
zAXwqdN0PeMMeQDOdIn9DhWkeJvEH5t563KKnaRdFkEJItQ6+7YTmPanDaKGpldu5lpqaPxhtAwU
0yG78mdDToLkZRzc1JaFLlO9a1Et0aRXS+/FSa8N2kkS2jgb9Te9c/XfqHY3o1J3+dZVDjO0vMuf
2AsaBaLm2KrzjstHEg/i5UxgwoEZaFQie7YH17QAPH7xZ2K9Pdkl9HhxLX/cOkcjED4ye9T0rhFQ
86WfNhWvt5frNUzjLRBPZIjgwG5IW39q9yZb5TNOkXeL69uiiWznS4RzUBNWY7KSorqC5aRWV7mQ
qEqL93F6CFitszu7SYsD4cPtuaGiOF6BkBCJ3rWhovVl/Se54LvGxxRoRNMIXVrYxg+SrH2LbGBw
OBx5ErY4RLaXI55RXo33BUAbVa6sxiQv9IrmsOvS0dk+8rBtcKmUtceOPOa5ZT8pc3YGlWaeofsX
+RM1Tv8FX7vwvqbqJTQLQPLZ1xQugAbPwa0FlcnupoziQJ4LhcRdC5Yzf2nDDFYFeEE2NTBzqmyp
ROLeDWCjNp3lhWEGc9/CdsMgNgdeTYWatZvIRWENi8qhOCUUflF68M4clWM1Sfd8d7n8jvi37Soz
TuF6LV0ZJ8EShywi9XfwEdwcLTshNheM/laPVXk0gFWe2GU47s/JhmbAgprnGwL3n0ivevIK+esP
yrD6+da37WVqdqXMJnkFWxbvR1Kq9x2+RRTXCboy0ZetSGTuPmP97aaFYfR+U8DqK4G7GBjOLjVj
XmsxYp5lLdFp7vNiIW/Nj5PnnZ9B4gG9SQp4VI9mokOy8jXMuZrnlbUTu4/B6OBM2kQGdQXQy0uz
8w62g3f1cdPabV8jrdQW00w1Am/B4Qci1DMWfvpWBk/GqIjWSwY/NZ1uofeUacDjLME9EKOfrCmQ
kiBGQvOkKv/FTNkloj6mau1ZbDeGwctAUZixDHQcAF/4YjTr6XoapoGReCe2nmks1AW5HFZw9n6W
tYyHD27XTgWDiafiG2K8cRf3UBmLDULqllBHtzTrfI0ULvDsPvgZLSPRwO2jtJ4kkUtWwh/XBAEd
M8a3S+NPK4UDqrsgq83Q5rB9K7et5omHSheROeJtQZtlC0TMXy85wRLAMTQ7Cu/jqOt+nzk6c56r
s+7Uau7rWcAgnj4/nQVDWTeqYh/+4n49ir7yX4liXvzDXKRp6yTQyTnzZSZCjNCF6q4icB86sNqQ
nWA4oDRkn8HkFC4zJVk1QLxJC+P6jfuWbZsalzOB1ag56ZwydtpyLqXXlM4H7lDyqiQU7CNocxph
xgJLvUOZPnlcjeBRUohNuKJJHsLHu5V4qW54OsuDsHp03r+K6Hh3Sfb6nramiNqgT/WJzpBsmm0O
0u7TPhdsGhGEKpHYtxm1+Om/PsfmIZfhagxNTh8qKLCj+q9ZA49v/oDtky9dQy/1tS3mPbNFHFe2
QmPYBD4Q3DLWQSusqZBiVjNn6kIbH9jdlOVnmg3z9AAg4VpN1pd/Tai7iP7SSi11SPsJ5fzh5mkl
h3VdgtMDyYO1OARlwdGopfDhGHb0p/3Ea7eu/xAcFVId6MmUyUaPobXqeWJVpMpj9S4u+ep+XgFS
y8BJo1TZS985aX2+7bUtrV4Tiwf5hL1D3cKtUV9ncgK5o+7kom/QNOehWd3305tb/JBNwZ44hYll
lQPvZWcwUGXLBftkF0SW3fYz8fGBhRYOy5y1nF15JAiGQF6ObxkfF3Uwlon55+76EWrWBETPiHWi
qF3Gjry3xqDQu/uQPSdr3SQWi5kkxROmIibMwyXDA7Zm099itZmpHo+5RH2hDoD/tWwv+k+QtkXA
qs2angNLta/MakoCTjvOJp7JLUlasNa+aI6bM8wem7eyYH79bi7vVfyFNYiwAfN76RjKRU5Wu7wF
sK+vJP4zyJTAH0dj/Rtmb2cUkmdHQwtb3T8i5L5eoGK9yGaEYcQwsM9v3WNsVA3kF9ANfER0kmbi
UTashbLk1oezuj/87yh23+7Dz2kpuEgJ1CKuqVHr+fkNQvR8RgKgGFm5o8izMOBr5LAIPPL6D6cV
ExkRnEjtks06qkfzKJJ+iSVwlg3UYwz7HxBRW40dEUQfqVlrBOd4885PCzzNvnDGP58lCYYxyLXg
B4u330PjWyczs8kWeLb7qCs9dk4gi6wCcPFWWqCHqEkyYvtLTFPsmb7TIqu6eGqe8Suk/bCS4Hk+
8ztcTE3b5ud7eETpU/3D6UvcIXLdXoz93OC7Ea2YLHccYFMNIqdOk88kr6T8t1GAr2SILABvH//Q
rjrYkHUblwW3AnRZfLTqlaz8xA3wqR7Fw9uwD6lWzuKxqyeW51ytp96J90vsxDqDZ6/bRpyQ5zb0
pF/Onogg5tE4WsvGSCuSnNMuNfBM0orZ8bbjxAsbyOjBh1yofh8CJ4q8/ppMBZdiJHVoIWyyd8x5
zQtgiW1EMebXVU4OtXEiufv7p4v2zeyAHX1sgIGFEHQxONnpA2L5E7Q8Mmk+yrA82a+QjVlwJKo4
iXn+yTEJyvBxxz74Uli9nMKT2pvrjkqpg6OIfVm7OMW1W2cyC+iaPkZMMJoqFDMgybeYcSd2o6ay
P+qj21wcHul7ZtGa26+XDYYM2VvqOiKfu8SA7B0lbGMfIu979/YfVdgIqD5sHg6bAfoMhvogm2pP
fXxuLKrT0MpVYJxEZhbgac61lfr1DFxzBCb9gTPfLt/sNUawiWju+yMPy0CGvRC38l+t+clSbhnY
owrCYglpPQGYExmDqcM/Mprd//ThzB6qom/zG0170DKMfrNFQEwc4Sy9L5f/I1S8/d2THqGXsLal
BwK8FnpHsmVQup5EYn/OVYjpxY7RBcSBh4Ctp1bmezT4PI4+S2YmuZpt6JZIFF1/9bHJ9A8ssOZm
ZF8nsKek53Y01xW9ij8NLIYmWoRAz7IvPvWTVehXyHIFI1WM0pWkAjiGvicNqSXmad/n+01XTrF+
WCvuMC6KSGvYd12naC6yTu0LObg9GNJAKAH5i4zD6OMlgKzOTueyF3KZOUWuUSdEI+ff8w47o+JO
sGRjMzB3TriJF8v+k931lAweWk46Fso8HKaaVQpwEcoebu3hmyhpEd6yvp6fTQr9WGAiDcmiTxTQ
vVQAFHxoNvgKg2Itj6mzkVN66lhRYEO79laXxkhYrDZlKHXIUs7lDnRPtFep9YQi0JE9GCq+6o2V
23AimcUkG4LC8qEI/EBAoCpZ8hBqLQHDrIZUwNeakf4k+4B5iMvOQyoUEzX3buVq998RqvoNQesf
aJLugO/2xZbM35bcfWp9DqNCdfd0FkW5jDx5GdtgzypNu7Ud2qjmHEW1pA32f94Buz+H715lieg4
du38E9k/RAzPuzogbpFL3sS8SvOmKAtWkXuK9NxVWMoTrc+AzIYw6HmiuueivI/umuwNqvfX0uS0
FB4S2gliyG1MaYRIawyffnnPv0qMY2gZoE/kEFaiu6fb0Vngi+2LW3T1Pk+AAlmiVI3zCc4+MIYJ
oj4ut9gFkUBy6/xAaktX6IbqFd25uAmrcljfwF/rVYayi0DT49nj01r8vV6iQQinC/Rze8Iynw9D
vNHaJoAsnpvvSdhPPBmwKms7tp1OnbbjzD9JY0p4P2k6QwgJdupdI1EQiGmWeZO4d9Da1QdFxBUA
EiSTe2ZMLT6nvKzI/rSq18UC3t+onxxdwHeg1Lb3kX2+1gSSPhLvuqPd/8PTPf5x6FcjQJiCPDOz
wkTjx8pqqrUhRWE0GgD9qozgPA66CxSsOwt89le9om+qnSHmWO5S8ByfnKBuQnSs5PA2NCgPoPqa
xb8ilAbG8UFeiGYwmWADSTOOoBs1kPQNMUXY09ZeAi3Qz+cBWJceePkcmLJ4DzIZyrzeUUSoVNTh
BmxVBtG32eCc24FGfLevYSsA3VYsFkN8qNR3d5ehUFgL8ulfYAKehnD0/L8qW38ccMKC4LT1ROBJ
0H0DKitgy7hfsOH7GkFO/JAITotRUQnK3wzao93LCaAGohNY7Nj+q70kj9waA3Bo355V/ZHy9B7H
8hxr+jhMgThF0JG9cnuURoJh0sqG9jBst2TVCPAtseUVJiOKTsB2vZ8HGE2PFr1b9xdWANiSsgaA
uD36E/5GNJ3DFB6ux5VA6WJoTyGDlg38/tYPkY6OFaj6iwpsoTJlsaGTFPuucMjrNPifOSIITxeK
a3eRwiFV2YTeNHN+NNd7fZRZd/aDe7MHij7+DuaPWjSDiHL8kkBf44q/KGIqtbDcYUJXOVXZymPS
QyWTc9pAleJVRnVPe8OYM/6Itm2pfPdvCEGJJZskSAo2gG2E4vAynw2Qe93f6FfabdDuGLK2Ulzo
SMYHqKV1XeHGMTnxW//1OGhtXBcBSmL3OyXFmJ1VBnEjcs4/0SHjcpT8hya6johfP8l2+Rcolc4A
QPuHIZq2Vat4Tc4oM+CQzbKDJrIYPyZ3DH25uNQJOU5KNpQPu58t3poW4rQxJCtYePB/jGdAIjjW
H1ho6NBLlrnjeiE0WM7Rp3ZhwlesTL045/j0OovGA5WAu5X2uBqYdzuT+Fc4qgfUTJ+nK5ZvkEyg
3Skmp5XyFDeCJRPBVTfTxw4nnDmkObawrSda1nhShnU2SWJb4D8CEOCZaRP9/u/vC3ZeuJbrq13G
CHjWUD43eQhtFzy6zWYuJFsw4TacH+ig0zE/1JA7GW8wENge9+Rxgu/SSHxNvEG/B0pMaTWNV69X
3RMF5eO1cUNkbE+QKvtnr5QKIEiOtSSU28esjMWKPVoZjwOmu6FOnJQILXcUZ9SwHoGUwT96x6b6
BwDu2cupI96HO5RBHZrkRQLJfPk79dEd6wBquZ4FSqZxDKssnoN9OiPi6qStroI1Y8SQT6/LQWZO
bd8y5U6YW1PAVmNHKGnB5D06umrxMYpyC+PR6TNDU790uwLZJIZs5kpvC6++OvdOtKiGMpnaeLLG
vgYd1bUHci3r+W68Ii2rFUqg2pMqHyjfXK5wziM6GEa7sRpheohdsP3qreD2ox2Vvh2QtT99Gy1J
cJpf6rYcgiQ9+JN+/9oW6q4jWNksD/L71qMMTcsfnkdREtXus9QgMSxJoe7aKal5jxAE5RJ/9MHe
jABUwrR6Ym8qlGRgHskkJKPtKwyorvG7Vkt8/ZNsZit8aPK8EwxNzw491OokUnXIWbAl6WqoNQVl
8IP46TJ+ATgS6gpWlxOizqWv2ADFSF8buC2YIIzyI+Arhar9oDCaC9PPP5JpWdxXcILfp1zpbS1K
94RS0DA3lF6HtOAf+sB//qHHLacn1IoBlVVCs02layuj4CY4VizsWNeeFyWTSJoe0F8XTIkl3dCM
dwnZujLeRB9POBK82VTk1ifMtfFptS58G29iCf5nhGB6/SEraP6q1r5cGyd7Ze6Xa89b9PpPSSjf
AT57Ak839I6XT1x3AODii5+2D1+kLdslRXWpJ1ud5+omwDoObMAYnwqwS0lGW6JfY44ARTIlqFIB
1BFkUJbAdsLwgPxT+CKwFHGUwEAST09iATJzOJde7SBoojCS1x3ktFpmwGT3kpqLgTyiFXOEeFoY
QAZce7yFOAaZue5puc3Cemujn68dV6HPoqaNMay+F2wRqBFFYcZiMvnxRJvydSmFiaV3KlX2FGny
+iNeutxFIZQ6xdteml8TUAhiETawiB2bRZumXusNJdwCOKp4Lokq8igjusineRsID0FZxgnjbwYH
cOYWoukBw4H65EH/NpilvWdKQvrQ6rEKOotLwhNA7hBQmUMw7bzMeJWo4MTRrqtKmGntwTNRIwuM
uVGhVNIfGfqcuc+WvPVujnOnRnp5lWF2MAVxX18N6cb0hoEw2fBj5XesBsP8edBT/Z6hXUxmCEKr
FHuWJtkL+4QueN0yAMpub94YbPoqqyB0BloPFZy/oeBMxev0UL+oKP8e78kUn1n80X28okK5bcAI
WbPdJ7m7rJCTV+sJmmXDyinFdB+ftwPu5Jak0zaBUwiO+zJYvQ5Om4YPmZC29c1uBaTyOkm9Iz1I
3P31BEjY5JBSsNDWxFlA3c3bX1RUR0Cd4sqJQ70IyACC50OC79WVuIflCtgUxgLiSWZvLTtgHZUs
us0vORqTMwqDKzgXNQ+d6ztSx5/xU7DlknYbLwrix/htu2c51ZPZZ4nIMHZURjzsEFFo8mN+4GPn
vG0H4iJ2Pz9IUr9c7Y5QrdB4RCS6NB6mmqzALL8YqYPeRn0eyyK60j43cSgBSsOoN6vlOH2jpIOt
GqtvUfN0ae4Nm3Kq6eVXn6jUj506hCqKGfoL64ZD9Un68ztOgzwm4hfDMDmSd+6BXm/eVCZTZcHo
Jzxl1d3pUXEfHQpVRokDf0dWYTWSgvt8lpPBz87XjgBCkT6zkChhY+/gb8QuDlHHX5C4tmXqAKkD
4CcXgTepGq8+8/mjNWUinM91/MOXjtpyjgf/7GkcjxK57Gqic2zGP2Lq4hJ35LDwQ3UIhdWEyuT+
jRBs4v7BNogS4kUk56C2wr7L9nrlWGARb7Gan/VAJAAC14NCqYrE6BkR1m57g2kjCVyoRu+ZHdy3
xEFYZIhB9dQTTmzaW1W9SxjGt7Ez3uRnK52694izDS68M3al0LOT81HTHdT0bmkeWJIsDja4qEYZ
QkvFnob5Lq1jftu39Lvr3nel9mWkVMABX/+v1p0056YApEsSaTKGSJEsJ6ondsoDdttG/teCChsQ
X4j7xTiBKI3tCaRAwlgRcIijwJ7JUoRTLawFYn3yakJa4Qi0pnZBzNXme4Tz4j5aSjgbSwrT/TW4
rSPZ1KjnbbdLlw32vp5eXQH9pUEVyOW8m7145jAGCQ83S+kwJ9/T/gIhmyxro9Woqfl3a/C7Lr5p
er/TioHQJgGaiiL9VzygfWA9dukuOjvBLClLYrUwhEGgEnMI6R4TRUH6VxLuWAKvfxqd2rXlIyTt
QTWYMCRrrr9VwXbvqYywQ0G6B3pPSivxR83D3qiqqSyL8MsW8+If8rCc+pzKi9Bd0jOz62G8FqIf
eD8H6IIM9sFYJVSpvR/18XnrazNB1knNzUkvDSxzEyHSWgFI0ENbfFaNnDbOVlKUWu1bqENN8Hsz
1g92LqPhUsqmbN/RbkuxYRxfGeH97s6PYQFrUXSGhGwaeYT93Njo80dmY2+luXtWKylZgSHotjoG
VDohew+aWOcwy5Xi1J0MGN+rffSOIYPz1ODKv+awmGQj0fGE1OZuEhC0aZMpgjeTsCzIpTKPznxK
g6DHmqsFbVqa5DPxTXyKR5QyZXnWg9UiuqPaEwww/kyi544LnAiYilWOBX6pTdhutqZKcxKXUcCW
XfWWC7iMhB+G64ceHCF0X2M84HxGKY6bcwWueXlhWp/JjsOmvkSAiMz0j7VdkX5G+O90T0W9/f+H
cR33PJTslGHWvGIa4HTyNKdtyUcFXE0Nepuzm7c4DzFcGA8gRJ8EWA1Av1UXXRYrtMPxWLp0hnM+
PP/kwWKwj/pNyZCXXEUycFmauOWj2Hcfa4PZCQXGazIOeFdvJWPllL23x0s4EyrPKts02sTrVtpy
oDkacDHc208Gp319+9yj5fHNt58eGtosd6qUvxCJKYMWv9RGWiYqzINdu6nWm9INoOnVweHrbcEx
/RFdmiQS03iqRCZ0Im7iSKqa96VmyICO/us1dy8prY8tQHsSvWSQ5ruWDJg8G9Ag+yzrMvcP1CH0
HnmJsDsp3Px2UHo4sVgwUAWP3BqsgdbDmJQz/myZWKlrjvYjiZ+pr0gv6BnnXpubfwVpbCdlTcK1
nME6LPlCAgqiOV9diaegRvGZ4OyD1YNCwjmKvPmfo3bt7BGtAVV++RtKbTjrwSyKxJIJQ92GsxJ1
dXwRua9iiqckaY5Dk5M7gzZiA6JGOBgKEwFnD6sIw1A/9ryJ69BMuIaxR8WG3vE95Pp5FwGpN/oP
+ipYbAKzDVGOXsw65mWnrqX90u2pXSnpp85PAFxAYB23xrSrl5eHkmv2WI/ilRCzGeA1rPRyR9aR
4gWbJan2fmuCYzTuH4ME7php3R+h80LQRomj4YvGKNaJFNEF6W7zTufslWrUcGxeYTldrBrv71Q9
f0St6LVVoN12oY1BKPz6tceujH4RwdacJwMIhLDCrixKPNPKzPM3L2/zxiJ0DLERm0f36iaIi98L
Pgy8OPkAXLJm79NMWzTEUVeQADQUfk7jTwtTBmBdE3ROOw4VB/vS1nRc6lXT1dqDq8c39HZdrjA6
gBkkQjRzR+0gn4rgjvejelRf0HV5itGMN26rYxWz0Y8LKDWFYWVXVIR0s6qW9NvYwaEeIsAuudK1
o3Eo60lkFkbyhja492b/yLby2wLaxXFR8b5BO2fgS1uATy08DyT+ejIy/NXvpi78V+6BR2ChZO70
GqULWzNs46dUoGMHQtyllwvu0XRSM8Vig6HeU4udRWhoYkWJ+wE2R7Afnn2ZC7oXSnSisYHtfCCa
KhC2WKLeBafUWJ2wujeQYmR046UZaLCJRS+Z+3Qmm4iAbJiOTFvzRJNYMeRokRZSB/wf2Z3568nb
U4+BeO0SmaBUACmvKwq52HHteRWd1ZhPnCJK6xgvyue53GLHjDayJbih7zHvfwH6H7oEDQ8lGPkJ
kP4Pc0EkfiEUazQ6zwYZhfAtTDaYzeFzv4iTSjq4jdYXXvcUa3mVuaeGGUFMoefPtY8Gn17XfoJ6
P0GVNMOS4+d7CvI38UiojvXMCRYYIyfUVYvyOMKUMMgJuIAnLEIIF49ud+Xwsl/vPYCVL3dEOWvD
ACTP7XhGM/ERbRzYKCigBEHETSML2n7pbMKhDfZnJAZKGCAm9HOpkiUT0IiJNiUi+jNrtdttUwk0
nZoIFjWUmT2b1K8GGScuyTmk6bxcrugOwg3fHHs3qBEkOzdigpv3l2wp/1NWPtUY+h9jAh3yThzB
I/DHqEZ2KebBy8FRIJklEiLfKBHr23T0MV87TZqwLQZTrtWk6OiaK9OEasCv3RnSdkUbx51eA/Il
UwO382oxAfPqa4k/bZhVySQG64bu+jwyekxMRJD1vDEq6ZB1agGdPTlNedzNSkcydEgxXXLnWg53
bbHK81gLAkVflT2uyZkn/Drw80jilcBGMo3qhMxxlcAOQS3T1a5YBWqgBxaMeEyYcjmDSjxyXlSo
karMiKLn85vKr9S5Bbqaf0Yf0HZNS+hXTbCSd30yveCwaK8kZ5AXYVuzbTOMuqZfdKTk46wWsSfN
zkIAg2SIbw8GqewIKKqFNinZwP+HBINLwosn+YFK7y+ve3Ah2mVrYD9mN9CxdN8smsf2WKPKm9rS
8WVJ8kcLUebx1POF02F8dbD8x8LLuTXSMl8V34lEhrbDkYkHwS1S12+N/+lA3P81VwIV8cpjAXeX
KI8QQKArbyif+TXZSADxbkWIK/uiDss/o+/ZdGqE+aomvRr0i2Es0qHuZeBcP/ZpNfQtgUAQa5Rc
Eu70JWk+VmpcAIASE0g9LaJn0w5RedWYb/jPEFJ9w+scqAjWV3Cb+M5yMkde8V7ET8fnew4kTD0R
I8W1CXzzO+lJXI5NHS2i6VAFfLbhNZt9W7Lao5vowkro5yKA3eZATTxSJUL4mM8/bP7d/or/W4FF
JQw/43y5wDtIxzbz88raS94eov8XKv7y99M9POcHljh/uy0tbKq70yrhudkZlfaIjxPOeq4Jihdo
u2uyOuqMgprvhGomWqVwmQvyDVbxBYzVM2HcLoN9/QHVsVv7MAermbe0rOf2kbtWbjYhQp8X0z4Y
0vGWk2nydZAQdqLF6cZ3o90NNbAqb67sry7EQV2aFokWd0Prt1cGePzAuBbu0bol5n7A9NLa8e9I
dyDWC3W3kromJyzP2zO6AADLvW5qZd1w49QL439HEGtaL2wwFFDBVk9iXr0kI3+xgVB/8gvCLRoJ
6KvfZKF4+wAwbDtLke3tA/BujK14TuMDSP8zdS/5Siu+d11znRTOXRac1kaVOTaxZ7VnyKe807WH
WW465JJY+TzeDq71qTXXqsSHg9pNCYEK844SdcN+l27Vigf3vcfGQbv9Yp09rTX5n0PSeYfoY5WU
VZ8HmqTwhSlyJdgirPdIKTqB0kyJPkO1J80f22qEpoes8hkyZUfNTHVSs6NwEavzzC8YCnL/b0ky
3PMcb+R4UO0ODOT2YvTpLDQATkgHU9m89OmWhrDvZYg/zjxz0us3wts9Ec8KI2FadisdMbyJ3ENI
0EvJ6eCqzTfodAXrx0ZXVW3k1RmJdqYT/lXDFz0Stfo6NArNWV5NPENgYgSahfrI++fwE9drFHm3
X3zFjmMFVJdRGyGhcxqEoJP7HJQcRuu3yJcp1uECqAqsQjmVJzjTSpGHv/+DTMLuFMCtGxeBq1D3
v7Y+J2/IMP/n4LxYiROzJWbkVfI1Ho0ibySCJBk4Fz4OJy58lro12JV8T58I8xbnUfUoTeedWshP
cAOI39j/XoUupXNeVy/e9BKj+wFyM8BoHT2xZi/4VNbM3kKlE1Vo4qAbhZ1BK90iZSNJ47B5p6Ev
H2IP6Jrgt7NW/9qaf93EXaQUhDQMIZxEXBowp/ew+qAQdaLgxVxSFn8vFEDQWk607qp6UX0R7+tH
Te0UwGRoJQjKtcLb9IbJ2YRORkUIEUaQXSSeCZV9B/WwPuXS1htHXsXGiAsNk05kpH5uNUpBmR9V
8aNfWxLLa+twj5No+KflNlsgYD3kd3Dfehc1DpMglwOVKWpry0CnncM/PsLHasw6a/U3t6MuQ+Ez
wliojqXWH9vWlrmFXau+TgAwRm3uJMMgctDzs23jL/WzOkqDX7NMDs0NobeJWza15K141JlH4ezs
V5O8rBh6d2jnKBc3Hc6SbjRMeYNP6xbM2jvKRa2D+x8nr/4La7kksBcLY6XRaCJ0tJHmzzja14/8
9Op04MHOzA73libpqL6yIbknvz4ac7kuS/PAwi0W0sfzajnpQiD6FBLjhfko9+wPFilgoiPLTw0/
SYo9vyjwBG4/kp7/m+rZWH1Z2hC+7ijXRnIllgxHLsUHiGKEcmugu83gK+koV/wTfWQGDWh1Xtkr
J2c2P+GEMYzu5qRlFmvPop2Tl0VpkTb8jphg9g1Ulku1XO6WWso2QfEwcXzNsnSI8aT3iVBY4gJ7
61oJMeYUJ/uhzcG9LagrsxT7v5WJbdORDEfEqYSPH5INiGrvKZKqgMQgpOJ3uiYO/FSpnyyf6B8F
HwoeqFLeDSLocGCea/r26iZhia3CoL1nGUPTp/zFLX1Coc4t9h3o+URSV+AvHMCHv1F49KntfuNs
Wxts6tK//U/b1errAX54ANEKq2b7KziDF/5793RWCK2HfkgDXYOc3yn4OkWxCTj7DL3o1ICPtTFZ
DWwcDQEPzlUccKo3kLLwH9U3xO8sj8EXG9UL09UbnVLFqXbTnhM7grc6rw88VUtczLuBR2iHkaPw
RZgF9bBZpIkiszP/2m8c1G9Q+Mh3gm9bX0kAhPzI0Xle0G6OtlE6Xu9ZWExI8g5iRL+8VejIjq8k
WuTZltk9Wp59qI/ZXE/GyHIoD+4Gx0m7RHSwHhmhPiqSuYMelZ01n02qeaUoJsHbKwYMXOwzicDE
cdDt0cbcDbLd+ETXwlmNv6MtE7rfaT1fRCNOoaVkT4jWKWAYSg9XqDOxCcMO6eitckSyqyLSdK+k
AlBiU6AB0Bo+Ft01JF7MIvBW0qLvSutWEgcndijbiaM5ZvZY9tSR6BaLf8zJxvhS1zXCYlqZKoPJ
Sx4kYa41gJ62upLYDa0vKTKMYqnlKEiuYr2syNW8fbY40LYzObz+xCa0APZ0H1p8RKaA83K4uLx0
OYFCBqF/Ma9pzZAp0FrSWigGEXY5dOnlHIeBrxBLbaq+V1tlAidnCsq+6bjqr/WyI9QVRpmY3exO
UNiFP4ILjotF1t6OEUxC596orGBeXx5n6MMYshfx+faYzusU4KJ+OdgN8Xyl4S1tLtd0wwt0PWuO
NjsQ6QXzRUvIBa6AeQldhtJEpR5xa9Pd42OZFzerIYWOxTeo3VqnfWLNtAvUyQQlq0P9m5+06qOz
Oh8/py7m2THOFYjT57F8knAoLMEIZVqfRcDONp6/Dnl4JQ2tGGXqSnC6zgAzcaCdbLlj/pNPnBiA
jytGjQx88JYzs4Cg/bBRtSvwIvZYaaxApdwVYgSKnUm3alUCN5G63op+J8FPRTsYYgw4JROdH7hm
1/rgnCR+D9uj5pXAEurHE8ED85GUE89AZYGcoi7lmhHoR24w5VUMm+GQOz7mlCJeyc2zPwYnWUuj
Bt3sQBQBAb4Um0VSxcfqV4VG6R+R/bmPXrnL+uhV11dnJ3YshkDjxeGmno2+6xV12VokGcyuEzge
pEmYgL8afcjA0VOLwSxX/v4sr7J4F9ReySej7Kscj7x3y52f5005yuzA/y/Wl1C8oRQysbE0o6kZ
r8PALw08A0qQSQ+5Kxq3X7BJVUPY/ZxmS3guisg9hPltgs/mMdI5KC/fo8Arsh+JyjnYrhyYZb1j
RJETvHTv++Lb9O7vrTF5JNbczi9WlVBQj0leBr+rHcgOVhRlGj5pNYsj2RlXJdTpsV5xyJXoncRR
XPDq70NWL/CNyvKxzudSXj4KYPyeWPnmYW6ThmSXkBNi3637Pc191yqUDEUqUP5Vo28UqrYkx724
+nYlqb/Ld866OSx+ZKpYZBF88QeRnBYZuAfpkwhYTQAmsSYzPIozmweuuXnT3q0rRnijJVYEwJzR
Jz63nBdMvRvXy3Tj3veomotmJxEzy3gJ2eeDsH0ls1Myc24eZokmQAAAq2QWCzEEDcD//eIKNxMJ
RX1U6V5RQqKfnSFnQQf5ivJmOGyCmx2RRxR0QGNJQRtjuRbMgmeq+2KYtWFGf9jlwnsZ7kRFi3dS
OAsDryXYUfNuO11a+wDwHEkVRW1y2yXJ+1wYwjjVjuLCApEUqWRm7eFWvk/tLb5ad05A0FrgEHkR
pezwZC/lTe0/AAD6il4Pn/+W4jEtZo9a4Xs6sCaSbrOoXHOMmCANTZ2pD1H4Xq94cdcuYktgWLp4
1bFoSRfHbDFNoAlNVIDgP7rmoBXNDyydg4i1Y7kpJHk5JgRv63pZMHKG9dkd/HI6UIfNrJkXu32q
MznFxDXqLsoy6i0Mztsz+p9ER0aDHk39rjNcWiEtKJLgdDydmSO7e5LkeCKvkznvxzpc6lrVRmsy
6zNXOAF4eUOMy8AFkJGaHevVqMy25UZW9RcMUgQN4V2M5lIkJ2iu7QBZ81jJ9XY0XEGsWVrHdcNs
0YYkPKaENZZ5SKjwuHEh/kp247TXl0h7UnImRR322QZbdGclWguOSUMCpPaqcnYZxapA0AwVhHdL
YuLSfgEfUqbLd4VYnp1j7hsr2zbbRVtzVLEVYJdVJgEQE6LKCD5WBk5FqcH+jtg1Itz4432tR2yz
khzjQ08YkuqXWRzNLK6rYb32/QBMz1IOD5wVc8oQGOAnpgotpA7wVxCBixkxbDSj+lRsYQm1lHsI
JgHO/rkgipgzPg95T+oylHo4zgIE76NkrjiQrNUfttSJqiu6RNCYZP10FKsL6qLjDwtBItN2A0rG
oGnqgIG7qUpMAPifjI4uspkXAWC/8P8jyymNqfyYTbRYQVdrgSOW+DJLiV0IRs61W3nCcjkzL2dI
ECHg55j6BhLF1Snni/WIeYIjCNdld8DaskpSN03wjxm/IQnxARnl/1c9xFi400omNAAVH5nIC+EC
W8y4jhRY3Xhl2O5aoCiA2F56I6MpJTZqTjg2xlaugzD2FMx1U1Iq2pRUy47N+NBY+rUylKvhD+jX
5NTmtTdfma+iHekA1f+XzdNhAPh4dz2AUIYE/gGka388s6qs6IjQwmODpFlsx+01cpfiGJL6PO5P
VEPHjvxF12rji4kIcL5RD3K+2kXN8ZBBzjlC5YVvNwUsksDg2JBhABAdfkGKsHk9vScsUzMXOBJ1
sdTOB5wXJrkuICKyW89KES9xiTn6dXNcpk1dFUDLiPXos4perRn2fT6uBv4jZz8DQ5VZLPfIgYqw
ap/lM2p1sDLclfJAw/UFAtzPwUE/3woCdbC+2/NIU9cEZl/+pv4DYsmQ1dI5A3EeYlEnnK7EGL5K
3HQzhgY+KMoJMWJcJklLW5WL85unGM14/5VUbxfSsAWYk8XkOhFMFr6bV7cipLQUzAV3A8p9Mk8r
tg8EX1NZZxeM7sZhNlB4I/ZdyfcqciPrjOdvEsFmfv9PJwg8CTtXYR79pqZBnvcd7dEGtvwfs3Hs
huLiMzFlkVryhhAOQf9/6NLoH7Z1WHyhGcpRi7aCcQIIIl0uSskvxFqMgN6x2pQv/p/SO4H9kDFI
ADZsf6MS3/jv0Lkh6XcRdHV/bOj8K+FgWsoAqPAeJSiu7JMaJlg6LSlco25b7G4dZFxbFaxVVl06
vt3yWeg0qnjAEBiJEBw5GpLilKD2ioSKvRDPKCFv2lkZM/zbRFTC6AmlhpKWyQCZ9Z3xcJ+NWCVM
o6Lm9JlLKUK3iaGjKHPAxHkYj1cjoUr8S9lzlRVGFszsAKn1wei4juD92PLCuWvS9g3oGZOZDd09
kyO0dLAK83Yp7hLONPDHUYP19x9Ppaw1ajicVRM3+sDdFJsO4YMB144QbLvfdG9ssZlJdmHNOqWS
k/SW07Hlc+qWxsGuztFWXDUHB1cj+JACdaowlXhoJ/WsjseF/1gbJf4YawfZTfYFLm5ZYlApj0Cj
gbdT1O9kwFONFb/+uC8VJ8Tp4Er9c/2NP937ubQRILQ0A+/EbQSryRsci3GfvAP78iJ+6/FrlJYT
7+RwhNIHBW/bwYBisKLWxcSJExuWrv+j6ulNVasFPUbX2DCaRrMzjp2gfCpRKqAt1H0MicmKk4aK
jvt4j6PH2vO+ohlrO7qGQlcz3GANHX0bAkAkLnEVgbUfzqxsonYmv5KA2IkGHF5eWx4yO7uRZcnW
x5v/4uV3DInAcBDJZ3enTt2NAQ3LJcxAk63lnL3QhkGvXZHV0MzhIU0o9MkpXrCMytPX+XXZe3Po
nGrR/0WVdsvsOWy5CNAttiHi6xLBM/FW5x70FiszVbc0KWl2KkucvJbDWt3dAA46Qgi+jZM5QnJB
SRjMKeLwec9sUqOwr5zhLkHKLQi/ewtYgITT9wH5ApSiilHbmZ0vVviKR1QYTI7wRl08d+ZdEV8e
T+vl6jv48bzICluO7tb4P8mmgMa34HHoE3HclfGbf/EacCn2K67x4Ygyts4iR3qXas99oJJx0fgb
PHBlbOE3K2g/HWF7rmnrLJRMYC89u3z6alY3Xv7oerpFlhKnOjp24moFe12ZSacl3/rEqWq2pWgK
yErs87Q38XAzqLPUBbwwZJql1GWVUwZrUQ1owwP2U5WDY/8WyOLKk8W63fau9YKmR48LEgcLxA/N
NCCG77Ah5bjys1QhvYzJI71GSCT+r1xzruH8sfOEcTApCvxOFcXYAUqeKUmfIop9MJccK+AmKspf
vhcP3hSrBzgqqnXz+YI2htj+EydjoU0ZgT9jB7ApOhbcfuR3ef1PbP/GfDBdloHDfFBo43elcpkp
OyVkPbFASbrLLtQ5S78t2nfW1dY7cOG30cLIt0c4a+//qWuXuMF4ByvmtCPnUHvtLFw44ZxQOvA5
MQMNGRcnSMaCvi+2aEjKBPTg+7aUS0KRFqn24yGQNauZLuvYEmP4AT8J+bcFy6DBd5tPA5gTcIXS
0dXN74PNoNGC4atEeuJtZ9FkCsz8z6xUT/kwNWLYfsYNQnzZSAZib6OwbojJdb3jSclWnZjoG0ky
rHqnxF9l9TUy13HXAUcrYX3hOXQMFmEYaehVsRM86CXoYygP5XffKddk8rQX3/kDhAo7Fg5yGc5X
YqNO/nGRLCieDMJZxcJKqrkYMWD6yzW/YZdFB4cBG3nQDDjQliKIlpNSRdiO78JFOwr1xnvSQ66w
lq4xUUIyh3t+AyJGIhW84mXRCa0s/HTnGUaD9q5oNpcbiu/ThgOhWaj5Pg2NxjX5T3LbX2inmFjf
BdceX76RjwuNRXWyKaD2+ZKLpvoQ+rmM3cfBR/Jte7XbFTAL4PrBYDS8F0hN7avOnswkZio6+Z/r
YOQD3GobUQck5QM9Lr2/80ZYCcOC/xo5Ui/fjAlmivzHIi4+/mVYdHGmGy/LoW7uj5QmVBBywfDC
MVpSFqSmgvRvjeoDPask+jTqFDdT2Cfjfij7/HCPY6GbR6WXZYykxpoLjP1AM0a2XNf5zx+vRnQH
3yFNF+QAMlzSLFlPkX3U/fK80CdceS1r3TZgKO2h3/ghNvRgJQ/SywROFFuyfd16PmAMA/MYNJPx
WM3hCiLn9pTq0w7UOnLbsIO+0jMXBeSj0FiMhUoKNvq5mF82dFW4wv3xxGVyNjTRjxcFsT4hgPcS
6FE9VGksrlMY9Dv21rlI/MHgW+XXHgRc9iEmqHzo/BP3jkFzivaFjXPXzi7Rbq5zPuoP7OuRS1Jj
jiCsw6z6WxuxyttnqcuFtT4vpcpiGXSHY51nJ1BMmT3fwrg816w32XnLOuqZnBSm5QoBZ9JGye8v
AOBsSi49WA1C3mcpPyXwejZ7TooDWYNBVRr6/gdjPgPLasxSUV5hsmpuoQRxvvyfexcf8zLv61SW
6HTg6en4MfMZZdQPmYqG5aDErnPyzgem3vO952mRP3Mkr6tMdGIYAe0zsZltKdwtndG7ejnwVmS8
Jtn/lgCRhh/5VXYLnO4k/UZKs6Y2BPdGW+9ic7o/7HS+JDL9a31ruPGteNavWg6rlMTWiZ69HmwO
GvdnFhCUNYJkxiLKKPcT9SmX9zLX2Wt9bKi9cMavjL9VtnnVl822Lowt4HOBDsLF5honKY10RTt+
XvWmmg2g3gUWhLYzn86lr9bkYxoHLMUYNHBZdg0N3h8eVBwDkY0W6Vqb1mLUP4O6jGbrn5/c8B3U
tBcuY1zLQjM0IH25O7Bzj6W3ooaIHnisoOfmlaDjQ1mrerWLapgWs6vOWNN1EwDJ8cdeCq6WVvNi
K34yN/46MAN3YcT7AA9E1diYeDWer31SGyULJtJlhhI3hyJHWQGRQl5Gt8Dnf+Blzvu9qixQb6M0
3RU37tDYfwu/MgoO5j1VCRyyVhRXVqLJ0TSNEJ0KN8OIIVphwCJ1Ty4IjGglpZGPG4k7HJKZubdf
yL8OTlEM76r9kdSdDy6u28sWzWb1BaQJl13KdB41mbyYVA4xSZBzoiDR5icq2OjQdBkFJTwlBuec
IbVXO6sMln3K8wIJtgXEmwQ8UzZQMHoWv8javJVSXZ+4zVhHbQTDiuRogqumIAseP+WAoBDB+2jj
sARxgiam+At8zQR+a2TAK57tc2Dc7/rHZpLrKH6zhtVgPVumme6EZ66g65Az4fHpRTV2do9wsZlA
OuBsRm9ERrH4gulTUGNTwSHRlM+AZM8G1XUIxny/WDwQIlvdHuINVeiU2iIoWCq1SPAYvPxmCVNh
ZPeRKS1uGb5/kR9vB+/O3e9f0jUnzpPG2NVuFhGf6yALo84wRQbgzMsYpeuINjmLnMHHYDD6ix/E
6TQHTzTxpyPeFAYX1D6YYhgxp2l8jbPRbf2Dl3sLRlNFJ6BFTiIchKumEsx63ggJgnTcFZiOFujR
o6mtVRtFt2Xk+uJoAKsh2QjYbriPMyq72EJQdpJlDKj0craKqcWcrqTo58Ygvcau0EFBXYSmwm1m
AuCNKuW0ujDh01o5Lqrj1SKebcaEhfas+enxD0RBuRer6MpSYgWkh5DiZQazl2dEgWrscTLiBpEP
FXQz3BOB9dJIqidXYJYgyz53rFZnaxnnKg/y/c0fIWJRGXlaKM7A9SGxabVzMG0ceEMNzz8MI5Ab
D2VVZTpQmviJ9oigZuPj1y7/Aqbe6mpcUEaz7cIcRcxK4OeQ6ZHZKn9mkMPmH1BSek5OsazTC7tE
p6IIlmCUsvPSuDt4I+NyYZJJB7XiwMx5X9u9CbKrlmV5aYuiGYJGlK7DjKUTxdkpQRjKqkfpxmSJ
cQ2vRZty+fjFqM8wP0IG35amX12lR8ngEh/WtpsnOZgjRTFzpv2S3fDqM2P9kOEXVllTG1PUw+M2
04C6keVCCvbYCUowHcqh5LLNBEXrVD5fjULRr2xSThRzQaYtNYLpN7vjUfJGG3xWLKYRynDfxpkx
2nUz7XZQjsCwp1MSYD8Id6/hTipNC92UMlFQ6fu30EPaqLqbNpLAHmUIhEJz56YFcBJM+jWyFOPp
NV5cJiXUHXLvoDZJQcau5+kt8ECjPwwCixd/6++7EBeOw4h9MBY8GKvwIfCEd1t3wYbYGRYib5Jw
NZGcEC/3pmgaM+AG5dc3qiPm/mNPuuZFAppK39gNGgBvFRkmRNdI4TWrj93GYtTzfkBWeulrFIMl
J7pKvBsTCYhTjl+kvoHYZRJp3M5YRJbc2vwPKXLSfhiQ3IkbSMjFkdVZ79VqKFZOVmc6OL/xemOj
A2P6X1dTClr/f23sJbijWc10tpU74sz3aBUBwgM8IyW65F6j6Il2MoWjabL2mtuKPG8/rPVwOiTu
EQ0Z1LrvRh4eqT4yThEBUFfVFAcycZSSQE9k0ZVoT4R3fHzUjy3zuj4MkvYUwSeEZEpdpHdv/vjg
Jwk/7AQJM8scLP2FLtHZqYj0fdx8OV8B/03/fRQCAXQHbT0DMNLrjiiPtiEr/L/rUNwNtFSYAOl1
cPETVzDy+dbvfUhH8Rz3iupg2vrjyR0TDLP2NCx7Y0ABhPM2VvTuJWRr9yZndF6CL26CMtKFbccN
NQ1mXnGJ9tbistIbwqrLs/A35P4DfP7mHlQC/kvQXaxW7ZR5kEjQm0OlMum9eZ2i8sUtfk/vq7Yf
MCWaok6kQgsXShkw/57nIFrN/D6vyVuOrcenfMU82wsSjd+nv1MiRJMxRV3ac4xdgabPuXknE4EY
d9IV2f154CHs8v8nnZgJeWibwvNUKiYBZ20AULVtEq5oZ0s5jFxBmRAvxBNJaPklbpi9A0JwVT9P
RrmwU0pK024txidjJrJvF6nbxhuTW/eP84wQ/xHit2P8RqutINHSXimdgRSGJ483By8AjSgnBZC0
JTD6jgCzfd5IX/PN3ywfrUmNtuuupwsK3LM8m9NYcN1HI6z84LLzMIEh9jX/IPqdtkeCgTdxmWtf
GLyRPwU1WfQdPArCfogdn5ejFyeZ8XLybs89lLof2PMMY0QMEh27PEjWlz7S628SGsnz7Y5XOfVu
brasvB2aVWDf5Ubk/EzxKNvfUrsksJTWPu9YCUBfdVFfzxTFnjzeW8Ze6g/Rd4+grhnBYhNx7Spp
Nq9xMbrYmH8gVo/vozIdcOra7qkdmIsEhn9M3jUSWgjJ7d22nTZHHb4BlFz0uLjW5ZCfBtxS0agC
7bOkxjt2t89PcovJXjfvmO1oUJdWfHX94/dUsLISh/5KMSGNeYVSOld3I7P7U1Aqd6Lv4l6U6d/x
WbfGQHF/0OjLtOEj1lmPhpC8lrg2j+S5Z75eQyoibibMeijR9Qy7+DXOSb55L7EmN6lauw7MVFeP
HAj5MnzFJeJ9K69yHDh7dDkav0y6wGcF5K5lcRrkUV4uT2IcG8tCp0ioFbVZOiayX5BOcBL/BfqL
mu/K2e9luLYSSYDImU5g327MOH3CKH9qXUtVgqs7171wfRojh/qE9MHixjSOX8DxOgNaiU7nCs6C
wcqE1y8Njm68R0NDDH4QTsqISz3W4uzzf108DivecuauASYEu0ljbBK2599jLyulHRjt8eXUSn36
BYWrad89g9NPn1o6qijnvIWEaGQFW9LnKw5bD1F2ql/L42ZWPQZea5Fp0Jt37h6jWJYRFuyAmead
sMoQ8FqL/7+3WAKUGZeDvjiPMWix0ub8TI4iloQVwNUqfB0Ag2VU7NYF9cH0jN1hfMqpPGtQWgiz
8q5ZLZd59HM5QQbr/n3Hgts+iG6kbBLyf7Ge0/vO2XjBc3NF3g9nfReKZNeCxpgyfwAmpO+fByBv
+ycbFnOYHRMTZA6cmm3oRi5+XcDOggVTQQxTVqXjIx1eeqPBugJccQYsWwqkxP8UHeTlGJVxzoIm
gzFiPSNqN0L9cZktq9JQjM86j9xLknN4Qg5+YMjFEZxwODEdVgGsZ5CRsH58erJZSuAp6yddTRT4
s5v1gshIJfXRcT2N7NnVYJM4pQIIGoTKgC74z+0PvMWypQqI1KsSIJ1QRQrElRq4Zf7vit3nk8BZ
45UsZ3jLuw0bB/QN68v6k+/zrvOEJS5HhmfF/QFB6EYUPgjpX6gJx2QqtIvD75+Rd9IyhKQ7h8TO
Nti0rmK0Hx/gbAirtHAffJUxFNOc6lljottXU1PKnis0IB+nXOcuRz7nijT/p/OXyH83s6G95A6u
Hf3HF6KoWlk4ZtWZxQaS4mtPFY0QMLi2oRZlfYQmfrKi9ii59CmveKF5kutX76/T22ztmYs2ZjEr
ydDlIVfSRHJk78mEHiCs1SPm6AboxfqLA7b3N70wbrs9Hx9Qbs+4FEqShdTqGgnCm0TwoOa7+3NQ
fYGUuNHt5QdCVjffCYGkpT+XNs0z5ZAZWHlBgpMQKm75+K33wH5Y+3/7FQcHVWtFHn/Qs8w9Dr+6
FkXW1+bw+Pym8Advye4YlqtR1ci2m8a1QylJRdLYQUJTCBe0YP/GjMZdjHkbJaWRlM0pRcXq32Xk
AtSd/KR25H7fRJp9mwvgp3Ua9Wv4MK0MvAxYDu4Bz35Yz6q7/HSPM89blDnAucjZBRhags9l++Yl
8Z8VMwbozmm/gmk1F1ilWByn1+gIddwl4gRtCnChxcDxIxyUchmxnrMB8k+SeSGFIQMfhUQaehtx
rLHAcycq2uwgR9aEzSqSIvapzly6vBHiQL4C1BXh5VyNZU2thZUQaSSwyD3SruGKq2gtUuqXW7St
HB4qW1bX7W1K5CHS1Ew31yXAQzJL9zcv1s1rBDUawTt5tSgCkX7Ck1Mo/0NhlkjyteaRyh4rTLhA
GDwaQes6GYV2Ri7IFODZY1sQqlhYPpUBaTKAeioHjcYhw9B0YAiHWgsJGoYMzrhFCjWarwDxHrC/
1i8hbSDGtUGiEvU2hvT2WWKhGYPjw9ESRe4y6nq91vd/sx+1TxWCK1BqT+/5nQ6iooSuCXIdyDH9
XBtRhiG7/3u3eC5Lp8jaodk92IREroCYStoaru2A2jTmUI7VPDRWyg/EFwoRTeJJV39XawMK7nGV
pleNkAcqXoAbL1QV7w+z6M3hyras0fctgkN3Aiqo/Ek4ZxLo5xcPIFDPFRvmAc5kAl41FVhRkMzx
JfQEOA2lKhoCXBcc18ThWq/rf8T2oYBxxJX+b2/vfFJxSyL5VmIYtzCWKYkVctw9gxfvJN6TjiUv
qjCzfFK5zoVLeozbqdiOItBFi3D4LSe/psFkj7HFtyk/l63BSP5KCa0gv5uQBwz7Zog9lBR+DnW8
TI2ZdNn7uArsfXiNPbX+hNL4TBxjttnOdn2+S/6uXNOdGDuoe9jMlQYDUN+zeslfFvsjJoiSS24P
8kqxs/UU3AgXlKKH+MtTzKXzbvRmV81y3dx43Vqw7oBjA5PfeFHX5eahXkznot/spS1nRxiRc3rj
8MZlUuacl6+0djP66tGhWSkrM1EkDFZaOIkKqjk716/I0nfWVrkeg6GTEDz0xInRV3AIiG1oxKme
Lo2Zh8JYw5lgyftpjtiQzsyuKRe1AbKibaZ4ME1ULHk0/v0pJ9UUeHQZZYh3UaWE9i4qONjGjZpO
P3BtMKZF25ZwJPtjuwIID9f0KyT3U1vH44PLXdOLZvG7sobl4DmB9mrTtt43qhIoHXCBfI4gcUk3
NirVAotm7pYwidYtQusCyk4Tj1mTiAk75x2rqzRSgIk2Yq5/9r4bvkyPL0LFggecPp0P4LCxksD7
3eQoFEog2EeE/VKtKUx0h5KcDa9nJm+sQydtNYNZA4WCW0Lc0rhCK6bd8NjbUY2iH4HML+CAaII9
OjzSyXWM4Lgkc3UG5+VAHvSQVr8XpKY6YHTeSB/zwgmcyjOmTIrTk+LC/9FD44xAuhRR/HNWLJee
ly5vfY3di9wtXrnP9YOErNOwTs/IaBeUA+SazebrK6EgP1PSZHYt2vUf1RWQMAnqUZ/YgdRDveXp
3FDeoQzwi8pTqsCCjlC7NrcErkuvX6gR0o3sTOUgflD0hgUCt9v/cOSbHN5eSUXzOlKx5Jj91wXn
5GWfOdPhLo1qWchsRA7xsCrWimCXsUXNnDpNOwzFTqedIoIPjYpLTJKIFC8JBDdUHWm/ldI30Ysz
xmvmXrMyIijIq6NSkRz6Dfd2AwbDHgh1cArS7tEsBdLHpnHYoTh/c8mk1iQgqHougn4QLD9L+kKs
WMQtetBXKTVk6joZGSX5Wf+FcYA898effm6KHbiTkFUISW6XpMuOaLRivsbxK/fcbF335JsT4qvV
im2dwmbllJd+Z7Uhs4m/gFd2xwJCX02LPOCeK8r22X417WRuP0wdxfkDj+2Yu5hIrDxFIyag8n7C
IafqJE0PawNY7TAWzk0wLRoqrTo98wFECKYZ0/X0IaUpLazWrU9m/uj2PcGsEao7d5NlD1WGLt1N
D2NxuBBWR51tOxkQT6fSQ3afly4j2vlKMuRVz3W8H7AzrYJcj3MqKqMawnkpblPPZxZFoxoPh2WG
mN+7dX7qnT0AXsJPjEcjBlaCoSZ4dE1AU68utNtrqJKfhT4lb7Z2rAoSfE9qBQiPgvkD81CjcD28
4utch60FGBeTEZMGdrNx1svLc11+EWjmiAbxwp0c4Y2gIpbjOifCBmfxFhSpJEHF3V/6BLJcwzFQ
iPAWugTQ0oWOvbKKrHoHTBsHgvyPfd6u+eh+1SSIMWV1dKj+3KChq5I0ud7gEam99+5FHcDM8F3T
EnlaiCKIAUap5Zfz0iCIDl0RIpTCKORmriqby5ir1YH4EO3K0IirWY+w039tiQhU88wksIDhsNYJ
VwMloFKQlWymB3lWBlqsl8Js7z3JjT3rxWS3HMm5wxOlBOEyH93g8DsP2soU1FuG0viIuaPA5em2
aSffIe/mkj8mG2kLTfFZaHUtUzX8jSmTDRIkZFf2at8XmMBjeTVchdJR6aolp3Um6o3EPtQryyaq
f2j6heMmSZu9jdSql9N7XxCXaL/ez/TvzqMhxX5izJPlNm1P1K4EjLEi+xX3pjBt1xLvpqCKGYFU
9RqL7opmxLdRPmuA76E9AhpS2pDBQX7HcJkAVV9QfU5CfKAm9GVHn5GYD0PmChrYUPt83XS6EL3h
bZxMfRuk19Wt+WZc0nDqiUHFWwv1YZ1ltu/Q12Z5FDQUboPgyM1fFy8g2vTroxSBAL/Ve4Hzh+B9
k+h4ze6qZfkIRaqk2jZPsmqd9f1DYFDn8BCRCYD6n+46KQN1ryAEHYi0yVyg58KDXrcYCSdxZiqK
WUM14LDL43sapL47ww1jAMMSZ3tHGXKcyxSd83sndC8MV7cj0F6FgNySYqBi0xXjZ3y98IXJC9pb
/IRZEdxtJ2jxNyLoOy5yyRwsPdZ/+Pylj8XIcviUWI1alNOv8puKYaCII0LJ3/bGAepTeAP9ERBc
GT/o9u90glpbYXaNo6c/RtebHwilDkElSokmIyRrR532YTL1nKo8HrLTNehn/e/LSdxpezlvzGY9
jVSMr0w49kw3zFgwl/2wGD0Y35X0tbMD+B/2uL4QBwxgJhj27bwj3pNLQaaLBZLK+U+FDilTJahT
HuRc8FwVHvHv/79jTrfo+4s8xro0NtD97EkMMZjKilPyu4Ha9V6VuCfxN7Q///utC03NEbl5y1+h
7oGuei6XfwWxkuF4HP8/0d2Z637Cj6J0yZI4bgVnKEuxiACJU7+fpO173VA1cClOzaXZBXXrzRuB
HjbZKPXzmsrpaQh6tLKAIhvXjReNh+byCosOcutb5Kp4R7D5308wHdy7AdQSd/A9J3ySuexxp+bo
1YYUksyNXRinbXQ2Z+HyzBxsJ4VQfrQ1hIl8HPbU4UxIPJsmPrWrp+ydTin64pblbHBjylX/Lsg9
WcwpoZNvzyb/6s7ze0VVM3ZV2e0IoCVcWwyIkrHCPrJLFh8HGgeU7bzlInul8XIWjw2ZVSYdT9Na
w95bBLQrRfFiOcvtTsov7vlVWBMpEhZ6C3P2BrR6tJIVij28QZvxj8VwEPfxvHh+ZfeAtl+U5D5L
moA2yPYCu0WioB3Nhgb0O4jg6LdbJ0RdwP7CEN6Cv9zh+qq4RhPRtzU0e8n5qu7fSYTgqt9mcSB+
vEDC/wHUYqWZrH++DgKg4PYfCFJk5ZS/W9PDgpy9WlJ3Agr3wJ+BdZN44RGCst6Q5Flh0/0K7Rbt
6LioXLw9J2ge3IBsn/6vhugjjTDcwqMMc1q8OFn5eQB715lJJR1KkXDcBr4ihauaRbFw6NIjtt0b
siE79UtMZfIYir7kxhv7Oo7LuR4XLcLUZlMyNO8ESszZPNYymIS5BbOXx1h5agsu+J6SAT1JeG+L
7Krju6plu6c19DTtNPvDBN4l3EdQ7Mh7TTHg1k9na/l2V4uHWSfSMez71OeM+KBhIT9MtmYkt8N9
EjAkSz5+6xIfyiGLwp5gkU3EOeAO73RbZ1RNviSisInxoi8L4EuoODX2iuVyfG7FAjaeTTveGpc6
UTjKpuOvE6TdeB2xmvATKzvQ3LEzeNBarfNA5ZWQBFQX3gvQ3YmSR5ysZstBULTZNZTbPZzHANLy
DoSQziNrzSUkACOKbO75VdKqczhOIyhqC+MCcUH+yu7VNkHG/9PsBnh49z6VyVLxFhTTcxij22d4
DVublUY+coRtHYyj5YscyvO+mOiu+2I36PNYdLeoHtVfJG9Oru3DD9WvK13Wb1wX7DaJoHuaNk+4
MvarMFqP6r7Svg97AC1xIm3QioyApMYqCiNAcRnoFIXpZsYj90zDrG6/SLns272gFt6rtP17lcGH
4u8c89dUADvNl5/wkHWWTcSdH7ftxmGhoGp2OQM1zk5hVR5pZe5ONvyWwSvyDBXvmHSldbqrXRyI
diC0cfqZY+vgaGYhyk9u9oePzHOa/huIz762mpEPbc4ojiIH607l973zD4byVVRcP1N34Tu0DUXN
nwORHiwWZb1GLHHVXj9hOC36Xofr9PK4DKkYi2bTFJo8S7mEFFBDxGnysz2zIoubat0mjBhri9Yv
OIAiAIaDfcL+fQqa84muzEwN0eqePfjHJJ2ZHO2IXKfqdlIgHppk0wQIhkmvojE+jT0BzY/JlAG+
bT7ycfcEN+6IPRmuXkgHnYjf1iQBbTjTdZc3h3qSPlYzfKWqQka2ylywyBH7XNzZCfFhqL3Tv9az
Vqsb1A4lNO60deaieYQhAARb/S50tjAEp5zm4aU7lFuREMKpKSZB0c17o/ClaTFW4mnsO/OyLzo8
NGgQIMVEd+y+VqKncWDaGKUvwptGRab5SxGEP3qmE+s60/tF1Mfm2hYOArH+0o5DXJyU0U5CWyn8
WZk1ChTokNPYpzfGUOCjGJsB/jrCKO7pUYVUbi/35r+npzMeaKlAsHhLDjxDcXaQ0Q2Qdia0/iJT
15Xcue/nhPCkxb3y7+SCITgb879Dn2pT0b0FnUvKSJfYZv53ERM1EX0NMmL+JajTnlWc57TyaigE
rjXHjHA88eSaNa/mq3KquDzRR4/+gwFgWvrUowXhapxkUbKf+jRBxRUQsXwp0wbvQmgI+J/nD9hj
Lp0Gwpeb4dKF5dSk9uTSYhXywzn+AuRjVQ7DMBy2gjs1QgJ+NYMh4TFszifo8Q9Wqe0mRkBPZCFY
ZHp/S2PMn4o2FTCvic2NAx6tKK2tqu3h8H3B4YUti6weNk9RkBPKf4GDMCIJ+4HNy/L2yEW8NtID
8BqBGqkIcHf8A4EiDc+boyCGDF2suS3iBUhW6S8WO7Gk4uh533ZZeCjL4alcyc3N7vEqJ1hSm7gW
mzmxKhei+iCWzOZSTulZ4IGOAPWrefo4lO3BjB8dI8HsjVeAN7N4Azzq5z2bdgh7osChErsg5YmS
atdD6tsx/dvL8ZJPOHn889rkHA7H1xGWFzJ//haI6IroKLgfl0/B6HMzagAFMwQAKLdiG7ltgIPB
y4Hji5GgmYq0WfUSRU0y2d5B+nsv8fAELwA0QFdSMLpawinSY8+2GXWxwT27mTb60uYUSxeQ+JaP
B+1YZ8VLh5wDua0W6QkQ2XaMZmhqzzZLP1ur2AHU0CLIwFO7ghoo6yAtY2RWUh4w7NncWmU21Ocq
6Ja0UX2a88MpGxUZhGEuoDBEqD6sKmzEkpaP1T5VLFcB+qgoTdRcfjnKa29VihaHR4v6TLWOGGFc
j1YnZ3a6JkxoiqmHPb2Q1u8DyaiOQPuKD7jN3/GHPwxBhs1uX6vpTey3k8Hpa0A0bgOhPeeIxg7s
wguzi1yaz6/UDQs8TM0FOjAoGs4mHPQXyfJrGIyqaFPdYkUkSSPIP+bSKWcMZzAjfUGo2sTMhGPx
DHBFjtE33sH9CLUUW8x1vR4FDhZHd3TuPRqlqRsHnUWmCkcGfDwKU0gg6Eyhi88FERSvRhuyJ8Dh
ru8qhVxlHznyFtB8DT3l5OggePcK/TdPLhCZSdcFOUTlYbZQTb/PKOVsksgl0DBs76FyB+Kz6Cbl
SZjl0bcvGwYlV1CdIKnCRFCdp8Q6nTc0q1Dyvy9fdalOANMi0McHCVUQhW7zSC5E02LZCoEMxao5
b/us8nuFLDP3cW9TIKQImmS3KJEVjbAaf8S65Wavf8XC7T9YfdBEMFb6JKIJXYSY6PZHDM4AkIxH
Qfh/wxHAWEpbo3vIUzRsUjbDMJRxsSfVOkluqSCvVsiJV8BmmXAqFdRPR4Oe4qDjPADX6SjjecZV
gd2uW+Nx1keCoAierBvq3C/KCOXdG4Zs5E4VYHwu/vI1GhPWKhRwoqqN+5ZM9VGnXTiYWwUmODOB
ADMQqEA9SzaieqgAfBHpPBgIJ+2dYoyPkEmYF/bJLB1UNfVRt76ck3w9qHa9Clqw9dfPnNIlyiZH
+0OD3dDsIeGmiMDn8FLPWJ8BC+vgw/kAwx3qohb7mBUPc0yrON9860uuhCdgWsRPrWuRUeij4FIW
iOXhbdQd0I5lRjrRLM00r3qUd7DB4aWOOscLDyZh4rMEHTxLymHCAdiUts/QMqJBIEVFqC0srKIS
KIuoeBM19jQuIO9heNP1Wym3/wQZUFbyyRycwGETZOqlGPgehsAw5PE2JEmoEaLAnfcY1kPnDKZ/
va5e74Bg0IkaeIKKRMq0AUYyPLMpnSVEkkO/MpNdaxMO6YsNXp7EYqu4i99xUc9qcY+f7MjyDUuA
GWW9x/ZkGnx2sPXy8amYaSfe2i5j6FOEvyoSAiiQYcoTU5AcRTcAtWlBUA07SebTCZUijD2QO4UM
TCd8rUkPbwkUvjpK9obkuRUtCya8rPzijay4XopuELD06ozlQlw5DwNmttQCC7ynr2FE3KZkgIfo
Oo6ITptBwNiQ8NPGBF4HAL/U3cwzVnve5ZTS7yIaVxNsreslWbwjCLb/3ivgM4sUCwJ2Dm6fCCfG
e3VZAuDPeY/vxkkX8u6M9p/f7UtWMfNnx3bTEax3gM6YX6hjcpoc2mRDyLI/0PDgriGxPO0nsVwJ
RW5EfoH0B2/8HmdISZFsxxEPVIIbhgcKjdVH4CkkqPmEnLOG3Ds9WlPGxs5TJdUAqhcdRAcq6TAW
DYuOHcaS8xg0iVheAREdmsUtDSKNz3oCyw+BePGjziH9LZs6fTewwC1jyGngw8svsLwfxIoU47+f
HouUFL/9YSNaXyIQ2v18zygDzCvd9i6r6IoPd1O3VTIQu7ZUFeR1H8iuPj8GxZNo7A9zdCWQ7QfH
Uv+++roPOEUUFIkydIydMz2487DbAIHiVx9UlZEzg6f+uVC07fddV4BFZBp/kKnIIf9iWP4Ghy8H
oXP0fUMk26G4V7vudkmyFcqGPb7n90DyD0JVFFacvMqSvprsUrFy9m2i1H0psijFGxQzudUUYfUO
skallpowJ1+N8G3iLpIMvqjCConR945ZNsXTVP6tAtFZsKI7V54I4/dHJ0yDYNXcXcJq/hin/WJI
4cEtAIilAgWqeLVH38Zr2MFKFoOBm6Lnw2rJ0XgjvR1WwraM8Xiqu/JPAhwqY3m6nCox4Nei9nxn
3tMvToMIV2Bo/ornIx08hgNxY0WLhOfGYShbsegqKKB5mb+5VT15DxfV9WK+x+EUtkOdaaCoJUV8
u18w2qT0c9FEImJLY2APAtkKqGcXBYKBYrOZIJZ+CFIZcSQI3WojDCW7XbtID/1qj98aQDKXUX35
vXf7On2c0qdAZgMg4j4mNIaLdS67K012NxTbpRuRdFumfDyPBwzq4rObspF32ocVz0YfiBqD20Kd
6Q8zkjOaRlzLiENqMVBVrqA/hx3uxTKAOeti+ggp0TIeQQ29xZz5EeipTnoMKFhST4dGHK2Yy2Fn
R2kIWiBMSwPkJMDAskaVzk0Whjy6MgzHK+LxptdSJGa0kfLRHkD11SCMqoyYQVF9NzSxihHnigoG
LRuBoXUJuAQZcgCTQ2Ebk4fZrXSFyYZpMg0T64Yls+O/L6+Mz3K6al3Z6OJ825S+oQX/QUTZ5vNX
oLa2wFkIM8Stv++cGpGShXAZlCiaqj8jweuthTBJkzTkmHTE3uaEqOKAV0xqTmBxINJhsqCBO7zv
QZDNtWCP0eXxy3ip5emliICHWiVOzR+tYYfeggqmJ6TFnKGDQyQBX4ti9zdniaAoXY5caEYiOSix
jB7gV1tVG44pIz6ltehFLLmQvGVWNel360KJC7305q9A2adXmvjB2z3Ga30gaALpTUAgSsTXBpkB
eUaaM6tkG9tprLCPqeR9Pc7m8FU3MOlpNMIjVQaRpxMJzba28PuwjBbJSLMzY7lWg/GC4hwf1V8C
roHxqfnecwiu0a8CHalQy3x/ZPh1ou2F0rDWMLa/ifwK9jg6SIsLjD6F2dkUiTqSroRDW0gAjR7A
m3XQEKTHRJGpkH+njzy7nhQ8gRKnEbpooD3WvJGyJrPfAs4DFlQubTWGI/v2RXLMByg3C/DshPlE
O3q4UsxVDovJkBUq2Bk/Co6YDX5iKbPNQ4NvlbkA8HXGubm6FxbXHGEbk4Sws8jxGQIDs9dPlnB2
+xjWBTZcPGTLmgYVfLT5BmM28L+gNi5OFWh43irzczXh2D4JqXL1R/4MCCIJaQj1C/tKkIl9egCL
dnIavl0udNuvrpfVCp74u9V9uJuz+urLbwYJ/1u9hIHqRbUANNHLV0bAPJe3/CTYSGTYgIEMR2ft
dcR27c+BTKNqxwZYM+GVgeKdRA6P5IOZzhOfLZxFulurmbdZjitLmjulmKL6kz4vmu+0yXrnxrIL
5rR7sy5va0FdUjBuhnt4B8EarnJokfkoGLfrIs/KBK4kbjT2C02BFfmZbHpv/32L+UMONTfPZkFA
zT1hyDc2t5S2RJHB3CZJRiFYDY0DfL+f9yuFiKDhG92QdRBhogqALNMNrRSxtsA9uputbQ7OkPOn
1Qh7htb0YT/ea4I+o3ziTMfe+yKd2mZhKTRJGP+LC7RmpRTb4TM07pd81etU8l2R4G7dws3V/M36
ztgNLe2cjNgA5NtXbQj5GKYrUXfBEfWXYjfAXgfBm+QF5kOo7KVmqKuhwaKv3vWk12RoCwWs4NMh
wcHCs8LGpJq5TURwkllUYiqdBK8S43FKkPZwy5MkViTZqhrZsdDGbnyNowjfH9PX6xXfBRQ85bny
eiMSdbOSupbLDWYpr969wWhvBKVl/j2UHGXhX1fFmqO3UwSPFIOmXhgu6MlCNku+y6OSPOJo1zwm
41uSLaMOIq3Fvd4o3oDeugQ6Oh3wqSq21fYSmDS993I3DQ1SCzACT+kTbzFeeSqcn1v7ft7X3cme
3eXu3bWwKyW8y+WY+D9yNA+pTBeBmpj4FkRS6VLx2M0Pbotv16x13xdNO9/BfxY5Vgjcy5Zo8zev
sb8yhYOL4tbpYS2HawkQdHlwMEQvKqZKDwX0RCaiuX4DVereUnSvtzM9dvqRoJxU8J+SmrVPcxzR
gNK0PmGZD8lRZPpkWc5BDORpt2X2B7IjgKKY/mmT4EveUUeym5PMHgXylG1xlA/M/Cwx+lhFootq
jhHsTtVvI8NXfG+5gqUAZYnNSqDpiMbIhsenqjjrjfyc03JO36xYPbkkob85+GTV0GPLxt5myNs4
VZxaw8OGPn0Ul30xdcQ95O44pOUn7bqzE7uDfvQ7YtdWifPqMQrBFhHgr+c9gWi1Xdk8RiYtClG2
B2Nl+yQWw+IUIgCNqGB9MbA7U++n2QoWfOtXh72qhSwOzEN12w/cFEXu7mnVhLz1GhF7EOqWhRNh
htwPSE+ipS4rK5laWCkBW9aCcj7z6JZ5xtWIXb1vc7mMT5b0EA+nJTIV6mxUc18+SR2Hr85zqrGu
bjceLHgGoZAwhSWbrzOHbVGIWzc0GQooX6DNFYQ2siebry+/sPVjk3C+BPKzePWBb8c2Gwmsc6h1
DRfWGGj7qOyKHF2FghxhVLkH9Ldpp28470ao0omPKRo9QYnFi48G2CBbfLBneZdh7KxbINtYQVKY
dic7WbiAxZEz3d5Q4Ncg3YjacrGcrIYcLbojIkN3byv/iclkvAdlPWkJaA50JE7BUR6Xic1UTuC9
sPp4I+2tEqyYpptQKK41427pBPJBsCPRDkRwYIp/TWsMzOTS5QTy5ho0LXnAfEdGOC0Gb7Tn/US1
cptvseapcVH7D7lumx+8f7lMGzImDZIRDFiPobI1e7CgXDiY4FzewUP61OWlnIw+nKULg6uCmZir
ya5IehxmC3UA9Lck80wqLxSFv0XbuU2SBkRL3EvF8tc1RS94gagtB5J/bZWhelkm7tMaoeYzV0Aa
dwSEtpvUUVuxlLnnqffZazyaL+xXgiTJPmN/fuYLZEmxgQ5oDrAWmsNg0Kbr2EXPkeKTd9jaXY5W
iN4Q1YyOgW8lXFjSq2/VS/1vBSIMi6Rqh+fiBnnPSppttst42u64O7cmq+v6dEOqEXyba9LimvQt
gulvpmVdV2gT6ggWdl73A9NRG1hrHpO5+4qcmDSvZAUwjjJvR4O8UAoHrmwWTwV3Vf4MPay/KJZ+
cxqqiLauUnEOS7WV7vdIbM0TVQcGLXvNLKPk589eB59gcBB8VjVrbYz59y4S/zs3TktFFv5ALpZK
RDgjeZ3Y/puFnzii+qhKkyxxXRXlYBlOwv84/XmcKVYKps5oRTSPB0yy1Bh0VZjMbydM8pyqC78l
Nvlrg1dC/T1qIn5AdJcLDT0oSFZ7EOOt5Gs6exvoOhqgBaOuX6I4Kq31A0qUQXKkPJDsababGR5G
KZyzbz+s4GXYE/fwW7ShLMxnT0JjbNEJqQSbgMaOsVq+E9+hfvSr83kgf+f83ugwXa76uUmM3HNj
GWueaUUYtKo2kHw+/rDJw3w20XHIJA5D5B+nfZ4UMe9yHnoAFIUwYTgaeEap6tTdHZl6iVntP8rs
v/8/utGQ4lDO651JKazjjqW2of5nxjgDXT3Hj9Tn+f+EEpiP4I74BzdCP4gQD0fMZqo3TVjKsiOT
FQLX9ikmp26s1Ig+4d9yJq7yUTf8eu/CdKYx9cgnaASH9UNLGfBbHD3mBoqdbUMexPVxy/rvJ+uX
nx1/gJAw6dBQHwufCxcPLJAcaCejgnzc4KRiVQGx0cIvBaNGMcZ84Aa612acSg3vqTitPTR4GqFX
tt1pbhOGTNeyHIbdWXqwVSLJBuil0dxSy62IQbUiC2+aTH7XYRj/80cpVeNwTScVd9ODdiTYCUQy
H8DSmDVxur9PlconSS+qDBdco8Ck6kVYLTMe4C33QuM0q3mDEULy/R3wyFPbt6dxL62IQ/TubaP8
7n9NH7oOG9I/esJOAXiQI9Xnmp0VB+Mkg2onl2xF9RJjM4z1v3FMp1eQunpFriRJ/mDn1qJONbJW
5n/xRUFvKeAGf7ZKzJy0ZFr1NgFmiAd2UEpgUa5h4DVMcg9oxakMMFpfNrcPYggoPv2anR0JWoeK
YO+tKqvuZL718n81GSlfbb/aWfcSe3Ma+WshpoS2KMqwvhYairC+uAMYlps2mdltiLG0hkQlTaw/
wOSkAmzjCV9k9JQK96KRwUwYpk66djuXvBYinDbgXp+iE71uxIkquONEmg+EdNvJIWh2ygQtdxtw
D4euVDO1GVBa4x/SB8qI2R18MH2zTd7a9OAln60p7xOcCJOfAbOjLieU3nNNxlhfA1W3dvMfb3+k
vj5kGaqEHUGAVrnJJubBw2TimpmtEbyHF2NXOJr8ad7FYDpV6ejpFD4r4VN0HrOGiPg4/1CJsh8Z
dN2YhEtA1tqsjlrthuZ2L8y8c1x10OeZWrDl6f3KXls7tc4kf7JpTsrNcC5JgaSRUhHcbO5rsCMu
NvmYcT0Y2ZljpgY8iqiU4rYB2vP5HurMOTcnhC93L/hjjKyFfTyt0r0G9mkgpSpnVzfj/roRwHdC
7Gdn/94pY7nmgdYLrKggFKsx3t2c652NH+m+mLeo09ABN/z1TEbFSFWrEgXVgYAa7WWZWH8l1FZf
zZ7ZfOhsmSMWAS47NCwaVBwQE1NQY627fXJvJZ7wlnVoZbbjOPNfz4H0FA2MscALCrTdTvpZ4tAy
sTwnHhbwh5XD/LpEPUzQb7aesRFlr8QA07aIjwE1P1iiJUWFwjByiFeylFBmik8SW1nt7i5xrng1
yl2j2920B4owwPqvTbbvEC8JvsqSrH1jqIcslHIYWdaqdLvHDwQGH6c1zz4kvvegxEJQL9E2FBvr
RhdI5X4VSGkH4E5UffWe18iQPzksDK2lCfcOpIG+6uXzc/re1pygjM3fboT+YUd/nxoDw5Bs37g1
RpjPa0LdmmYCxbqUfzUP1NjmDtingEiHeBBKu8B9/I0h4zppCjBBn7JQWoccEiSeKiiach3u8Z3Q
6V1Vs/5p66xMYlFfo60XwC1ZIAMwa1WBJ8sX294iANbCHxBExA/SDl80DaPq7SJEed9UCyMLKu2c
W9xtkFT5MD4pHNE00GZvTeyMxZYkE3edHCQ/0F8KnG8PtTuciQ6GFF17fM6FYRBSB+vIt+heg6NO
qHzwexb6a4T7bwCqnDHZLfsQU1R1kpOSddQYuA9ZZu+g1EIXFs1ER1wDWl1pVoDbBkEF5y42Iidr
PviCZTKIsU5oNtDSgUs0UQLgcfR0Va4xXjb70IvBupN4kpLJVC7qEoyBRqnc1qrb0f3sqe86Ay29
ANb9SO6uGahQu3nBCdc1agb/ZIo7XB0jyTVZkMEjtRwPcOH0ORbbRSUME5g00ZHq39+abuMIQkuV
aCBCDvThoBToH6Uyhz1iLdVMEI/h7qVUJyIsKq0FebBpl2vZVg1sD2TSCzzfD3Di6Wbkx9SUlwdT
79TNYZSX3eT5lFYqOwpJVeNRygdfYJf5QtgMziwAaj8yyrmPZrCVzTAL1ryOv7I6EFGhra9nabqB
/PX1aSfZ8ZFDzBVzoSkkiHCukouYvID4gQMhO2aG1bdkL1brRZtn1qZA3z/AIV0x9MvGJ8+bKj3P
Hj/iFrTbfVr4ga1vy5QHxOP0zhAKVS5AFLHwheUhaJgIapscUUn3i1YiNUZXRE5Cq8+Dqe2KA6+L
ZzSyZ4DLSz8aFAJhQZjtoO8tilg4TLrQ0k3kTBYQtGZ5bMQZdTOIiPky91N70WC/beDyshIh6yey
qSIa14A5HYtvP3qjFJGbxrkd4SRPlPc5hZoRXL0y9l9kLa2wQIZY+/6jYJVJFl/ZTMdjhSM/jrkn
pM0ev3+u1u2AwzEk9RIyE6ND/N+DVJR4+3trCENl620ydB0q2C6+7cbYvH1LOISmSF2V+NE+aRcS
N81ZA5A1tYh4eeHrOzHFnCiOzDRG7d8liz47fIKVNc5nFd5i0DpIgC8bSZwg2zaGWdVc4rJiJP9+
PGySMeh6HTddmhHueoPKVr4+QR8VKjYcOaRhuQ27sBYAHoRtiTo30xJID+IpQRgvU2bDXDnwYvZp
2Y9RSt5JerPZ5+W+SW047T+WPLQEJXfHdfNOAA4GaW3IOleFg0G2zYgniWf3eMOPLIpXAq3QeRJo
kEctrL5cdkjdl0YghVlnbmbEMOFkMbD5FIXQIHVOjBe8u9/0xCRquuhgmt7oBlEbOesEUnALsZN1
sBMawLSSJQFn86eh/0kAo7ZMJMT6y3cosJis9QYE43MuUws0Bmt4TTeXfEhxYpH+YWK9fh+4/uMC
4PslIpBjRaVkIBTgR/4KRVjYJKzCdKFYIbR3vNeJGo3LhG4CG3hmMJtALU/BcDa5h8bOPL2yLO/3
B2TggJntnPMA0zrg2QIb/DSJy13eVmShAacPIAnvG64i9uDxRTw6i3AWREj3jBJXQxmNmnAVTVwq
VbB/kWdUDtwStdYjacjrQYYxH9EJGlI+v80sRMozOzfbR2yJ/hxhPY2bsBncXjJ8FvT9Ar51Nr5T
eovh09OnzMz8ySNKZsnJojhX6LOxMfGljnUngvzsLMGGj/pQkXY7C3fIltZcSTKxfHCBimGuZxco
QdaxEGtyy7QZLTNvI8RN10q71tjC4P2gWH9ow8BzSpBxKLeSVEZ0OlBIkTaXeRcCsN1AU1iC9RSK
/wSqxaGCMCFYVoZ49fG9VAw2QeviTl/uzUkaTuuYAXJH0Q2XIul0M1wBhIaU/WBoO86J7gvUG6pR
CJjqcLXfPw+C/jYgaQ43E9OuJClzkj0VwfFnC6gUKVYswn5WRVFyIlJca6LfHfQLfc4uTJVgZoJV
dXcYHe2xOUCEY7Hayec5/Bymanoo9ynBmXMG8fIcwdsKUB1Wx3ZKoZ8dvnO/JC2edfvH8xO5xGBY
c6+20ZDV1tcWzRbdp+VWs0o/AyHL7jNDdGowLs6q3zqCZBd+xhVRqE82kmljrjadgW+1obT7OXYC
8W11vDOMpEkABUHSX+NRNc/bt6E+xxgbmpKocNsG3QwXk8O/R7SQOokMenk8c12iFZkwgrl2XDe3
Z/QUVha4vMRMk/KtWNOD++5HQLAZCJ0ApPK+Olr67Djkf1Q7IO6kI7j64KBlwzCUnU0QcthpO2EO
F/VUIt/R80HUp8Jpq3ft49TJYMC9/xHMYJUsXpQBqo+378t5up5c13ZlIOUsKSbBF30Oaue2EeM8
m9aV8ivcdmNr0UyNzIhNWs2CXWS2wqy+cvTl84N35POkqNKyx8JjO6rWoBhBIDZqd8jX6jokUWIn
9vUrvXBamxOwcQJ5X6n5G77VLUqDEsKDSTDDz6IaQjdyfcAWV9eOZMWHon8Gpjxb0Bo3nXGpcfLA
+aGqJ3qdPcoBiYij8EOZhqvtzhtCG7buSjMt5JF5fSOzxG3vxSQznhELGu9Ehxl/rHYsC20oDrqC
K+IY2cbSM19RPonzFBxWDZA4R1vZs05rAucD0L9Hd9zYshtovQNXVr72XQrdEy8jfe6LACGEClGI
64ezZATcWAaxkl+rBzoXYj8RVoWhyvm8AvF0UuBONyKmBXxLe5g/tZd+D07EEK8MdF3Uzmj+6L71
u9Z+HXloFd4L095ax+OzL9zoWlfmUL66YCJcb52ruu0YuLFOedGH5f7c+QIeLX3sgb8LpxysS0m6
XlD3d+CeKPnJ8bX2I92Qt0KV4P2hWBfS8WW1O1xUrcQwvzUYIuqYBYYqYpPgZBHj6U1HBOOPVHMd
exMexgzawo6HI97qLrTmMvDdwrsKv2IDLjw2xBmxBdTDAOvteg+0wirHLzudFpoBh7UqvaPIe0gw
fwHzS2JcD4SSfdDeCuNSKbV2UxnPcGMneDn+6an11to7jOmdsH1Ga6ekFwWFGsoJkRRdJYS9PVlX
XakhoxyqRgbcTBl/EwxIcxTeESALLbrRz55lapQUetDaV+3tikyomDaZOqr2J40k/KkjqO3w8dda
Vu1mQ23L+ROfEQsH4eta5RFX8E/Drpk339qg6kSWcwKehN3NcB1kv3XIhnwq9sL0b6UbRZY4+sNr
V2QwcU4l9wS3SXxsIJvcOrunsfEi1i5/s5tbxIHKZKUJstfW1kZHuVws4aVHi6AgwqI1X4mS5ASl
F1sQYzwj7gxOLvskxN1HJsLyB38MS+j96tfI9rF+e4rEBVduMDZkP8hWQ7II+Hw40H2Lh1z/8Xtk
pPshbNYkGzb+ybzHiISdag3yTcoVmKUuLlcEaFQBJa/kZSVC6dboY8YU5VcWGMnyt9l4nxBCTeEA
9U2lAY/Xj/nFp5bAyI5KK7Dy5tb24SXwxfojzBc/ThniTyUxcLnITAZ4vDH0h+FwFRVzoHfVM57i
V5is70hcPFOZwJ7LqBP6l9siVYjd91u5+BEA/j3+/XXfTEMugGqlVT0kkMbNYdcMpGetJUwQTAJf
TM+LA7c7CvKOvWFDg/nyz3P1bNUPoTAPbt/aOuBgUUTQ8v6uS8/qypqo+Fdc4GJzcgJcmUBHqn8H
vvhWePU8YPfwxexe/+u6oPD/OtyaV0pzBej+oVKx2jeCpQVWuVY1OuJrNykTsRjMyL90224IWSmP
yRcGq50rO0kDKu0/Q2O9pTduqrh1S8K1ZZSTGMA1EPfeAssg5HrtWjpAfoT7yh1G2w4zytGoCWqf
PHcdEMDlZaapf3Le0oA6kKrs/Z24EEZUSzRQLQ0JMH1IyYBx/iompxLAxc6UEDfKN2kBHcMBok1I
+SxBe3+18fywO69VpZdbMHXXwXZnGTKYDSlIYlbGt8LOv8lJTK5qSHbiiNBOl3VJjdSUR22kj7Ek
qjk3iNhu1h8cuN6YBa8kLudXsOBc4hpKLDj/MkvIMOcoOfwjxBaKbyMOsePh5gIQi8h6w42/zn5c
vZ33Jk+JnnZk3SlcD6PG91QUiSYKjA2L5/Pk5aqJnhe8NBJohzET6AubSWosMHBzJsnwaGwS5oMH
B+5DXmyOX2MGtcID8uMsu2shj5iEQ5CSD1yyzv4JR4YRrUZGWxnOVIoh9Z64zZPM0hBV03mhQwta
TVj2nEMgS/29s6eE5kHX+oCthM1Awyws5h7AK98iTfvV/oMiDrOam9DsjVyMFuNDm+X9kkZfxaNk
LFFUzwtIqK3PbzCRmSebTj58o/UV4fCx8Hp2IAiNmPjkk6Md5LaqLwRLsTVVnGSYxdBAu/OiMnGE
bwjxJfr3Ts8GBOlCRraZ8xZ2cC4uZEty5d2mgsquAFvg36uuSKgPBr0kcdeXEbjwBjrPhLOYCmRP
CRoSN/Fvn1AnOnOlbWhMR+4/rH3OTj80VtM6RrFU+W+WvUraxWAaVZkcRK5vQ1/F9650Wsw4u+2m
CoD0fGjhUluHMiWPiHgbjaX4dq8t32r2PTWcOH2ISBaJ5IwGVY4ba8Dq3J6WXHyX8g1aZDpVdryQ
TM3wuFn+wimBzG0ZrTrxzR84AcmvBcIqzX3crcFZ/3IwUuF2LwoRib0SNXJtgh2+/RqIA52kwDaJ
NmAipUUBqMsrZcmow3U/8mXtk4mRwr+L1JBuUUzaIAJmR9kWtOH9EqrSTZuEUb3sOA7vIcljAWgm
b2/Yisq7+lb731r5PvKfnC8wmRABSAn36o1hk8Zmr8X2SD9VHcGg0KnfWAUB3QXjn5A1BLraoFKa
6YwqdwSaduAGSTgqKYnhhjCpcM255rv13M2XhjBhJgwG/7TDnLUiCqUlgf/Df9so2jfo92mfxLvU
Z4oRHhNC2qn3FvXpkZDeH2+DOhWIcy52VUw2FodkInEjxqKVAMh+z6uVkaPSF96tMF5DZtzeHBFi
MyJqVDdrVCguIK4ikqohHHR9lA6ECnTnv9d3JYqlsVVpCvZGPNtLIba/IUw4Nx5BtKhv/4LxmAYt
N0bmPBWDOSz+zS6kq4D97zoGxqAUNqN7ciB5FhiPPo42uFDK3FDx6kylS08wm7GaNA4/HYKUGLfp
QJqVza/ZM2JTVj7H1Zu8UaQnkxj4brtd2SARXinsYyjZpiAbVZ2WpstxTjhsyoc4fIXselKgnyd2
7j+dG4SfuaDuxPnESZEJ7jsezcsV1GS5GjZHVLLsiiqr4SUSBFitHcKh7j/u/wGlnuADYN/b8H1K
d9H/Yr0W0gpuUgtBugOmhTYasYHfBarVAR3b54WjspLav3sbsXgzGHOf5z60H7urT9N90G/6zD22
Igg3JsTYwZt5EGRowtFk0jnNCWLzlO6LivbRH7eNY5/dd9tabi4aC851c1J+w9FThYqyms/aY0xK
A/HLKh67Vt8aCdN9butMPoHqjMFF6UfmJ8v/dvhTp7HdcZHAQe2ucbs2vdTkSq5VuFcvGVKirkAV
pG5v32PaBW4A64kYLEIPm8MmdZnWelnG/eFqUxs7hQ+WvBRKVRnlH2FPg2ge21sGkRGbhBQcixpK
RcHSjHlke3GnJLRcp1rzB4PEDguAGFnkJpSg6L4trUhlL31D0Lzu3sWqTNTGSjhnLz3CMOiiplHc
2uQlE/9I8kdGRxOnepcjZpCLTwL6U7NeaEa/J7m95TXLynA0EGcof+H2xFbbbZYPIJLWVxrR0j3H
zsgKVa2JCGbGIZ47G4CJCERuTR8Fi5XJLwwMRxuXY1OgiTYERs9ShoqIx9sqAtSY9SOWuyoRRNoH
wkcHz4dUkdNu6dRRhgVI4rwQyes4U6+B+N6OyT05KgrdF6I6aWDDc8gOXOGFQgh5fv/aWptzfsUz
Cxrur04gT9u2iYQ9ReIOWeEucUVOncmxc8Xp3GaIEatcSlLBvL8/sfoEI0YEiAgQpHlidc30AgSw
am+b4csuS5+6+hyXbDHM9II/VGMjnTTWSaCsE976Bp8lG1r0rd3+34Mi0pL4iiEsz0FpyAK8qQ6R
YH9l+X4VYPV9nRg6iN9QlVEjjlgCuyuJuxo8MmlQqdEyOxizy6R5gnBog8j1BqpZvPeqJhbCKB0y
nXPKttQxU1pvbWQi8kUr1t+XXg2DFZmxknEXmkZQsKYTY4/4yuVg+k9fkkRvdcRtTLZ29Q9d+wcL
60txBkoAToK5+RcRYhVoHbNtzdsdlRpW4GTAdtagNTNK9xI0fkSMSqm0prpcVQfLDpGLQh7Q+20O
hoqBe61l4kh+kghv6UcH6y1RG7aTiDhpp9Qft9xyxurbdMiWprCQQY056w6REom3o901SWR6rpIs
I0ubPtSoUseeRw21sMkIT4VqzJuoEIoCeQrdMTPdPnYevZCQof6t1sKN0bEULmRBBr6o+5Pc3quy
xHepcq5f9F2YYZooddV5jZ78sj+8/a6W4UGXLbqgBjMyN2XYrDq47U1PR4kN9+uyGjRsQtW0w0vo
KPpl8672XI+H/nbm0CO/g6vSEztQuzWn1qbZ/z8Fu51EDHsz8fOZYsfWdlAmWMhJS/FVbGqzueAj
HlWkB15ZPHEOBa8Cxk9qILnDyJwaXHnab/lvHgYBbj3vl9UrQBBG2QVnTnpVtXCpOMOhFQX0HtCM
iNG4r9gu0WTxlWjh3fiJL2nUVwug66QHVQnZtAdd4XYQ6fhpIafiOkiU474WhUuP8sXaSZn9rSco
Yq6rNerinruHHRMNBzzz14R/Iimk/mmZT1OWkKb/gv0BUctlIYWNk2K3fQmCek7oZgSna9T7XPE0
FeBi8tL9Xolv5hEoUiiDGzGgdFN7blzPYLpuFnOaFPdyM0q9VbGffMXeUQWk46D6SPfuu8tX0PeE
3YAFs/3bihRhgwX/3ejEIXSP8YkclIapqbwIP+ygOMfU09XCJZDAOvDJ+qcGFlAzDk3vgd7x1roC
GRUhbdXDSDq9cZeRASiQ2tIvFxPxasp0gZMOx+P0JjIIbfCG+lSgw1lSw9PzmzKNOIlv8OVwGniV
heBObO9tozlQ6d+FPcf6GGC4E2EulUd5zQaA7CTc2iVbkJFIziK0+XjcKRPq7xW8i2I5m7O+P3sC
g3FvAsc8sft0l3kaxQX/N6HH01W/QkkVXZ1WMTJNDxe7dNE7d2VttOXSrX+FkiycOvT5yrFMhjpL
Fm9mM1+T0Hzj0eBFdWV+cgd+KOl7xwCph+UX3KtDRnOUD0u9d8Tcb7VN5EOtpen152t58pof1Lly
L1UvzxOgrZImSv+zoko0bA1pK6Q+n+6Sf+fhQPwyc8Z+11MARAEDEWNqYHkLSb5iRy7KZIO2GIWE
lw+Xm6Inb9omSd3a2U/xI6RFbzWpgxDPlypXIxhzPf+9aIfRuhUZvdfzDGKYUkc6ob7nIm6RluGl
R85f1T4RtykCUJmMY8uoKss6C3zFRl9VFRUzx2Od6GAwrBaPpaJ+JrYtnDZLPI5v4lYA1T5pAJaJ
wrPws1GydBsKaOxFqsbIvnlFmr9MbuMX0UCpN074pzmWg2wfwCp2q6I6YjzK+XM45HrzTOHGthz/
IkF9wiTB2aGBGkS4hi618xKmgKiqWPB3oRFaP7vtGew5cTaWefKj6vUrm58Jpmgp1c2sDJF6cbA4
uu6W5uf841C3LiTWSRoUNndmgU+TnhZP5gnT8nIdEaPkNt63D6qr0aupX6ssRBP2//WQenMGOLgc
Cim4NJDbqqTsP78aEt+9d+Oegqtrm2x+byrB2MgPJkNaGnkHYsB+T0EpjYpGa9whhU9Rij3Npc26
gr/lbfhn4mRotmnjAfJvEMLBB+QYq0s0cdQT0NIksF8eqiSTTMhx5d1W4R1B3LNF5B6nQO8QDOgE
75IGGoVrfttHZkKGPJWxvK8ESPxdZ8v38hbb7zBy0eEH3/PUB+JbhIA4YjsIXGj04wFQNZF3G9cp
fIGO7DjOcRmdTadm3a4o/AZ+pkaaAzxC/od70CQzn1aetrbDzshfBl9fIcuIIAb7HcNK+XUf+fAZ
RLxbmJKVRYXHbfTmNfrXqjiEk0h0AlFf+VKVOE2DEx/LWxeuzfZwhFNasLrqu44VHj4iLGjoLqyA
BfxbhqD3Iw6rpydiR2RwWOLLd4124n3roQxfy4w/ANh/W9IyDrvxh9SyQoSijBo3WzezSErZ+RjL
DlzlZk9oMKmi8llSaSYQagAqLQULggKf6KO+R8KDRmz+YlwgYANc8YTVY3qE+VfJlPjrt6dQeZV7
8waJeUppEe/8E7B2opWs+eXrKkqWPPPQcc+BaltihmLbGkwZG2k2WVFjCZAHQY0+2Pi6JBqCb0p3
D8dcURXLiGbTNm1AZyQBvIsw4vFFbR2XhIPZxLJpmN2L+cpC4ikj30BrVwYVzRpmiJHuDcaDhYRj
ejpKq8VmhyhsjKZDV9UJsxDIhhn3MmASCvtXVCD0a9/DHMD3gp0bOEY8jtBMDGZHLu7/ltB/Qc/w
Gn6Qr6IjeOwD9iHRhmrfLB9M1sSISjdcubKDQZL6hYimm/S0Yk5C6rNICo1JkC7pO5BEgOeBD5Hj
neq/P1Q26QdTd7iYW6+GcNlAPR6V0zL+SvWND7b0S8J5gLe4R9CpP+BmTSa/IsUX9sZdGWmsHbDO
8iYUJeUdU+ysiGv+Br1xBPp8Vup+Ba/BYil5YoTfrE528pq+qYxSAE7fdVwDia2KJTjUJ9/f9hmO
hTYQO+rH3IzJlTAUgXCLPHXS4GxepdkBQ3FTOQxBH9poqo4ix5/k8tWxteWlG0rtTe5CcrWBZgzU
D5a/XLj3y/Wjd3Djn9vhLDGTUegFnv5CgnKThQj1IknjufaCUqQliBm9S3ovmnU6Gxcsyw0na7f3
wfbEalQ1/f9XbHHOnrSbTg3g2rlQ83gBwxPhn1El/pXZhJAmmDN9j5qXTS5ocS/x30QuX6eEPB7H
16rPLklrSaivtzmSIpabrdT3Yvktu6Btm6nmG4JwwYOlkzaVlaR0/3B2Z8P+RaRJfvOVgDqS9P9C
mZY0XsmtTe5iRcanWNcK+4LCEwUi5tBVHdjOeXEryLaNdwjem1U3z/rU+7J88JyzS/5xPp1EDedo
Nd/3xa3mGj1tsVArurB13qhTA4w+pSWi0JcHiVPnAQnx3H0egvzNWG6TdhPKijUScqlVvG5Jo9FP
NyyLZgC8jDx9/VSa8VizXqRXax+dTQ2hwLRIzCEK0N/3/f84qMilaOdQxVqJkHJ2hNpfjG/jqm5g
K/hpf6tQhytZ2GZzgrKZLahgaaWOgHTVOriasbRCrYVPVDgTpE81i37C88s5olz3wOr2+ul3llMn
Jnaqki5Y/ynA66MyimwUvm3KTme1LhfOEUyxaDowu390WBuI7ZanK5MFGZUxkUqxdUj5qnYj/RrP
EQX0fQtOwv1b5v7b9baxwtK3aIpIU/sqJAb7GMCYf/6cS05Bm+oi1Gc4g+c8yyEnm0UflBv8iUYB
LUw2ioX4mfPFsl6XvKYVLvd/QAxp5/5uZUd5/4B1rhtp5ohIUu1OI5/7t872FR6UTrPf7SW5yNI1
403e+GraR+w/tKxKjzuiDjFH4MzH3ea/QI1vSd7wpMw4sZYMwdFNt/U7Mf4sIBApxjECtSN7JqjB
Xrlu9vf9JVlrIL9vPAEweATxlOm+gA6YcJ6CaswNrg++ISBDEqyto8xA9vP9YW3xgJKXQVulqUoh
adwuVCBbISwjKtgOykQhuIG64V66gZStUYE57kWlwd6PPorMpZVGTVwAkJpbYeEdM6TvDXO3y11j
1xfUU0gPNiAJ/yxsHOKXEo7WYf4b03ZIKYXmCKHr5kpqvrBU4FOD2NRE5NxHmecfACZylncwhL7/
hpWEkkRpP34ECsBl/y85HNWADLS2UNurIGh6zhwBnSQ7hGyEG72xKA9whtCC3nAp/VvujGCUJYAU
I/7+0Auwe6YSgwQXlI5WCop5jKTTN4lKf3j2Glw8i1Eoq7DfAtKF2uVEGFgukS1F+FzU0c90DDxy
StHu15FVx4Ra6l++fwd0QFGjIp3Qi+2pq+v5fPN7ffIxOtw6zSL+l7l9i4jobRsiNacRDycQx4bE
xgNZq2Li6P/BxjABxtY6mQcDTk1mA1XuOMaAGQiUSFKq7ewXlxT2QpO9koxUXe9GRHiC5TktI4oW
fiP5/HiJktkOEplLYGWtE/LsDnpDJqlRsricPQWJK+naLyJpCeStGniBho7/i/328SgdfdyTOCK9
7VEGxSsjOniQkTwj5t4gtOy3sUdePYjYv3GhNgRyCKBx7HZsJ7tWRkCklaQAbBou3WZZ12m3KsI/
C4i34w71X5Zt5lARtfuDKr0h73u+gkCJL6S/Wm9wd2cwUvYP+RSxMhRiNa8zY99qPxk6Iyy9lY5f
3O/8YmQ5UrzlEfEKVx3ZT1xYKIDVBPTEoLsn3LtPIX1M3qsvpdM3J0EVzY9HowzjNoTtYpapgyL1
D4sVbSQethA8Rp9pPnqVzIeROqBMg8Wd6TPWcbWXb/2zfXffoYdv52me9xQl4SPUWOyiDmb80a+O
oONzQKW6vFAaioYuFfCPSkAz+caMqcV+WPPXht2U5oaB0JTxh+39tr1ueW9uAp9pmzlSia/mn9Ls
YRR/ARXIiiyVifIRIKw196FlDPzMHTgTQUvKqDV1zMEHyGGSufW+tPdGUWnS/kPWkM1DWxk+K7HB
gDBFxqT7lSoRxvjdv2OKDoXsM05A3BMq2JXM++u01Jgip7bj5o8wroPXhv8163br5/V0Snli8yRH
5Hr2yUvZgY2MamfDTO2QKSBxeIyGyn/+4UkkRbYf448O2oi7Ix9Krdp/TiOQh5XcQ4UKQjgrjjNn
G5gsu/XoW5Qo0hcl1Nm9Ym5ViA4HyrAeAMJSbNpKlXnhisgGeQvKtP6N1CzNBf0viBrgE7qgOaSa
XXr2mPFVT4bTao8zUQUcmp83KB8wdTSMoqLqGc6NFCkCJMkuCB32lY3/0FNSbYQ0fmRVgUORFIEF
Uz3JABxHz+r5+cljt0QrRtYJF/axFUPfJJV7AXCtAN7HkBOdhKMA8mqUqV9FqMqtPlSIXXVD03F/
qGaMwwq26N/yJS0tQgcvq9+IxAqSk3rB+zECmoGkm9u31CdqxEpP+TmWVGY6v7dF48x7byYKp5J9
Rowq6RUzp0ZYpPxAgg1JRhU2SfwQxutw91D7TWG8kNbW2+CFoCviv88EnaR7PQl4bSRdmC0UVA2b
UD3H5BO6xNfPiYdL8I+N29eNCb+HwaTMJEN5QrbFabVZCJXWom9aLsR4fwj3mKcoCE7+D6P3GaUA
HYITc2xssIXMZKbjTJZhs6iMxbow1+At/wRZbFRrZ+EyGsvBwhuHwkD4arsISlopXypQ7jSWpUZf
zpid0t9cfuLf4WDVja6N4TFDf/OnMbo/SxvC6rndvHA3Fqv6zjTnl4N8bpTUI5vmbMtuSqeRVm8L
9wA6Pj9K6l3F1e8+ipPRQ8jRX0m7ORjCI8MSnNG5Z2+DPxEHvNUEz7nM4jaoJMtE4YzKtOH3kqjb
DO+DsMhpSDT7R8TA67xj5MzQOlrrNUcN40z8KDj+2bqCgUZHovZ21DZ4oqnzJGcuZSsG2ApU8zZx
jb9dwWtAp4vqOcJuUMGYxLYHPFkbOLzdvinj9EN4W3wAYDQr/Sj2Z+oPvYHpLFk3xz3TvD8pycWq
2FmrBsZ+IpXDSYlVtXFdm2HeJfMmQ4NxvA/mgP6rbpkNX/H/8ZrHCj2s9nkFXzWlO0TenG+pLZQD
kQEMgu65s1I3neoicp1RMv1QR5yBhfENZijizm9pXFC1oBTOSi/j4c7Qfev/mQ21ibkcHGplbJZy
HokfT9Ykyr38qVFZgdZokeNLgj5pyQnyiqgevwLUr4UPOcyGoCtsNI6SQXzili3aqaxphtd+1mAh
HL9RiBtC9xsr7nLSEE2SaquJWOhlIeCen45+76U83sKteqffvri8CgLyBlkYUpoVgGNobH0MbPEN
8LVP97CeyX8eDNbnkeZeUZeu38irpw5RIBAaSaOgHO+x2OpP4MEhOHdZ3iFG4PxhpTjuly5Ebz2d
wcEAFwihvBdc2pbq+DsYnnQFJOLCw17KED6HktzX9gBG+CR/bQy191LExDZqcOxSTjFkDhzMmN8R
JVxBJU6h1i9HBlDcWLLfIcjl7yGr8Gjnoiw35FuRX3Q50eYjR8WkxLIW7L4PFJH/y2ydlF4pTAgE
hQ6OiO73qMMw8wEzRmRut2e3LZkl4PuchgQ67JuAq+hQojj6bZmfE/UntIbtzgOncikLiCz/cn9b
r3f9q+8RoxIxhiBHvNprtc2uLIWb0N7N0T9Lwg1xzUJMKGu3flMEkhcNjZre8YShSY0r5xRTX+Vb
RWd5/NOKQ5BlE0XjCrULZrU2pRvihL6SSpU3cHRLDaIWNvEQ7jyGy5JSBAU4hFSabMK1oDdf8D89
uokYGNWgWwt9k4CC7r3RRUnruk/ZbD0GmhPf/fbWNtsIrXy7eMgvlcD+aaQ4s3Zu+tfUmmbHm9Gz
J+fSWqgM0oaM55s4UT/pbR+oPfz+iRa2pKVOxHY/e3iZ0DNtyw759G3F2QLZDfMbNmwTmLTbJBzn
qclGmjXdjtGcrs2stJok9jUWjMF4DtrSIO+hEAa6flwepo5cBLYFSC3famWT2wTHUX5l+eg/l3OF
+kGEjvKILr/qESrHbxh4Bq53VK+JuZhWPAmjhtb4ZcVLaN57BCPtWMENTWKs1L+kCuKQIlimqneD
tcPX5eW0H6LdkN+D2Gc1WCDxfF2z6FHq/FV2zV/x9s2BB+iVUrPVOKOS9RQvEyJWdxMEVd5+kUzy
flAMYnyCB/7mmWONG0KhkQKdgvsKVE9HSuiKZt/kLsLGTeQhq/NazFR2OQSmPF8OiD6JgbScn4Sm
A42+zvVUE+C7M+9z7P3Qvkxjq5/BbKWMy6CF3tbKtHWECoTAKAnk7MtVtuOmZCxVeqLhk0pvBUWX
mNm+cFslNlzBv8sMgOKe8DJBq05nn0IbYpxqbZuRecDetf31KYM9IJdp9uhgHRK58qrMxR7BjBdN
HlFDsUSEX+BwuSMSVHli+wK1ZlkAViHLci8/plgEhg1Q3NMD9ibig9VlCnUL+lltPEnYWaK0y7YA
yZNI7yCQVtd1Vhy9t6ISgEbn39k7yy5NOi3QYxvY6M8izCaitTTouwFhQrmm9RLP/om685Y5uKuU
rbwJuYVJVdToLWhZNLEgwxCZiGJhSR+NfNW/K0G9hku9cwiDGD2kIBJoh1airjTAub+62L6N6K69
Z3+DhPL0Qks8MvKJYifmeywiI68Upv7UcRDmQPEQjXZf0M/PT8z/N0AY5kH7y4OfaUIlV4klEe0B
ksRPyjm/5vSdawLZNnsw8+F0BvJ8LiknQf++PgMkns9RBB4d+6ox4FH8x4ZNOJ3i80mqNTNHWpg3
PEnOoEHsEROs95ZDSeGrghXBeveUT38VTDSSZc6xu6N8+6M846CZYt8pK5UOumOo05JdDmWRcXYH
kuYEX2w8AqEeMOghxIJRxSlvuaD3YXJREpA1v01ujRC/nSnWW/QptU+dAM5J2RHgk4gEyJqjdOPx
r2PgbVmsroQOazZWIPPwGgmuyxBDCJIg7gZ8g2vYysAR1FBMeOxlUc7eTWTBa9Hn3Uq+voGHO7u9
rIVROYyUI8A5Lt2nszlNY9HxTVHz2m+zyPjXPrcCKZRSP8kYMZiYTk0feKPfchFYeJ74LCauLrIS
CuuTNnfUyXIoQMhX9yMSFRux9wiOWP4AQab1DNgRGvfSIcwvsPOpjrs91FMNTKJUKSsBuw/z3jiP
d3Zyg4tzNGNII31NwSOUknRzXgkjoOcv7he4znp3yukhjbXQDs/4FiSDBVLz8rBk/+zPJLxx9Bt2
hLIvOYgMr/jz28sTuu4Tj21nbBeRFS/CI596DxY6vjreEjByupJQuGV0tGlDZHl2PzUBdrOG/cLi
0PwS8XJCoSiWszfcQ7amjmjnziadf2/rj6OCYEptgXq7xmWFBQHI5vOQbwj1CG99RVdGuD6PWVM7
jL8w4zSNGhOMgBCmAmMjQLkEb/+uGl2LauZG+kBB7lc0H2vXhdWQnZwnuxlT+Om7agKFuEutdFVg
LGA3SYS06Zu7iZf5+rLnbb53//f4oyHAdUbqN4AxFMLDp3OGpCLrC/bnyiTVqEuOBXKjI9cMvyI/
YL+t+Zms47AIW35l7L9fucfm0BfWXzDy18MHqTLi42jGyKs7GL59DLCCGX1xIRyEZ+vxxGabCzZN
ObLR4nEqPkDJ2clUhG6hFtWkwNAuvTEx/tAWolfeBG/GwIfxYOKxptJY6sa81QIXOZLdQ6CooSkv
eBj50PknBTRJFFpEA1Nno06gfeTa2Mpl9IsutoncBUg1xZ9Q0kU1JiVzsRtTdk0g55APL3p10o33
6ddVkAF2KOm51xHDb24eeB187Dc0iIqz8Ilp4lVVT9k7D4mQToS6LbBJ4Erpg4aOHqI9Ds6efETI
dwt5uGDfEt83F9QsgwKKTQjjHr6TF/hfNEGLkH5pGhI69lJvt0zPdlqrmGPr8c5nRnShLJ2mL5Jn
4iK21OweqHydXsFD+/4Lk78wpnYuNskug+IM418L8FhlO2eYgG8ag5a0dPvZlZ+OR6nHp30yhhqv
BDpekdf/VZQzPXYX81cBcSEhHSaq88sOIsKggM0rnuhltM1YkdtiMoeny75I8fdsdNo/VV71uTpP
eXfDYKHqbPDVWatUacIpTpDF/DJpLvEX8Fa2KOnHvGPU5Qm2GqZQzUlTkl1FDsqi1ZsuKnQLjQ5X
UNBeVdLZJ8xJCUlJ4tUavm6KCz8ESsinNzyjjGF6iMo0wIDxVnKcAEWuqW/9K3rpvSbJaS5VYwyL
/X0aPo44Q3LhtBBzhRkepfgGfg6lj6b/bI3H13/5t87KSp53kuiImL8rCVu563pQjjX9pzFkYfPv
gAumyAVCvxM5BWbTKB8nyBajUigK8qSO3XM5VuSLeqfpVED7kdiBtwuXvbqME/VfDB1BJj2vCyIF
Jevxg0556BDxg39ZdRHf37F4hmFKuRgdQ9jvAVL/TVd5T7tP422kY8p/wVncQwWNJkszTUq9gqub
/rbv+jB8FJqjTf/UTqw4Tz+i+xjF9uYO3tyL83dCBDTuP+xIbeshOmqNg1IP4aMboReMpv0JNexA
8U/Qie1X6OAV7Nz93Ct/xHLbbo+VnTSjLnKjBZk0qrfVehIua+h4DmkMJ+ToR1PFN1AKDDZMZJGe
qmfoL7x5w1FAlhnxCIE6SmRwcfgKWkUa72f9p1lYQ5CkW1IUKLf0/amKdy20zlSL+HiI7aMyqyTY
LUJebeBv1Z6AlMqQid1IIqA0VnzMxjmSH0WVIq14gMBBeawHyNGxINRwDJhj0e64A+sPn30Un+/e
FwtCrm5FSkWpn9wQSZcY2gCjpztThuD5V8bH7dTV1M+F7LP0nQZAlmcyZlXIVHU4mzoGNsjyJVnL
aY8hVdJTkzX2aHgdd+aOdO2WA6F92vBz6z9q8eLK6NB+OnULP5BXcAiiLyVHsjqZ0PNsuRusEi8q
9jQ91ZEOkhDt6zZcsWsTjpNZgF1i6sxxggWQNYR1tD8la6LqULDR6bVwd23qK/pzawB9dWjj4Abz
H/7FbcT7/BAvFKliEGi3hGUDNhajzme6w8/qgVQqSLRde0UVx4ngCPIkhtk8l3HdBjYwGqrE/in5
m8qCJAOSVo7c8OgtXnSTo94hBCrSg2ele62QW4hnuHTF1CnI0o6ZBWFwMlfp6SaO07S0QNw0QSDj
5dAokgLe9mNRoFSR5HmRvB3/gBZMKx3UvwDxSDvGXKlGdV7XemdSSG+hqKNgdN6oa7UVzoH1X2d8
yZn3z719VbTm/okH4dNeR1OiRuY2F+R0F2doyPaSAmMW3+QAy9biPndqMMSZ6u95LlhV8bSGlSeM
XNXZpTpJPG64MhxMbc9WYZdUD413KdyxkXXmiWOFL7XnHMSBRZ2JSRc/qX+wcNecCa+P8xY4m8x+
eAA1mVIdJcXB+fYQunHJMCI7y/lvqROj+ZhZ39u5MmmelsWxKh24jHcgsSxVbEU4SZdPoyxcS+aK
EuY1l8jDFwKgJLka+qbt9B8mcuEp/NkO6kZElR3TBhtk/UMQaT1offlZwIwhHZj1uFS3GrYvjp97
WOEMl5W1a40Mah00nALEJa/h0ECGUm81F+LmIP7FyvqeMR441PCfIJw4LAO1d/NCiZ0zKrlHEZ1b
iN8bZz9v6tr04VnveXNqRVzBEXKIQYxzUsKS5rdr3vkKE4gSr+/TYKmS0tZ/9h9Oze52AaWFGhsO
chhuk/eeWKbpF5LM720u1y+l8AbAJ1CapkTfvhydefNU+XWh0Fu/lhtBZESgxd1BL+Ai2GCVwcZK
DliouNc8oAzaV9Iwuoq1bceTJJwgVmo2JuQSSnncQfa63LeQYlMJ4WrA5mumnfc8F4jv9ZAY4A7Q
ViGdq2tNoraFxS7ogbqS+JVeU8LloPeJbSTT7t1TrpgfY7Yim/rvXpl+9ZXPVswMHMfIsvCUdAJ/
QrNGHJSdaNjib4Uv6Rtbx8v43wZzA0cyOxA1DqHcptoMpf7GZNR6fVqPD3vbJN5bTeK5fIdG34Sm
rqECG+wJ7Afr0N7EEYneMjeslovrYwetpYVlKtK2jaayCWPCOt/3PBc38ZzueAzIhqqgsfocLOWT
hhUQQBvt9pn8+ph+1LxdSL1YFG5EUvuAuJdAxOymOJhdt7bCMs2/ecGvTwgxfBUlyZ9fBTlPhgmB
vhIjLfpcN17nx2HwM131N1XOyiJOqOTkR32OAH78uhhupbABvt4fpCUJxw1hegFazcAATLkeXtcS
OvlKURl5EKuF41NMTn7J9E5KHh2yt81J8ht1lNWPKBRyWIy/EEqX7QeVrOW3xDgat5H132x6AUSU
RpFSwV+EYtlOV1Rp7ZKTh45mwzloRu85AOuuXbay6bK4LKWNiIlS4QUnyCMhr7ifkZJ7szvn/Pb2
iP2T/t6mGyJBbsM0ws8eGLHevdd2rC+acThh/QbEiOznw8nXrmwmnQQOQtxQ6ewzOJyWEMp9vAdd
WraZoJ/ECbSnmQ0IVRhBv3n0V6g6r/QNrg2OJ4yZRA3LRF8/aFFqjR1r6AEaO3sERHwprtwjPgkG
LnWI6DguqUZzS2FHLVcj6Vz0njfZ1qL9fVeZR1X7OeqJfY8RczSAu4Ge352gZUd9EPUbNkTcm0kg
0uW+uO9QwO28XKxGvi7oIxC5y8dZPpakjH9dfqf6OeWScyJVGg30su20O9zfdZOXBFSlwaMCNy7H
hkF6VB0UeoXTBUs6T8fpLAggYCa/2uCnkqzCzwx6YvLicdWwMb8mzRcl0RZrSFw8Casgw5ir2g+L
/zVDMkrmDYdsrCShwg3xgKBAlPz0XjLWeErMpptDa7QVxxoIqClneLV4CORtt1h4t1QYTfIuHeAl
m9pNZtR8EHdDM0RwPAuJDNhCOJmYF/4NZzP03SyJsqTan3msqqbS064IaQEN4Tyh+hCxKqC93+Sp
s9PfAGh7fFFCDoVtgJLd1FsElOnZQa+RBXiTuFwQgnjSwbI3uDWlMf+qYvIxHQWHyO/rxEc/vIPm
UiX6GyE656N/iwiVl+Of/zNuUpJWaOqfbB4maOei1jJg4JSqhRxHOQqZGoMfhudRerVrjArH8KA2
6X/gXtx25uAJXclFGqo/CWxfZlyZigxWbTfxvA3kq8vMRmNRQVGitv1Og1/d74L15MwboyGKPbNE
w9PVinYhgQeB1WcL4/r07Wa4byeUGEwJnKoPNGRqpbIiKNRnQ46MYBe28gETnglWdkwj2ZKw/AUN
nocCWc524uEaq9XvMJbIGaKIS4Pt0WDkK7iGa5R4nmoyydpDmjrnh+UPOjhGCzS7htQGP2NmDi/8
ZNhOjtZskOx/ItlyyW9Sncmg2+rmdlSP3aUTLxBzrf0kGJtgfEFsm1l08WmKu5z+ICmqFgBltEtT
IjFrXqqgxz/b2RQZHaBemi9cYJZUW6DzvvhaUEhBLLG7ekNWpSWlO0UGmXm+gcfr8TJ8vaOacWCX
u3fDva8QwzsbysRSKY08CbLVI+k+3pDzKRDVaLi4lu06FFs//gdGkLvF8nhBJfgA+Hf16T8tL00L
Df/d+2h/CyLK4Db/uAFrYxeOJpjj/yPehl4vjXkBjVa4nQsqohfONi1l6H+pjURVgZuDuJPk0E49
jEQ3WrBUzxN8uxzii8O1XLlcKH6qy2EZOttyFu6NekYjS5ZUJDtqoD1mkheJhKFrYEKIpynDdzoJ
Qaif/80oVKTG0/8DKZDtM6qiPNsl8htrN+zEmsiTFtvnzfPi7oOZI7zqP75yWX27CpptdsiQV3wO
Sk09kO+1e+PC8DB2gtiu5zV+IljxPpWP3idi4n0a4q80N0hMzMAnj4zbYRtEfhitr1RpmaKM1Py8
7YldoBiYgF8oQEwYDbiSwePSbHQQrb0lSZfbWKtQJmH0nInulFdWFJRsN5cSTO0wi5Qa5NxyjcBB
0JzAJWVHhPqB8rZaGYaD3m+si7e+hqOaOsEUGbmOFoYAYgzFTVYlJ+BeQjESeEKvQt5HZUPqPgyl
UyLCK7Wi1n/AhdmUHFvLlw0B0tc0gYSR2vOHqPUuYV09+U2ZUAnRZULPoWwEj2ak8rxYePVqkYZD
qhf+OK4YNhA+mHfJghgzssy+uiTkmhGahEcuZUiPqnQ9CAgjt+MehviYMHFCWDjzzxTzNPjvCBy2
/00syqfd9T3lzBtoSqWvud5uu25dI5ZHrXSgsP0vRIWkO+bX0Ac71258pkdTkV2FPSCLL2D2k1KN
OIm+uI1C8111ihxKDbT1SdvAC9yj0Iq7j/oCmu91XRbJVgDcv9t61U3sSmAR3CRaTxiLMgulU+T7
y8pLlh3d7kk4xE0TymFBmT4w5igJN/CVUhjHvSbKuEbw/FKqdOE0RvRIVptybumHAIwghhArKg84
2FOqNaiU5Db0e041OvAYpXEoQbx9FmHm8y/tanaxee+rxRvsjy96S8U57EHuDbvlYyLdr5XsgWhm
NGHNbEFfp+NgVe0GnLIuZotgQCxo/CKZQ608BTDnfkD84M5EHLSzuC6QXCxr39PBokPEGPH9HTah
Ji7aOgl7S9fCvpGiPSOIn1sx1oPtEJgVjSo9JmGrvniEryd7qIA/P8Aywn2aCVWIQ1n1i9XzwOGV
3Kr8Kz1LAmzLLU17kptQYlCn47dUdLw7B5Ndf6Mx4PvrZZOcY9Ka0KAhaSGiPJgNad6q/oUv1xJY
QeVOwzTZ6/GC1YRLYPU2GOrE1+g1Pc8vNBxc+xi9IDilQFNFXC/DTtBD8375BKKqlBequSMY/27u
/LXHGZi0xOTx1AgEe/xTUeFgKKIqFnWn90jm0H031rn6qOMX7FIhTPUOOnzuoD/YCBhSomCdvn9a
ITw43MrZwSGwRuI5ETFxJwk7IQ48RDPrufX314VTtihftCkEA4MzoeakjnUKfnKKdYmiZMIRlin7
RgBA+hU86zl6LNgmEo3fw9udVSpYMpjSeuG7WG/XAyxFEEm8bqS+myLjkzXK1yjmX1nRzcFIpOeV
eHXoxUoBR0HrvImewUtFz1jC4H6Ain3uvedON6Zb/AoXylvRyELn+5nPjhafOpR9J/+ElC4xzheb
cg7czd9kJ9P7KzrhLiUGA7kjiwtA6Ll660inXjMh1N430r+6jJeB+lbCdrpTKsOsAVNOHESrc+9P
eDAP/6C/a6aHzdAUmHyKn5hncHuYZ0dqaWiemOKR/pscfu6QjKVAYHNMor87Z76qFjtjgZCPiIJf
2xnp4UcRkCN+0juOKavx4x9Jssa5Syobw1SfiS2oXw19BquDq3qykXeVgUGazm/zHEUWm7HE+bbr
PwSlI9domZtCCpYK0xy7/QTICqQhgf032GkScdz6N1oukXQ2kk3hKCtSPFzFOrYGKdOPcnWFM8DG
2+DrnKNgWGkGmReMkaA1aA8w1Kixu7VF4S2ruqYV6gUy5hWr0giGdGuTLxzf8mxS8SOEkFRXUM2j
zGSk9CP7g1B0C29YHBvjjCbpNXibMRb7P2CDSIBb0UHqgA/gmvabwpeeilZCufnSQRoNS8sURqHh
KQT6xAB5vHI4XKLyztLWJk+CFCWrRRQV6VURiI/efPLwgecysamOYRkXHbZQGBRo6Yzi9nTB+pBD
0DhBcF0WZM0leFma0+WO8B8bhnwKep4EHeOb1zDYeI6qtjSAGG1YYpH1CSpeM2wBhq0FY+GD9oNn
RdiQgMgCzYq+zTRJ5lm4F1Bn3SAtX+fwIXcbZ1kD8NwrliLTzNoYfgIKme/ztwiVM0obEk3rSQiE
HEv1TNnF5QVvuAwTYcvIBF3Wp+KO2KzKK+qC9F6y3pALHvg64eadmR86+Q3lc8sMoaSN3gZA0hc7
ZnRkn4zpRRax6EepbEHey8prCb3G2CUxrJ6NyUmAq7BLtw7vVSRTOCUeStFMdu68R5hycgxz36x2
ryhaTF41Ek3TH7mkov+KzmpfdX3cwAcoutkNQSzNR7SfViExgVOhYZDGhyCe0kz9DUzhhEGTpru1
+jFxx/yKpohf6Ch70xYhGKcnyMBXOqIKyz0Ovfa4iCp1NM1uceYsuc5qjUiaMHp/bUQiaNnfG03k
JFdGMFkHphJkz5xXcrgfKoVeu9YsJ+LqsbDIMCtkStVzHrz9lEbySWe1JXhJtwig42dayTA8WLQm
u3Q5KbX0LIbZoC6M+PF763sPV9m0A9KxWEfxv/hHRrixOudDo1ntQTFyubeM1sqFxeYZVKbxIPgd
RwOxSbRYlLV6w1aMtU0yHcmDwSD0Cr4chGPtTSCGtUK6cbBD8P9RqQeOjPEiVNKy2726h6oxO0Jh
ZWPbP/dUjQtmNeDfI7yh9AY/QK8p/furHSISBmhZWeG6KqxtyEPX9xQN5LXgIxT+vFp/Wyit060f
mcgAlqQ3pXZuHV5ikbcytDfJpsDY8YWrfmVDaISR+HotKbBflgK7HcN8HPg82+kqSeJxJ5RjAIZm
RcpvwtYbjwj1F+PNdBK2gnkS1zt4kaaPEe7ETEagICdWSZfXKD30brhl/b5frqE/mz5pdARhdcqz
YQj3rgFUmb9ngjRWKI1gRbE7sPyqKCzIQIMMnIgRtdjjB8iCu55px6t4UvHyfriCKNdEa0y6KtCS
Z+tSaY3MI9U31LslV66kLyQATfqKToOvuNXukQUadGljodZtp9+GkwSmQlzTWT65ZXryZNgg2s1D
0CLMTTlbB0C/gDBvWfwkyf716KGhOvj1Ae38WLR4ByMxPNTMGaIrJvLXqJ8DNbPyFDu1Mj/c+RUe
XOZUkUOWrLYY1cgLyYG8eklxC38EvNEYMsSua7kngtUhIOAuL3/AQmo1y15AGcKz03X+cNyu/cc+
dGstIIjPyB8TEJ/kTxSMoXKwViRgIJYbzQXg1fgkh64b0M1Sm0h1GunJQue++CyArNUgeH/uS320
jEPdUD9Zh8hZYwPhR2hlGt0IJ6HFN5b5Zr37rKTCUAOdZ7fXE7afEEsVsKtul0aUZMnO6QIgBPKc
Pbgn6Wnm3I4IXLpIWXx2HoijtFfFDpYAxQ7LLipP2ghE7yZjuFITQU17mUtu9fP2o19CWrAD3omb
EbjVcwJLnbCBJbcXk/k0PzHr901ZDwN8BO5GfozSLk9z6iAI6ekgshbPCQ+r052ggW3J2sj99KVj
uA8L1V0HlLnRAKkHOVas2Wyfnzkp0gJIyT1+mi9DEiyQ93TobDHp9Vkz43iB6dUpYBty2lh9em5P
Py41CcsNuLORTFhLM0D/i75Eev24D6hvNiYaFmd4z/wdWwhKHZJIsgCL7xphdfJVrKx6OxVCVLDr
q/sxgyZjK5ojyr2AAhzvIT05xCrofLFrneQJdR4rP1C04XdisSPPkYvnt8HkKQQHDbNPLuEQ/gB7
qymUmrjm1XBXy5yJ2fSnPC7u33LrIOOly5Diupnl/H2F326slWeu+gKAaSoD+SeR+VJTLnbWzsvD
3H0wlRfdNcCSTZAZfwGEJEegffbo1pj3s4rNeTbkxHAZraQPYZ6k3CjsxgQBfVNbIUekF+qGCY1L
h+9KoElWEQ98adDSyzJ4Wy+2aLS+BwSGKn4jx4uR7e1ARnJZSjmIVm8volx1lMnFQrwvTLmka3Ly
s5T+HpYtE0Z9VmHdShWDEeg4mlK2V/yPGfvroXDut01Em0ytPGxl6ApL0tt13AO/lMfrJzCM3WzN
VrpmEHtRpQ99CnY+QC4oxSVWX3b2+XVpvOWgJD2OHJl4JL89+Z3OiPHhHg1USWt8WbVGMWERJOx3
aaC8lA+tT/EhmsISYy5q6e/WABAGMVt2uk8f7v52YD+wFP+g3D0wCe3H1hCHzfOAyEN3eI9iILmd
mfQOJEK7HgLFEYsGFqnRED8R5x8VRmFQ7MD3o1Cal/0oxR+0Cd8npHGBBZzqQfwDkRSnmEFbr+xc
1A178jVym6CKf+gy7Z8vllhEgDwNvvW7ov/VHWcwCCAvwEJUuG8M4kUcW+GcDpfPpGkc7PYl7kjw
4J2GPYYpXfNt2qhtrXVOYhghazI3W3FOsUDDswPri4H1+Q55/jhk6bAkEW3tSuY7261qEw2vH9JP
41qWnT6nlO32QEbiI2vYfNpn4TSwxlj/9DKQMyTv0Elk7Idv4SMaZQSndcn2mmm2wBBXZtcUUDBa
akXIHDkysvXN8qWdVjzMhN/3NHVlbg8syllF2VkiOx01hJW74ghLsuiwc18WwMEfa7XSDKSiZc6H
B0J85PphBnhrpXKX3/gjnCCIVs4R+HbteV/Y4av+0H5O+Gq7mklunEo8OhkQIkjFT4gC2UNQ+RGq
4R9TtApSU6gQquPXeSF2RaSlDsx3NH0S6YouMMWMJd/0dLwBQXiJlw237pZ9LNYa6dJ2oSmWnMB6
uMNClu3Cft8JJb1t4hlSyOMNRPowGZW2p/o91VEwUujnc2BkODVPmDR/FjDVTAvNUy72YTz6j/sf
aS9a7oaW0WSH6J4tIo6zLIA4FIZuDcq3HZpC4/m/wbgI8tlllvuZiFWvYBfsfEChqM4mlhO+UtXB
4QSBc/4Y9ZFyOL8diFqxxzEg0C6Jfk3fThn5xqpFt17megPqPDZH0Q5dFxB8KRW+FE7lZoNG9WQv
Yb6OxPI80Qqf7kiZJIx9UUS5O5NbJiYDWnnugc8EFTn4TgH6la6rpXvsWX6m9oX0wN5w92xOEknv
5tKQ5NA0waTQVclh2oxoGXmT/qaAX70BIn8NbtPGYIazC21oBr0Er+TEtoprgfhq4Wj+KBIV2E0R
HPG142IwgC6MSd/J0xmSN+q6K4ggD8i/WD0pJdAxsmYrnhsPmFrhf8h/JuhfG8C2Epk10d9809d4
ayZJ281aMIhP2y3AqpHlNU5snAjXmZdY3VRTkw99r857upAEkZwtVkAIjjKnM0gguEkRaWR59hc3
BBCpl4/apz6YNtI9SuvD2LGKBnu81/fxg4OUGsahTHDv+RLfi2T3OduJJn+gQk8s7ok+Q5GYkK4f
mBwJvWa/RpAD2q4DcZMWuOtyZBW7v3fnQqtHG+uW8R9ouuJ8MgdbpHmtq+k6GHs48BzGia3UVbR5
ZxYx/4izzV0AFQmWgsplhL3QDe0GOOtZKu5yzngxjO+ELkPLudKurP9EewDeqkzf28NJyw4afpe0
aydHHJS2nJPIzufGs0ZPIqkh+BpJMeFW8oostJbysC08F/G4WsUwO6oOhXot0POicagJHzmKy8PU
3OG81xs2kRI/r4JjYFhEpqTo0ACWH4ew3BfzMgx6MNuHGbQKWYL3SQ+amFeKm2l28HH6Zikp2L4F
CDjJv2v0nUKT59bA55oGeUp8Cd/vS6S7dFD4eFCbm4HqAbUNqkbx/cjxeGwD8w5ekisRySLvXg79
XJtu4v5U96Y45REDrSljeQUD0MyksSaGrDFjIDaZc/LHYSar5JYrrmkfCVcT7NCs8YoPQAuANV5t
OHAodlVIA4OruOYgsd3UsZx/NpMKl3WtC+enZOTQV52bO897+mjFFs6HnuX8tUjcnQvDBlhF14ri
e6n6MVxaGI/P+R2a/aQFGEZedUosfjAC8jnWBbCSumiByyZLkpIPAkVmUlPg2ozjNGIvmJyFNNlk
P7DTEcjPmwbekcA2EJEPvrOD0lamG6xB995+mL135Uh29QR1ivENIi9ltVyOHPpX1xiQWoNWkcIR
XTG0SLh3HGvvs7mTflTSkRYPmM3mgoUTTRUTkuSIyPVEWPisIOcTMTLKSe7B5/F90hABrI9GQ+MB
nHoSjs5SedouUkf5Tou3sc0PXLCAuTm8/iNx1alvmCUEx1Zl3O6CiJ12hk49wrVyUTVjcUrW7xEX
G0oQwXNmJowZ5gjPxcNusgB/ftOfciDsO137kZREpoAccaz22KLguwMBBaH1bPZ09GvEyEDLvaFQ
9M8ODtwW8yvNxxpTCc0e3tOzIxwkOAXqX0aGslckC9ZO3FqPzhniJhAnvh+YUK1N0j1SDJBAWMtO
nYtyduOscI0wbyzxEuQ/wne9s4/kJ+v3m9HpPOf48kPdz4NbHg/QwVqG6U/FAR/oBsHc3b/9Lsog
JPrCtCpH5NYcrvJC/qpF8ob8/wRZCKr57KxvO1PNE99rkdn1/FkftIDMGQMH9TxallaOPf2DFUaY
PWGtopejFg9c4ioKILQzycJept0gOX/dA7OP9QJHSPWeVmuGCMo5uf7ByxkZN40AWy9RabZmnZCc
XTh1c8rnB0FOWHrJWQEmZuN+Ol55r/rWoiU8wcvUXGQauR5wtY/+sgq0sdteR5z9591vR3BXG6Cs
MO0VpO9rl0GBd/YsmXDAuoHeWtAfHQWf5QBYC5i+ozTm45mzKjLYN7vf1EQH6PcACc/CUl924h3B
otKbB97joo4ak7lp7Kby52sWKIPWgTT/pS6NDwKKR/a1BYMVp8vhToyiOI7GWKMwsQDnsTQ+QAF3
uN5j3tf13eV1I7qaI/7sJvoyR09mz7QsE3AL3iI5QVXDCL0XBC8XrXDorJTzyINsPJcBSStirIDE
K/XTpjY4/Vu5ODgDulst6tSO5CoLzeMca6bvn0QEbOuR7SeqhcEUBtvs5kdy3m7InGu0YgsWeNK+
dd425/o20DngKRGxMW9RG19kTN+lMaCvtQGyW4XO0rREL5lQwiyjbS54Bw/NwXkpSE99wOo6Yam6
2BlW6dQKzP+s9O+AwxR95WJen0CmNxrGyTPh4i7G16lQiRc9c2edMvUekWOoQSu/zgH0e/Sjld1Y
jL1TL/pL1hb2vcD8qnpOk8lLFDY88Gy+8mRmtQVrzSWQr++JrAdiGnlc2qABdPZY8phrrzkTPBJs
RDQV5NExzP5dteJDQY3DVZG1gY5PBqhKNVZ4SJD40trfM714RynXDNlHSCPaaFjbvySmdCGCUtQb
H0rQdecYUffVNEIjX1jpYgf1lMtO/GdOOM0QmyC2yUKwmyY7W+mSJsXzoUMX7ibH9No6+drTHDUi
ABUK5ZGLOzSjLHMjU1RCP5r4oUvDSnoFuGV1L6a6r3LqBuatb5Sd26HWSafT/bl/2LLh/sgFBYHs
Z5Ds5ksJqsZyoL6spy/La4xts5+dOtJAWNXbH4piIBykxJzZiQl5TpQRA2QHpEdC010mUYfVgU89
N7SwptTw2Iqfw68H+2A7vv2+9sSxKNpj6BD2bWWLQXv0im67PV47YCV66f5mYG8uf6cnQdBkMS82
n1/xwKRAL7XP6BV5ZRbEmmz2y/KaCm5JaZ8SKqP6f7/6eCcPUPG9tF3TvDgcVfveVJq81ovP8GWT
SxskS1AQMk2FwINVaSgPR82JipW6BDiVFijNvl+lwnEOeIfQ3CnOk6MWjzHXJAd176c8Aaj3BzpI
vj2FoGVoIFVwEmDwyWUQ1Pgd5bb69xHS6/+mDLKAXXu6ya47TYalx3z88HHhmerMIvXpRwbO+IeQ
MGvi29KkHqpRaB36zItSN7AUAxbGB2lWfGM8ZD5ELQMYg+ME5n5f4rQJ8S/AbRh5qPQRHSX+2pWJ
kV+va8bmcnOdIoqpkAgzFT3f3kLZQljnzloGx9wIUWDAGVMnIbrLJCXG86Ym4nfW6KMk5cMVfNKV
ViuHE4z45ts+L4VvK+5SXI54GbJ5ij8nBLWR+ym0Z/mqx/41/pVYKaAA1pBPWZ0EMIA/3o4SRlUk
GwWkA4brps6INfu07kTRKNGTRQVLHA78CHwu7JdUTaBSwSfcILquMefAeJEa0V5MtJzwx+d5UqKe
ZQBqFEFtXR21gYwbHY5vgG6PCEdWtdhyrhm9jbDQTZICZlpwafAj7nW96+4xrvDGSKggjM3GIMBJ
N36GTqv4hOkdqR8W73I2gjdhqmWkIYzfb+EJOo84IDdcbwhK4XudZ6SbRffEUkxzCd5UgXtCuO2k
PxICouHtN/mimah9myoaIPrwB2j1lWPq4PnrlgzOwfRJ/4EHyCOB9onjN4GCZvnaxhBDbS42ZdqO
zr9DoN5iMrDjJaShckgP0zIh96FRWPVEusvBrypNIuJxsSjqMKOtqtHy7+8EuL1vE746R02K97Ca
tzJJf6LQR+moicCqit1+tBok8En4nmb1Nk4wLsgUQaFftKc5un+LGWpletbztdtv7ZwE9UdTwPIU
UGzgR1PMUQ8C1cx6CBQttodsenX64wBdNoKiXGlDbN1vK3/nyL9fsfUVgPZd6aCvsOrDrbRkzXgL
SokyK1SNSjvC9KSKdXGhMGmmojICKBpufoaPr6l4LB1jf+zG1tup3IJS4FxB6bmhIoJG/Oc94qgM
5buKl4sgsPKdrGLjFCYgxuCUFrai1ldBKTBtgCZUHimRIaE1cClRsJNp267NJFNlTR3a0UWNGisf
TW2p6lJ3b8TEAks8rimmIgjfQITB+EIzhdRrAxkhTOxxqDkoGoif7P4Q7kFMpRsol9o5h+38TSgp
sYybsBf0PEHUltWOGhIYtsTp7p6NP7QPlC2JS5dMevZ30GQ9+Joo4hUB9QjPun4UuCLZKzTo6Emw
1tcQ9pgbtZCl0mDYwqL7zrgfxJUr9aIHmYSat6Bq9Zr9PKPYRM8IJrM/6bHlZIAL8+92+zaRbwmL
waUtmIeH9j/Z5MQ8LbDCQAgxGG7Z1/ycM5QxDmWBRRvh38uxg5jsIX0T7M6Efx9zyl3D0gbyFuKp
rYIz11q66AHvskCTUC/m5dMpOjMe4PDcEfaMEKmG+q7SHN7x6wgRmNwus1mNsT3g+J76RxSL3Ahx
YPRHMfvmSN4MtlByNgtorA7sd/TR78c7zrKRkAxfn3byVS4ENoIu3CZfo4uewf3m9OUje+eeCdN+
6XjYv7NhLHj9LxjT5IbCmuO5YdCsVv6WnfzNZtQ9qvvrm568bKOsqMlhFX6O5CscBdiLK4ITYISw
EpdRshn3m2Gm4PB2ey/M0tPXxMTmbq4DW/Uhr4czD8xEe3oHg4pYLAt29+XGY0567hHp8pp99RAk
tkGyaytlPouThCOTbuDnaYrFpfg3VTqzkA+NEkruQuocuBccKEj+PfsV2om1lpFSjPFrJ+tlK/E4
xZ6aCVL2y8ygXdeAa8YLwSQlakiFxuShhy4L8LR2KBDfwMGXK8o5B9JldwPo+JGc9WsG6IkdyR64
Hlf0zwzXudMyiXrGbstBHVqGxykJKTExsU3wZJM4ARQDnmLYscRm34qOI4aNK9swQoqxrsW2eU2s
tOSaNz6CMSXdihYlERCEX28UmodJvIFPVRRIWHVz6x7UCOOcDP2HqHZW3ip6LwxoAtPfH+2DXgMM
28D0uxiFGBSrTjERQ6kSOEWbLCPfaOkmvcL3PEHqjU82nEm0dTDQqhTVUOjob+1o23NJywwMCMH7
9YvP6Pkyyu/rKee3Xk7yEpe1QY4qOwBa12RT9kVzFSeDoX1z6x/sVFQ+F0SyaNimlOsLb/hIrwdL
+jGuF34Zhk8gZcTRDyUzDY0fgKzni3X7oWCE+80ZN5uj6mZxkFmmgLoTOBE7PuZrJ8dMNEvv+P1r
50oDY559KG5DwJEVxul5LAcQxx3beS4EtyJzasLaixGOEf8SYBVaRGjhRxFCxolluO1QyXu7CEwO
1Wuz8ud0mLuTy56XiX6MQPOhk+fzpNrsC797FdQV4SPBPI40V3sDS38pBnYAEEPjQY7qQ9I8wqPh
KI/ZbK8M6rKxGi+L6B9eO474I+t0fLBc0pALvK3VSvGfG0edc1VUSiLWTvRcg6Z80HdhD6tLAd1T
04wwrDd3u2+vyjBSwqNhX9DIfra9EVwlH5Veo1gPodce1fvAgOi0wHjy6Pyl+G7bEG1UdrNINNz0
d/4yf70p9GmmpDuF4LvngTzLvPeE0Ra1c9RHLUr9KXgy/juGIiNoR7WPIgNT9x8RrUkvOVmmzgrX
YX7pWiYX5vjl7XIg8isSoB6ufbuXGmvQIXOtHRc2W0UR5BefaU0JOvd/3LGmpEhkhaarXAFs890o
c0wN/0vzSF8KAKRDAHBmqk3q6GJq+bsqDF02NYXgvlnQKk8C+5cYE9jEB4DBbbyu4M3tGQr1dFG5
FD5kkiS5yTBlFjV+JY0sQmze/Cv/NUvVDdthH+DsgGxSWI+JAudrrOWkwfQMAUwu4fWkhuTeiwyD
lHMx2qHZLqYb4xUm+kPBEbIdzaUpHCu+5dFfxBMhCdyH7PUhPJPil6pqdOPzHs6bFHYmK7oAf89b
j2FrbTN7KqFniz+LB9ggZOgId5kG59bhlc0l2nQbiuU00rb2yJCHvaeG/M+tu3uMHgW+8npwXJeD
vJzQ03to1cOY21Sqc30lCNILe7dNZkWXWz2mSTM7knFCTHlYysvLO0b0gUS2nbyl3M4bvwr2u+q6
mMWRbXLRDGGXID1YJ/rmrNNQi7f1G6MApJJ9mkLUShglbSRD0OEkkliidUqtawVPzu68NkN1JF9H
N5nTXstlrBx0hRFE3h1Wcg3C3bqSxdYpX0LIAmY4914wLuj4iwxp4Z55RpXbwdgFRf7nXEbH2iUN
xT/2XJrNFAsq0+lxA3OWOVaGtC3rmfMJM7OVl4mdVSnn638UEUdiAhc2u3MSfX2idy1KukTphaEY
wJ0g5kks4A88K/lGBXvbiOuO+r2OibSzK3bsoeqI2eM54gQFjb+LLfODY3r3/R8Gljh+LYSew+SJ
4JaO6XBvPmhxehNBU1RNWPBqE9rttLuFbWILiM9iwXzQ5NZmMPNI9RhKZji8DzAT586rjSZ4Yk3z
svj3DJ8h8v+IUDJKXqVVQAusEzcXpUvOh+JcHBQsl9/XUgHHHdbYhrGoxtZGVdeBctsIAgRvD8II
n3jyukw10Net3XcM9e0K06YgVlgw+bVlQJPCRJPxMHtHHYL8HzVA31uUmkAtnmI9ASF9ZIxc/MVL
mgP3sHYEHXBwAKkWzujqGQkqWe4e8BHNrnARTAxe99RofdukFkp4LuMC9Xv+ATUeHTbIrWw6SHxy
FYIgijp+Kx5lOranHRj0oYcFR1wh6e+mUJ6vsadM5JAm7aJotUgzz5QptGdP2qxvi3BXbbjA66kY
ip6sNtVLol2nWnC9k03IVOHNt4xpyEOMHshR6UVHvRtkoVd9Xe2cNtvjQnbGqFLuHPqrqjiOAmTA
zRaR4vse/q3ejZrJiumrLnmV8EKARYzqKBpBu5CH4kzkRfEJa7w4vKyikwbIDkeoS9OVSlG4B2cf
U8LxN18qcR0VF5Yln9nkrLyfzXL6eMdX2NqeW2EgnvpRiveR3TTkdCxa6UqnV4+l1OpXBdjSHqm3
vB2Frmnp5euanOJqWClHvYvzdb+hQviQKqXUA64DOQhUM2F6UxQdLx9Q7hPkjLTQUMgdmm3Qpzrq
OLmz8YLGefdorxVpFImXFIqRrDh+cUz226vo82pZXlcytsOhbBr+y6mXzCWfTm0kGxEuK2sFfoH3
6Ty7NRUeGTw4TQyCF+AmsaMKLDnotkCX0ampbwo3DOeu99ohqDl8TSaCphYgDfrLgio3lGLIb9Pj
HQDWz+5cb8z1RfE7rG8qRKtMnSlos7iVY+0bXaTL/SY4ridGxbpuk/Vi+Je82ec16Wb0DZr38xNV
3YyNx+Jwe3eTaEHBMs/b4K6cx5OZp27usIFdH1cQ27za9IJX4r36ZJ2P6UCeS/YUcXawy5qATVPL
JdjuMqTMWa2AGOUzFs7SShiLFu5qgFaRXNd5QZlkzVCfTazi0QWkGW+WAME1gVFCWAEX2KBs7K4E
3jZzS74OyIy7lO5jIKpOsxHAnKFb1zj5Ho5Vmc0Krt+tOeAO6bg5iYSCmjKaFnZVCZ6nBSnbVGzo
9jVZB/GblNu6BV0NE5ZDZ5adiXXq53U/tAe3JC8J5pKmCM/b8nYgCwxpbydpXI4t+sNS7KaEvmE9
yzAOiPnoOq4LRggqfZ+8YIesvt3YXNzKfAU2MvGMqNvKS5NNoGsPcVfpIlBHaC9IFjv9NpcNrBBR
bM6e5GaQ5UgfJqXwOvYDlAAPRhXHL/CX4UlP31NwZW26laMMj6IH78nFyG1ghd7b8+TlCNBpggqw
hUW04dS5uzqSRbKm+WEw0pmDQc87glJxzsSGI3zClobBXrZvx/1jf8/5CXr6TVIutR2YdZyUplby
kYmttSSGj0PVMN/pdQP5Rbna/NRFIF7wjkGXB2jTS1KWhMIn20HlyaVWbZJTDXemdDLwlebLxsgu
GDqrRZ8qB5IRFToldtGrWzyx8M4gg0y4pZvyNRrL+KZUSXzcM9rOUSqA5pzFP1NLiKkrSAXw2GMn
ycb9pG04NTRCNfH0nixU9I1EfVkSW97/70pxSL+XFU4EtuBIUy+Ym7c9bZURs5fa4J4XxAczqrq9
lVmAeA/dI5p+L6hLBZyEPrsldJsS+Qt452ClLvW5vbz3ISD7ZM5vAcFAHHEkxelUjX0vD6VSVKre
iSEgDZ20sUQT/4u0RBYUW5hTmqc5kwvc/VdAfVnTKfgKAoLos4su9P6ZLhwIwh3YPP0gKaXDhsMT
DL3ISctdr3MrLkNAJoH4N5YrtjTWVUShvqCyAvwtvVea0xiHm7Qzv+eCIsDdHvEJeBGDTYiqt2GJ
VNrydXilkHIhOGIsCaPGmF/LTzOn0R8ldIXZJNCtz0XOI0SxOU4gGPx4hPJAe1/JWDkIrn32f3u3
KrHk2cQLFUOJoddrn/LgHjCDUdzoRGHGDAU1hXTRf8nh05rX2ntxwwPvBg0RP9KVyL0Y/o5v2JAq
aZsNSiPK8PXvRvNmyEP7DrRIUKJpY4xa9WqrMH7/45YmdSNX3FAKxf+u8TSgx5hy3O83az+ebQOI
S4J0RfSVYHj+ABUnAxPo0sYC61OQO+uWxF4B0IsmwoQkPMG6xa4rSdJbH3lcA3l2nwEYhpO/14K3
a09qpri5REX9YnyLziwSIk1IFaDqK6qIKBLnES0KR52+MFOJkDRuC07PaZwL0E/jQ7CfdI/cnqd3
o37dHz9x9QXNMnu+SVSq3FrE6s4gz3U4zqyoA1VhUGswyIzmiH1admLO4HPHFn2JQ4WI1CVGHf+u
7tp75QCcrTJMKdB9oCD6dK8Gq2KgUIKklkUX5/PW4j82Xnzbelkt/NRSVE8iQI1JP1S5nF4RTnao
nKQ4RkQhSYhkKJMmuE3DbYN7Xx8cvQWzfkpvTjdztn8DVpYqjly8pqBfniD1bJ+H4c5hoOV9RhQh
EKSan7K6zlHE4a7bfLPKJMOQbX29XAIPGkW/Ipbr9v6eIc6Kly1gb+ABJYj6nYH9ZxLeBVEst0vr
gzfstktz1bWc6Y8uk9wz9QErEiiSqd27xRg8MlMZODOFoVpZ5/24QDq9U6ME41MsTan+1V9V9f22
wRiSiuAtit8EiK9lSxiVQcUz2/Rk6eWuWGF7+6uiawLUYKVG1duuC65KZ2ZWwhnB8BhKCeyD0MmQ
5IXnp2qkVaLYVLxecCLAez6KsSW1FmwYG/NWbdi9UXzRWp5JCH+pbhgka/FgHSbS3tK4IfFt8f3j
73evdrvOHtjvFk1R+blZFOSw67t87Pk8JQ6yaFzfsL0y1i0DtKx5LYcb0Od8yp92yS4JMm8v8Bjd
7UPIDFNfdW8qfjvR5jLOLeinw2dbp3OJ/6X7OrcwyhH0kJUWOFe4Y0uP0BbPfhKaio8MPIolHheq
+8WAM6KpYXJ7KnuDIqemWt5Djq8BvIwIzI3NM5/78o4JEhebJVcjeKv6P86IW0iy92l8N23IceYJ
TF2kIyafE4crOHrSsfj3JSpjRsCWV6dLI7bKMbGymQTNaQhaFLKAWitpgYZOf63+9F6rv9hv4D8c
t0Tb0Iku1m46TK1dimci0maECr8nFBEeedItMIHKMzx59Bs1Q413R6bhdhtAYQ7KKplm8F21HZRH
k61U7AnTkF8zX5hqs0dyJjH4u6eAGZufpPrjw7/9KJ7qIs4JiY9HGFb3UDUcr8+QURg1CW720iXD
fCmsF05KZ8NPAweQpk7yPd0bOHBM8lGxMB4p/ITeW9wQdgOaQmUyupXjD5CEtxdlg4+Z5mGkkoZN
x/UKtxotk+vHTndtfmWzb96OnoLOHx68PWYEpnDhm3gCB9t9OV5zXiOJAj+fRAZGBYK3HXw3D5OE
lpqpIWXNj7e4G5j8IebZIHxUE1uPBchBKPBTbJNjpEy+yQxCUKJku+G/ccoYsacBI3u7wb0oSdat
6qzIsDgNi65Pk7YAs3GibrkqZ84tOK62cT+e6zxRS/wi1VFlG5GCwvtwOBNe848F8ebBhVS+27R1
78c5/SN5DN1szUX+6lurZcApSHDOGhJzRWmA+RE74ZtmCvZdrgQgyDBeskP9J7z+1EPMAtS5aMg6
KEssXQQezEok7Xq38fcH0cFZyhj/L0bXw752/sLrYaQU8AHHmPqmKA2qcrNe0OJqcD4GQv5rh2TL
ZM72v8XuUiO6Ki32t3MsPcUGw06o7A7TCM65BT8r7p/bCjs4eWncsdB5o62CW1ClcC5Vf1p+AX/4
bye5OCO1saAM9p2qhZl165/1gsGv3889vaqVRV7tI+Fz6jfqZGbwEtYN/fECAjeBEOUTf5IUFtQJ
g0ewayhrqQZDKjNBoZI9i6JRbATSXei0daKkk6aiYdWdq/LrHvIV0+kiT3v5XOjAsA66MUuxIWsL
IoMuBmBoX12EFJ2lUxEqnmx6xhbnsx2y3BWzcw5LQko68Rl0iPIlbUkqG9QICbD2hxwNQjQo85O1
t1hPwTMoR1DDE93dik3gLdVabLQDriy5k8BXY/eRKmWts6AnzmSZP52tFyYYgiok5PMLxN/QFqFK
PcvljCDeO5Fo3w+ehfkJ5qgp+ayJTs5BjZ/uihUjx62sCYKG1/5Jx8Tprw/NEeMh444tTs/H/mco
caKaDjGx/KVuwEr25d7UbDMG7SD9LssABRiEBKg/q/+99zwhBLF8SuBtEuVX4yLfW5GPsxcqoLiq
7eNgrxYP0drjyVZqonOHNAZODBwNALKVF7eL8Nz8Bdp7T93Qex7zGovDbXMSmYPF+VpNBjMKO5jy
hxNvlkarUuxeOphtON7edC7BMsmP8whOYUdHUIJR8jrZA1aSaipjAm7f3gVC4cirVPMe4dRiUWSA
LOtfxhebm5zyHce0Efz7M2j0kmm2VAjbDKK89B8tVbWnrMMiVt29rgBKDoQBX/nkd1XDoHxo+RoO
tINnSBwwygcpOboAeIetaY9tHrijv34TEdDtmxWm10Kpu4kfASxhJSo7QU6HqG3w+htHHkhcz+L+
QduLl/ZbqJDFHBS0Q5unJpfAFmTUCDHnLuK7YUBaTBEc2VLvmSqEPz29mJrrZq8cHDzMS2eXHR7V
Tv4aaNb34AbbIP/BVpOa7ZcXmxTy8wzaUpfo9aVfqe7sl69bCBA7v4ijMx1cUJGEVFD6ux2w0AJ5
7r7CDTreUOv1zZIrxVPFSwignWsCdj0HyIzT+ooyF+WD5F6CNWCheTNQfUnUqbBmfO5s9g2QSY/I
mmWHjHYVv2HkF3WwNpCsb+stHdp3QiXGq/Y+cRyyyak9+K4OM0gilw2yD02iTdeaBm7DZaO21PsK
0NWSFagJkqWP/X7qC/IHUxGBRv3WTCoRisUcNdH2FHQkxhEKqq1MO2cRdOERzd91hZlF8LRjDvdY
dIesjiaCKMxdbbGvbUbk7imtYwy9GxlD+IAuOzK6bEh6d9wi8I+ixHlcMnKqLsBXqquF0+KXqlRh
en1zzta3sZZFpxYSiCRglxJYM4p3PFPo76z1dIQp+OcyyRH2zTA/c4aG2YacUY8B6JJXYJXIwzD2
wb1CZxvaIVpHg/h9N+C+H7UpIfdqZ1jiuG+uYlcVVVLquQqQB/e30ignoWZlQKy4ek71sJWoL2jm
BlIPzDvS/PI/oOt2unJuGDCiodQePyCKbTlNWb7NOxxhDhTGhP3CpRW5L+7DwnL6jpVDnhjshBOo
06pZz/8OM6RbJZ4jTDNKcsX+BPM3OcW3O4hi7G0Da73de3CYMy9gcFrQefL+aIc0WG7VAMcn28yd
dcZlGbGY8WbkBwdeexdE0UyRs8L7p/i0K+UGLcYXWAbWFmIlGb0CcXCNi8N3LdEIYs1bncylGiPj
PavHiG2EM/ugTbGg1ObM60t/em1L+c9y6xykCPB+fbYl+8SaKX7n5x63l4YFurnMkbVPWTwtGDuO
GXcFoT1yUcqf2l0pXlhJai8ysPEF/0PsXi/ignwbXd6JWDtHFVgNuyl00c6gimhrMmRLokQMFCAy
OLbooSe+XkhLm1KEUjBJd2Ylcbh/HS/6gH7fP2nVdLUJYLjddCNYi0uLhdVlHBiJqJjfcfEPprq0
Y7bdG7Dk+BPi7Lw5zDTwuwRm92sPJmi7a5GvWBQmQ0DM1WYTe617xdw/DCwjgGVjwUXJjyVGSmFi
6uPH7k+lJcxdLBlSiFOy5cgBn5kPZw4yVwGZ0HtDg9VtG30gUHH5KFNHo7PsDafvwTfG0KiT7ICe
6oNRKCxG+KoUIG7Zafb8JSYMtn2KvBfTlJmGeGwISIWPS9km0pwT26FgilfQtLcAcqhL4Z6cBQh5
LmbAG5qQVG2wwapRFTgElWulDjLx7hjYNrpAIImnkRIIutNUhu9DPp1EETSXVwepEdOcwwgfidpN
QSvcn6aLbIoK3R72bGkJ9NmWsQjFhnHQdUZvx547bu3vJFSIvxW4KiNG5Wldvg8rHF5JcFX875/a
dUKWwFx56tefUGu2QzgVubsembO876D0ST3eku5mfh7X71R1h7cbrpCIuyifwQeXL92cjeO4SbIN
SDswu8mBUp/2evIW2B4gtc2xZXULd7GX0RwmkNuTHP/zi5CRr+ucRPUvV5q/DVQ9TJNAP5sLzZKK
xN0qpbP/fOszNjhhuYxADP7kFNTxAIwaYDZ4O5sxZy9lo0jOBhjVG/LM4uHDXU9GsIqpnRDerowK
MMJrF72Nb/6Coqr74M/ny4L6XkRL4ZEJ6k5zPmmn5vnlqxbVHoSYw2FYM5+N6DguKt58QABRBphL
c/T9q2vBTwCCb85Y58ru935GzIqTyneR7zeDt+OGEhQA7/5oHLaAqqa8snhjuE2scSCZuMSgAhXf
/fDoVl0IuqYWZfrz35O3Vl5Sm7ZbkZyfpfQylHu8M+krL20l64C/f54KyiZfrH0EX/QPuHZ63yOq
Ekg8E5iHGL2SLTA/tNRA9PGabKsxldcGEB2FAVeCik7WBsbYS4asFR/mxPIY/Mg+pzKLMgTASbgl
82Kn/AdtKfYIzl0oyUbk60xACs69rvPJ2eLYHTL1a7AQQjK7gk8isXSUXNBqOWj+G8eEsFyYxyLZ
WrZJUAFkRiyLnvd04eP8zslrkrTIVWbK9Ey8WHkNqDy32Ye469ijhqnwrKFfvKyPQUL7GHKs4/Lw
rXV6cFD5N3Aoqarko6EJbpnzAON5B8zKnrXlFtrJIUS71fc0SLZ+Ikl3hJJ9g5/oAt31P+ZAfi+l
qFkkS8RESfY99YAMIgZV3SAie1vTgVMRz/2+azFAfecIkG4dDQPzS0aHLkWFbdr0pv9MJffX1JL1
nhsD5uk68P1Pq0ZKIYqj/6KheHgBY4dTNgDDUMs0MKQWpOKmIQ4LL4TAd7TMxMcO9LDi8eMTnMcY
Osnwve3EhFJtlS1o461SbdYfUSTtKuPTPilLmaQCYLkBE8FcVx7fZxi8Uz6hns0c1YF1m4/tC1bg
XjZ+xbWt/ApxNSU/M1Jhpgr2yYNoCaWVTtskwY6LTcjoY2EjJaLW/fBf0Ze6C61/kPZXpzUn64ii
EgVSrg+i6V6pMwdWqq5Jxk4UIlZrMLXOLbfx1AVEXhqAO5nR/d3VS56EIixzuRzCfBBqz6+DBxtF
tAKRzEtMKGkaIRXPMTYJJC0fFnPi2nw0PBLKp3/862MEx2C57YIMLuX7sOIKindUUnrnRAnUexKJ
g8TLAEAlbbzM1QRohToNqXUxau1aS1eKe+xfSnQon30Fa03zIBsM7SzbDqq9VFaLkkyVl99qQpWF
2n+4epx/QIPYa67N+TCLNxcEPY3jnweq0BB0a3vthUQwu3BPpBddbHV62gAullT2jvEIxk/3JqyO
YxjmKvzLI3au6YRa7S0BqbsezsLuFrV2uwfX4mgF8qCmpxObUdfutqF7HH9sZ0tzpqNQ6RYV8R2X
fajZI+05HY0iItHmye/RY4Rj0yOxeDmfKRaztn+XC3Qaddfw7sXIpaLzIJ/OTnwHUwYuJc9zHHAb
FxHi6BTKt0eHFcNH94d2ccHIC1oCZbX909yl7+fQSo+A1ijh3xxnkiBYQERmHV4qHEhnuwys9we/
8GDQZuECkGZYhmVIemB7UqXWZ9yJKrukwVGiuL4jS4i1K3eUp3oW7hN0XWnyXShU1ElR7mWjCwJm
4OUMZYRZy4KbUJwb+2DDiMWyp6zAJFTbhsKQImk8O/3L7ONnsrqiEeJeoku2pZgNVVaGBj39rMFE
d+uFYyrS/VuQ4P+PR4BKrUSeznvzQzimhcM5u+aRMM4Ext0iW/hQx7iX3CyeZXbqimQWkS+gmhG2
9B1EJ29qx8t2Z6c+up773p0MUTOywLXgniEZmOQKPl9Vm+zfylMuzJsTTxi6T7EfsJNtua3I8ubN
+Yw21HTaDMlWjUNKR4T885MVHMojZeu/NF5PexvP64+1wWV8Vp9wadJyAXsaOQ12MsUrDEblOz0b
PJeXZcjOTM2jmNjIpT/0Y8gzPgp5nLP/0yK2qJ3L8eXijAoIyOOsqF4wrnMfi9+c8qm7eN4fVa/6
VZ6lLe9zJm/kdSuXlKFU9XRYO5/hn4+y4F0um+ZxxK/N/x6O8V+O4WOxWM5lHnBSzJxLttBMfhzQ
gRt3rlea1kzQkbMrBIe9J60TlDHEW32OXbsclsQL6fqKOtWYoIxxhFq7S6ur/ftwEyp4F28VFD82
PBAhAlN2MJPmNzjz8Tki40zPWrjjdEhR2M2FFYH4t82V2phSaKFWjhHGLr+ERkZNTe26BIhVLk4U
VU6OCQWQp/nseqG5jOxgywvMK4WjGOxK1iSwGUIch1zNPs60o3CLCOxQ3ZRE2rQYq5nVrcl+Mnru
T3+bs99xAyWUG3LJCfhQmDk8cOlg5pgjrA30sUQ3d7YZGlNE/ARIzioBkkmBEk1WP68zJglwJv9/
GNB9y8Z0/CADQbdMm6KNTg9ibdRSHXmAuku0X6dQ9nrl4RWU4Nn9fxyXYMC8+Ph/g7vCfJa7u38A
cGI8HCvdgO3BpWZfPZQWmmiftUzku+B7dT4t+bI9BgeXWrHupa106udgOyKPYlmpd95pOttWC9TS
HYXARS2ioESzKe31eaCWi+/TWEeHTzoft0XEsCHf455wJxYtWUPvPT6Lc1x74AXiCCXpriA2896m
eUdjBkDgnvgzxrzLgrLdL/8sqD51xdQsUm82lDUqkRe2K+rIINyhrL1iWuLqb/FhgE62Jc24bbrC
Ie7imzM/2QtbednhxEAzyC4oYshBIxhWaPpsbHX2vXHQxSA5a7VpOk740AL1qnZCKux3CTzTGvyJ
6M+51qxuT1iJgH6P+sLK/LxJgqvhBNY+X7nz9ikTsFvsxpbwvdVf7vf65ZEJIGPHW1QRrGh3+c/4
qOUYl8Rh75X1bfVR8cmbmAqndgNpaVh2fqRDmMBVjGlQi5iqSb5XSru8YLdIu2S/xUM8ySk+RKuz
IU2j2Gr2QF32OaFkDXWkIUh3AvI06hx1lJr2BzjO3K0nqw4atLAt2+H0DqrOQdMgEcNzrcaeNlBR
TQKb5nA7/wj5EgVKPB/HB/0+t1IvpqpDdZg7q6LUAoJrtNvEIiFvI3Rqj7VMzjtudGCjQ0AlqUMo
xAUsSSGnE7L26cftT7nPHy/dgUSdlO8WE9APQ50Ke2T55SU9+Y3flPPdIaBFit0SGCLbiDFk3qlu
ILxu0eg7LQAVLWJigtP9BGK/Zix52LlU4Z7Q8bKltKRl/0gR6i+R5bBNkoExHVLJMjxh3PWrA22d
6MTpyWpFmGikslAUCjGbe5az4pNfkmkJTOQDw16irJi2zEMA6z9fi/0eCbAEUu4pkJmHRmpIKkqN
GUY7/J1eQ1hN6KX4SV+AttyQOYCBZVI5vgBQYtgq8jHQF1yyWbvsfwsMWK6ceR2pWACXa01ynS4q
g9MfP8auQwmTUGXuo0jJNtDkao6fW42NRzdGUIT8RiJskBxeSVPEHWtrPWrsEDhxjdoEGKS05pbE
gtHKWPumalfXMKZ1itXOLKz8XHwgVP/5DhMYtdGCC4bKLvLj87NYeCkQ2wc6lrkwp2hjavqQ87VI
AgEnRxj9rfcQhwkTlqhCFOFX+xPBuFMp387sqGZ+4TIcKMKaivcqbcRVkCd7SzK358r6PedAa1xz
Qn+RXz84jEyrENt/d6ISxrTyi9+9qZLslm61taiH5RNu3Z4wQmskVb1Ua993NjUIzbI4VH3DQLna
5qM0hgPmMJ1aDK0gc6dloBloHGQa+yzAvDvxD9ANmSgf1nqRLalN3mvHdFA88EX7mV7hsdYeTQlu
4XoLpPLvGXVTxw6e/x9red+pdxKryCAwSqr3PULTU6mukk8VAzqnj8v0bEeFLoIeWqMG/aejVcDP
mAtqQTJVLGNgop4sEaRzIREcpYZdtAUIJWIfTB7qDtgP0y9e4FQ2L3136hqy9N+sSlRKpqqSQ5ik
wn/qhb38mXjBqbkVAok5BaeE6Qbl3pFDNiSWdKxd/DC8AyduNp03qOdDgKvdUQlD+seYZtnqOqlj
2N1US7jqMN+CfhCmXeuFVePRQbLnay9AjyD6A8KgjKaVaWmoma0s9qP14YvhxeC18awo3lTqBQDC
J3BnDNz3AmY9xLpNfXrytfsgCMZji6hQ1+Iw6ki6/ZLyPNa6uF+uh1IamuhfkvNIrLCg09MgU8X7
lOFTl69janymw9e5zrfi6516SSLZfcMuBcNctMaRcnrZl0PsAPXs/WYdyROVFFjDQECnANsYEtmb
YYrHRi/6gb+zbBDyXTtNPkMzwlRC9+LyCpCyRNbMEOyu/H9iOVCIaRsQcNaoisAxg3OhiTHBLwyb
0ukp2jAyNdFtNZAQ1dXRl5FJqBj2UfTLS1f70+y8H/ENPz9BLiOGj3ShTk2YJq/4NqPgcg7HNSSO
4KNix32Yf+HolgDqcg4oO12BmlW1+i5Pl161G0oAC2/OU/7M78nYsiHe/XrfJzZji8nG8q2bjSQW
aZ6W4CTkmxc7XcGVtIHLI2DZ7czmaHYkIKbhvXk/pQQqnpK8IjrKF4ZlQZCc5dBNPmRpW2H+iWAC
yjk4QBBSeoJmxCIr7lrLX8PyxKlQEWIvrayqRieL1ZZRtYh3rBrg+//9fvLn4dA91C2dfH3IrPVs
jnEvsZ5vDh9ztFr3OBPG4jepF1YhfrHAnX7AdV5Vbp9q5E7wlWrtfBBox0ulU+24dOrEOjIaIGu8
B9PDxiw4+p+bhlOpwvtVsIyvj7p+NL/oYKgbDiXYkR6gNPvNFPQ3+Hw3Xq8uAnLzwQImOJuYNUHf
uBvViau2sDIYSQnbnLJD5y1QUqyMUralUmUw/X1mMINL88hjyhfyBwka2jtPUfYIrNL/ZB9O+XrH
Ueg3WuIAYZjquSB0Gwd9evyp78dFOk3IHDa+BRyfbnhP08JQv3gDET8Qf05/KGtgSGlmX1FCz/KY
DYqUG6bSalAp+c+oOZWHMRjKYabDERM7NpxZzwBDSBFFVx1ETeblTu0xItga8Vk0kS4VMA/4Qkam
xF4LY0tEC5x0meZ5kGySo5OCczf+HhOeS9+WpVIuexVGmMZmALWOGRQvQXmiRltzJJAZLtt2m+dQ
s7fCCawfeNrIjId3vtjwq3B0X4ZMFLBwZlxLYKlDAd9Tor/F7HWXmkbIAtSIc50TgoLX6dWW1Aka
PsUhK00WNIZgjStYexG31g067l33PjNKGM5R7kTZ2O43Aeg8g767l/yaqD0C8gIrr7qcr3sHSac/
pbLYyPwRMSXX4Exc84noc7QH7FENeHwdZ3cEIpHSWtANrVo4es5nec2Gzp3bjU4oZDZbJR3Nlh4k
08JUANC6HgyNlPy+QLJ4yYBJgDNoDeMS2Bo5k1DYcBNnbvh+3rHT+Vf1Q+qGbfObJbtyoo9XL7EY
WXT3hUUPQvfn9noMADpB8ktSyjDV4bCk4N2728LlSEkP5CsESfG0IvOpmJ1XvEB1qALay6+4sIZ4
kn7n9vMzSDHh0akmAqToMsiotN0tIQScCSLCbKkN8ghIVaHKNL11LIeTzhwW+12aGzJ/ecJYBD9T
cd90NMsF2uKj5M75RiAqlg6j4KpVPpy5b7t/62J25hsn0W+4oZkrvgaF1mmJCOV8HEGkZle4QsYa
r5Db5nPhwlpFS6zedgdu1iJVfP8ZQZd+GmqPYczq9Lh9Vsa59RhjdbU3hT8VhEtx7UO/OTO4J/x0
hgBpeZ2djwY8pn1AZY6IQ4pyrN97y6up7xdrD/xaCORvgioBpvAQwFgB21eFgYGJygdF/Z5MS0UG
8jY4IMbMxZf3InNtHFcr1JQdnyzAZgeboQF7rGjUUZi3XCwPxJ6UwoRQk5D+6fqUrQyIp2/F5YV/
ZEAxAckDeWsZYKergnC9SlkUSL/7f4f0b/w6DahLugdgKtg0jjyZJtucxlycnXxhVircNvMvSbIm
MIbqM5dHYaH1EhhfRqsxp6CO6vW/HTLVUUGMc/XkRAUOXf0V8mLa+4hj+2kv2vykD+Xgg2RyHYL9
ShWuylUqI/xsRVqmFNnCdab0cN7J4U5kEdK9Yqi4cciaP+eTRXSYX/zliFwKCaNmICxEHnJtirrJ
pOAGmDIJ6FQeZiK9RgkPD7M8R5lf3qwMyYGgX5BsPw8RQ8feSjnwWhnMpeyQE1tLUTzLkzvEokBj
5dICfoTOveHGkR2oy9eCBlj4eduqUX4j6aFJ8TIqon1MnRVSc+uZm9FpA7VyWUoQzaIEauvJVFzJ
gOytC/HCa193u91UzGBkfIIMUAe4o9UXoahQ/wYWOC65XLIgUaJmt1QvJLclhXN1BK8BxukUfGMy
MqSJZEO8XkpkcFViyOmi6xVaYyAxr+Iz6cBZ/bJYJUfXCwj7SGwCfgrtQOov3rbG2yitXnyMflI/
cEB9PDNsaC/bTCZraQVlFYvubHUpQ5pm4yvo7yfibnwy8dJJqYMDE+n8TFos01p0esxjv/gp5Hy+
jhUf0LM2eOJl090jhYb+AvPkNIlm4H6vNK4mZzjtILAw8GaYI6sW83Z35hXkFP8wUmS6ZE+I2BbT
Tc0koOVPNKBl0cjFnTYVXB/w+72hX5gbwytz8J8oKoumyRTlwvs1f/8DYl9cuIyPzlXxD5t+GpaP
DrXeslSb8mp0gRgSM0qQMP9us2g52iUpwQ8QXFtZ1+7mDDY+OzwUqVEHsFcu6rCy0YCfj9CPo+Oo
3Ix+tE30rblFAAaxMHMFjq71IZjxRLIh1h9Sq36f/7lVaklfLQzTUda+zz5FEIGMIl0cRCjaG28w
w6izhbhC2OA3FL9MDfIxQEbrCJhEq9jphE6mJwFuulKPfQWUsMysosZSVeS/KcSidq85vUiQNXzb
WeyqQbbV7dcj3ZsefJ4kJCDItSGZxAo0iOhWNfcJkWugKLKGojtJR6aqC9g0P2eyHtyAtjcUwisa
f+jLIuNldFXofv7JUNixTwXG/xR2LMLmzJNxPudr6RcoZlHNH63JToIUu9Pw0iV1ivC3eDU1VgTx
85jjazND/eAfaH8OonEhm5MbUfsJOLJC5gsseOdGqiq3k5fqRS0tC0tA4t2x7dgBzt098qqZg9m9
ivShIFuSHUjC6SRF2vy6TCVoW/3qqfVm3OqMKqO+3ROx/40F+fcni55mmGMMKpPtjirYU2kWO3yK
IGmv/1m31/Ul48tSbrI+VxZ8PU2/AwKb+TSYYJtr6SYlTXQcA3l10Qm5A60kJyennsMw6gMOH4bz
MCj37xLzlJgdnyVuBw147MYQo8rbfBP1gmSg2sPOvxNpfAtyHwAgY4uy34rSdiqitZ5UeSh+HcqU
yn4SMuNFjdb6jO3cZM/bLvErz46WpWS9Nyowp8nl9AG7VUNnmGEXDzV1rtR4tGTJjGT3v3HYx6BQ
3ti/7SV2eb/3QoNzfvNt6Q5oAtAtjbOMOjoCTDTvZzXQ59uf+a7vX6Yg3bPP6B181HUpwlw/aMEu
SA79UfCXT/BetbYel4F33ZG+t0XPdtKiKTNuQ4XV57dczdgyYUcgDKFa+bvutzTQ8to+uUXLVezS
ILv+YcxUs7TaChYU/Uafe5bD3coceW+5bERpjjl+4aUTHIFeLjjvlj0WL3MLOCcZ085D9mEmMrL5
m12F7YaeMqic+IMJ/xsNhv4+5pgNz8Xl247fca35rGlzjE5sETy/mXhLJfpLncwl/2oJ9vbOw/6c
l3IlKfQjyAh4UuBlQ4q46+rywBneA/3eXLN0mBGhV/7eH8tj+8nYXagQzSoED5g2BzmhkEc0sSzn
B8k8O0rZ8ONjZUzl40+juFltEoy/7nraON7UuTs0FwDCQqo5/Pow9OZEEWEbDxMkMvFsdzg6KWII
PUFGL3Jm2ekbPOpz5/atfgeyIBYL5JckbmwOMFcAabbdfiWTpM6OeECKAdbnz4IqE4ZMNtOlSzST
7ufRZGFN6lxMBFj5h00cTGG3pqPdLyZf6Tau0liyxXFssP6rrvTF30LjlO9j6x6GfJCZb7uKmrLc
rhehEm8o0OHlNYutXLiuIsiwP/ehrPMZNmCEvhoTwMwta8AH9c+KsvKHHDhQbU2TLaatYrsnsAJ+
eczMgovYbcPFiScBJDJPayHq3LTFTr2PtXrXLNfA9pXsYJf05cx34oC2uTtDu/mvjUR2lUw81aRp
HrcApi8eSTWew88UJbcaIkiRdSZUqrdryYEcjQ1f0iDXRO8Jy/S5OSlJWIjwB1GiDH46gt9G4RzX
AJAFsWS0kyU2Z2R4ivqnwPBSKz4icXPtbW1PsVxqCRnVTaDk+ragLZnb8zA5nGGHmSRZ+d3Bcn2c
wtbcQWU0LWe++REz9b5jjBFf1+5Arz7Hg7nGmQzcFSksoGIOFu6Gr+SijmRPieAcywhT2Jtla3T5
nsmbVpOFgfopg3GBPaB72ax41fA1nEKQZckPljWeqIfK5bMIHlQrH1rIYIJk88/+Z3n/bt/zeP1E
2zVZmCyPVXoM7ss+9qNlXCYKn2Rwe07+yUTrs54CaLFc0i52NIGBGq9/AIqMl/Rot2BpOoD213np
1uv2bVgeD5NSDypdCYmPejSlsDhFbP5dQ05hkHmI2e4HpOALMXW7lGzmh6fPsUuDtd4gq0iBtC74
/np6zrHYs9rjOUPVuQlzIrzkK2zc2CwStUTHqPvm/kG2ui5qBWjxou8/v6mC+Gp0gBWFOyfHNQMI
9xKn35IP0zF2SAez81K7mxtuNX1G+JuD2vCxWigQ2E12zob0voLvOxl/8IqnXvR9IX7z0raL8OFj
RrMfKz47PEwfMH5o8Ch2vMPxVzbAGDHifEaeKoKpLcdVH67vQU0Q/7AZSClUVhS5bMCoFnI9w/lK
ViUduo6511zuSDc4+63ccid05SOB12th9PIbneSpe3T9c6z8+c5Fnt/aaDWRinaDHr1ZKu/0qq+b
kiBE4DLpU788/PzCp8rsNyNX3Opb60iTp6t9tRfrlpsAnvLNJ0gl647OeADC2yoxh8OMEnE9zVHl
dGIyCmg3m+/aJM321k+Pssv/NQgQ1yuLKDQghAkCOpXxvO+NUUkZZyTancqohRGvRh/32ksTTr1k
MHMc0yTKB9ZsslMlX6X8+BpzMu3FvS4e61/8M7isw3Jy1AKh6k/8hb/YLM5fETJPQzgTh05yOcIC
MVeSSjuveAAVEWYAfSE8Oocs+Z7n+UVVnnZKIlcrmyCVOFz3+kyVE5dT2g6QGvRnr353lqomrTe0
wLyjOYYK4Sq+qmkxtzWEv4a4zMAaewGkN9DMEYF9lrEUIotj/p9JyZDumRd0xc4xQyLmT8VL8XdE
cnxY87g2laP9F85k4xq4YrzRogC+O5UN5r6qWBh6fF5bQOAHdwvwTkOlA0kma3hoSXVd71SArIQK
aUKxoKpXPfP3mIla/CE2d3DBeFu5LX+zediOIfiuNqQoxCIuHl2DaEIrrpXdZ9uL3CX6uDaglFza
CSzV0of/UqQ0UuGu+KQ6HmmPKsZ3V+TuFKTXdFlHzdymC+th+XbrvEGhR3P43/mI9CfNaRfxnmG9
KzwqFtF6ig/GJEhkgWaD6TLOqSfSHWOL/54FJaDzAW+nTyaypO+JTMX+cmA9ckwt9Kyq4UDknlD6
cSxSTFRxppgUKzrRJwlBkukHWul7jjBXIljUZuKiKXLLqGp2bPa0t9ypkhdzK1hYHAQAtHK2HSbw
OJZCrUsJipvZYY5ypb1Ak1D1crl5fO0l3WYlpVZHgWpgZnZStV9r9FQCX9G7x18Usu4mVL1WUaeW
8NsgzHJp8l2drr5fIjAs3d4lb5eg7BOZaBJQmbVmUbwtA4hS771OmrQ5Gj5r3Hf4PIdt1QI+HGUw
5lDX9zbzhbqSBf5za7PWfeb53GYvtwJkzT1zKFMKW2W1TER0p1a+4XhZMpsu3LfFlKHht/ZYmEvI
6ugnrbUbvvfzQ2I0/IBmQEywV7wwW+08VmC5h0qI4Cdp12D1odAguOlS6S/qiq3uwoWtmoGGH5Wt
4i5oTLDgzl3G00IMgMh/E542iXgLqRmHlMS91YJT/ADJvRII40aJis1xUjk+qX+1dpHifEZ1QQ5D
Zd97hZqL7Cgd2qQrg2YSm7ZH0nu6Ti0fKoPqgAiv9bOFcJl6NIMXvbFIptxUGaG/fyMWHqgVImIb
qx/vEbGxsdYnbsgXGprW08f9SxwctxOLMguylgCNV4/UupTQ/RQEEhv1u+lrFK8v1J4WywyC57Qg
MC87Au5RgDtHoOlqu2hxgsdQGobfZdeM+/ksXYtc18l/gDl2CCypWUl3vsF7TUfo0J1dfNFm30GS
w2kP3/3fY/Sr/P20Gq4eFaOwE/WjdpWHgHA6hJWhFNJy310PYqMUOLbNR6hFLqy+OPulNouuar8B
N4XOERRU45UsJ8OOrCul5pCEiocvnxoRocUzpPdXlKeCP/CJkrzoTmoHOXGZ3xauq2AtEHZ96lmF
m8ExTy+Znxbk/Wen08ceAN/LP0/3PzDigzilssNvCPRIzbxl9vLuNgv41lNw9vsN2mTtVsBxyGlE
XTx7Fmiy+IYEZch075MM16ShVWnEZpVh6mxSrl7lys0TEEAMcPzIUcC8ikOOJabKIuXGmd2jY6+m
Ce2SHkcvbTQ8c1i9RrPnrnmxMp3zvgYqFi5Vx+czo+LLG2tt+US6pXGGIkWNomtJsrJ6dz4oY8Gd
vQJoShAT0T/vgo122UG1ULCXQpQkLX4wBD0vsCdcRG5cpiKiJL3zyy4Zrmsfxjwf/K4nmAOox8zH
Y087m30L6q+vHnLJsOaRjUxyr/tvqXB/9pKb4UIA7gcOPzVli1Uu/mFnMUMDapBWtOLnLparby/D
iIkN4IGetGOsDmBwE6WmlcJH9pBko2LbtMlnBqoUmhAXSwBOHMNo8nOvy4f5yc8VfZhwYf7uAkKd
iqJXz60JRdPEFxa/GUJfSu1dlbFwy7jEb1eNZA8DZ688jWFk3f7L1505GfVbSTgHaNB6QvucD/Sl
6gpBgrOGjfbDApOhOPD2xL8BMJlTbg8uz/Ft/Lhga+QlsCBMq1tt8S910srpSPOlOmYo8tJMXu6h
l4SuAxDnJ+Gp3xySSyJg0s+nHihEc8mS0GURxamRgl7+9aGUu5TM+2Bn4LDzlXBFKSCyZPFu62iJ
X/p8zM+ZGByUAiOFJRGanxs/4BkJsCvw8izId+dYBSN1NKMUTnzj0+8nZsYdmR1w5a7fS0GKLd9k
oshhQMxWPnuebQF991oZGVm9JATeoaG/81dMP8Xwfg4JfCaku0CK7v5ysv3mgCQ++/ChKlzM2EfK
vmtSecCCvjLAtTmrXtzlDh2hP+Y7M64VOFVq/aJGx14X6FiYcQ052d9AAx+1Xw0ZU7PydBczRAyo
MpD8wwheBgSRlYA+uX69BucJOqQK2lF9/szxt1L4ZuhFZAd7bK+gjqnLCp8Dj96ga/R273m4KbFS
XumzvoIBTnpxXe4pdBIdXJFU8copv0PeoBwYklBS63ffQvzXyC9BwdpKAAtMizgAxGfJF7eIUJBl
vNuYl9UQxuIDJgsTRKFVG+yk4tXr3ykardyK8JTB7LpcKDX1B9zKk9KH3OdHp2bqL5TDo/jcT6wW
K9ajmJdC42vSlbbUARWsBcGlv/9jL2GHcbLZucvepU1dzLA5CxrojPUnxWJC6S3fpwU1XNBxDMB7
oCtltLLJ68ynQPjhvC/gYuIOuUklx6Cq7/LOYW8SbDCJUHN6j6PLn/s0cvhyjnl5Ioe8TDlgYhO8
nG2HG4+V/AuhxRWwy1oIbeofvdbRNKYjH7MjkJ9q2z7u94Ls7x2q90yx8Q313s8VI5Kra+C9WA+t
vSej5YHV3S1KdKdplTtNFgIB0u2Sf00XVl/Q2sQA0mS5yK7GbmxJzqEKO8Zz4og0ZanxmfHqUSDi
2KnDWTjwLRSLVm/PNv8dhwaiqozDO0yVTcTEIuWAIiUWstj3nD/nXOd86znCt9tB44xBnzqQCv/v
GkmgYKMMkcFh9vU5hCebipju0iilvjYt0+TrA0mcP/qaE4e2z6P3k0PCC2vNDxravZyL4Gvx7DI2
1y5ogi4bB7Hn0vmcH31uL4+7XAg0ckF4ZU9NxUG+qbEDiv+dz/X3IBlZY/I4QqcLMIkX0VyBfmr8
/BEEFU4etLt4KfO/uX2SDqScpYTNo6G+6P5tcmwDBZ6ywe7nBMoxkLGm3lvsAsqVTIqFe6D+HAGJ
k0vKWMHQL5+WWSG1lkEV1SGGZlBt38h4ZHeMCDX3G+twUfnizIJX2S06+P1VVG2XbhLBX32oNx+V
1KFSpwU5tVyyQRJWTWarYiDRm8uSRlOsIgKmQLC+wI+twpaE6iuF53XpQ2WuvC01VoU4TdTqkkgL
Wui/5q2ahKz0Tva2Xb412JLdBlvyNHrzY9hcM2x7fP4yauuguDggQoF9OtnXaOSTCyP7E9DE8uji
YKnBl8HEuYvBPG3nMaXbhQYFKzHKIFoLsmcqF/xQ0m3whj4ptlyR6FZ5XAs/dZCYT1s4ENJvZNd+
Hx3RmN+dvYsaFuQjKKsvFmdXkWPWrOHqI3/hdjJb87HnC5I7ieSsUkYxf0cO4YjUKA6TgpXg9L0A
ApBnrrZoaliiTu0+v7D6P2jn16+aGdM4BeZMkKrVSdiZhmSN4mjNNfVS7x6NzSFyqrape3y3FZvl
URcZWoC71dX3H1MeyBDJAQJFks45WH4e1/r9VT1pX6mOYluZQnSTEJRooZv9aok0h3MCbPqmk7u9
iSjQ93EaWh1PcLb66a52tvOzdj/jKX7lcEopYvnYCGs1lDeCDpSDWsXc/Xs+IhaMG5nThX99lRqn
fX5HcyTwoPaUjBA6FatSa1JseWccjOrRGU7bNEyvmmnQeAz9Oj3v+UcLy8p1vv8F8oeA4k676mhD
r7tNc70RYWOdttecO7ttlRxOL3Bq0f6SdHSwI5/S2gyTXGou6n9aIllzmptRBcmWVuitM+zNg6zm
uOsv6gi+ddc6sOe/GMZSRK9MjwiN4TiLWKtP+QowwX2YFovEIDfc4RAFiR2Nhb/9qW+6j6aK7F+a
lh2rbR9+X0BE6Cgdv/nKgOs6+R9lv1KVPm2oeiHEFfhYdjXS+YgX+yBtHUozj7YYV0OTLYBN5fGQ
ZzbnTDbNf3z92wWMK1eGBva3keaQXbPk5xyuhKJFV88lDd2hhORuo+YMJ93JzBCcNUvSn9wRZSBd
f0sxFA6Qdi1mvECf5IbOx6S2TwEiZwZMu8x8khe575WB8qyBkdYfccwDCF+J/KkYGksZV/YLR6Xr
ThNV7JUpH92zxRv7yELIsMzisUgUIzgUcb15nXnNaLHKWRFt6W0tytIURKPS73h+xqOy7VbHjSAK
ft3+dbp6YHtwoIaZgBJa2kOoeJviLdLoh38kMfHy7n9J1FfAIkUUMVCcrW1QHy+skFTUFt5fFLSU
BFrJ2Vvvw6FxflACsMLMTsZlc6ESt/JGFA2k6QKyAdA1stQzYDY/zePioWhBrxDUbN7Myxq1rLP8
j4BgpYgefbDjczkH8CVaG8kPIrtUrxvA+qhMPWjkuHgUCmI7HDwQsYOfWEvjgQj0f7gWzggTv8Zh
5rXVsC5I0dICHZywDunsZzmtuqdL116pMJA/mbs9Av6by7nPysaiwrtmHU7PUmCM3TEXigEMkw1T
YUi5saTP5w4aLFhkErfc5CFQ6lBgdrW6J+phY2fczoi4VV6jQSwNf93fAqBzDSDyClgT/LjHwM9J
7nO7xDL7OI6UDCnxS+n++8qywnicuVXIhmITYA3Hk500Un06jBQWpZhDO0/zBwfjAvQN5RTP2jBS
6z0VFayVOP2rNyrnirw8A5ssXLT9nhJiq0M/BuOOt+8PIFU4leKI4VX4TXlE75GGhJgzjGhhD36C
d3eQhRbFlwm8QAte8YRcIRpL+B+L47aXSfSa6eaGhppcgYMXSKaJQt5yFSUgP68f0wd+J8i2fjAV
1l5ektRYOmVuZzNmInoZjDMvGSj5bReLFesOcy9JBi6U4mGG3z/GIpPGSSGDuohyFcvgm+aaabI/
eGwHiBWLt/Oc7ST4bFwDi4ZhubZobV290I2pDmrYGpnaP+a/LGcLjNl+o1p+St0oJivcBKb/TA1Z
gq5JVRAiqRunPiiE9vVQ0d1y10UYANc7Rh+wsvd7RFkQfqC7qIr05uBkZp3PR3ZxbQ++kX3bn1It
yld9dOjGfrzJlEd4/UExghN3h8yUd6IFq2U7c+bvvYFJInVhT/FAXaZL+SgrCiRjPHDQR8NxhmXZ
qRrGQM6q2FxDsLBVlutt1f81grstn/549BTZjAsRH/LQW+vgfzCHIcmBjk3/jAYecwmM41YQlIey
QIfIkQ73HYnW6goXXz4138q0lGA4xe+JgfNTJDOtVK1nS6WLJpgjzq+1RR5K7n4vXoJetZspc1uJ
+NhFY4CGZzx8UCYsmA+Thy3sTFsNgZcS4rNrc1dwH5rzYo5NGlStT3/EJDkfNEHQpjU+qytA94Ju
IJ2m8snBbf45Eqpgka2/rDWRiXA3dWLjHfJEICyIwET14hxGQbnwXvCSTvddAf4yVKtgNzWYP8qq
9GFDisF50Oca59qL9olk45c18W55M4J52ZftMZTuZpLZX0z+OL7mGQP1stHHFSo/+6zQ7owAAg7H
RrWp0QnMNAcHIQDgq/fmtP5qW/eIQqY6tmqyu5J+TjWuiUuu5Ii5TFCLjIgDgboV0eKncKEzEV3E
BynZnHPxL3DlH70ODy0oizccTG5lv9rHYYadKD/PfokhmmG05ZyCNxSigqcOLfz0k/eicpwHign9
Jr2Tp9Pa6lxTXrBu0fU6NFX162a1pjzxZYsDqsFoGtCSBvODqnQvcuxncUTQC5k+gxFqtFZxaKD6
yAL1LNJeBmDkY4R0mFcW438mTHLZlzfxZ0JJ+UB45IGluTdZIdD2GtREEOkFtxNdRX3wo43Ty87X
FUmmwF4xu4CbRZEoUvluj0yZFWeA3C5XI4HT5ANcz0o2RPPu5thWZLGHg7vNx6usjeM1QcSB5xnG
C6jyxzRkRAXh//B7l0jX8kSCrHlJS8krozGyE0P30jsMCCUrJ9rNAZVqwpsT0AzAiieVtIOj232E
k59tjTYN0fZIs75FBvNCnvtx7jMM7j2CZmI+d9BFmwN8F9JxJmy9BR37BE3jVp1dz3nlpu040tz4
DPJeNm8NcT5otRpAIp2R8R17kMfKeyTE1f/Xz+NoH0E9XeEvWlYeopY0HTvYcw+YiEgX00qLhto6
JCRwnOldssmmFAjTQCANI35fqF8FxVp3D07G0NSe92XzmfxmyqrxtzJUrLAOawX9FGLTHTYFk+YN
knwY4wa+U2o+m579KhtlnbeidhLB+vmihAetf3xuuUTnWAUhayVrnrxYBLZGtE/8HzAV8Td20/rD
oYlEZEwIxWRi0rBfzP83CgFd8ZcXpA0wrjyKf09FnL1Ah0n+voSNnLmo4QcI2ONMXsiXZBfcgpXp
nb4gWlhkY+FncNVlvIOWdF/RpX4WdigK7zwSepXk7p38HNcPHPIE9O4xdCBTjIF6ftd3YhlDA6o5
zj9WNgysMIpYi/jthKC1Sr8a9MCuHAIKhg+0DZhnU7Vg/Zc7T44CpCmW/zD6FShTPcNm0Z6U2wMa
UBNVYtGeDqkwGd3cQ4Z/Mzt1A/qVaR+pA2Li1wUCnCbLYaSUlW+rzZZ3OWqMvre8nipXyCSfJKr6
BGmmylNs4Vgnd33cjulYAnjQasNdBHGBoOzHRv0aDpKQsPgP57ecZNboQqFaNM1uh9qz0+7s98Rp
S7dykXXZrxXJxaGfdeCi5lsAdjwvhFFkZpxDVPsVC3t7FMYVCNf7QZ+HHQcHrjC7FcGkWRvaf7ir
mHN4isPmDTu4Nrf3rjVKzztMYsBiaGKdsfRziMK5ukYVdkUkiX8LySLZN1R3UbZTQ1RXZs2OYJQY
Mpf0AcesnhAAhqXTH0I2/ROTsxyK5bJbfzcB59PsqBjA55p8G/zDW0KNFeqY0nYF2KATLvOfzJqS
sb0pNfn/AnVY8F8x3hDfgkOm7gGgcjGgkDbo3bWmsggxY1vsioGnrVPLhnT7Ruwj1RMkd4Da4qxS
We5BZppkPpE0hdz1sseh/1Ag2R8l7uGUEXuuXy9xqpmJ8OXtICOzFPB/72WpyKU7wssPszH18vwx
v3tRSW/OWvoZ4W4F/sHKrm8r4dSqIkU5ue164pmLBVhJQpQTwLPsQvs3DrWbDey7DDNZrNiivQPK
qmtuGT6kidRw1keI5scYWlIwHPN4FhHNai8PRpGxFNq/8YbidNEOCzJU1DZe+U0xXcW32wJXvkMS
ZupxCqsd6K9KktRV8Oh4RpjpO1Sn5uqMsRPUy9dqOsRq+Ll9LZAsMMwi2cOVfEtWD/sHYDdILbOH
U0Ij9ij2MRhw/hSDmtZNdnhz3b8JEZFyV7az5XGwpcPmK3rQocZa+nWgb7yxoJrgw/fLl1r89s8+
SWTpE9GSE/qiBKEm3I8ek+bummbaPPPs3ip/Cfj1VJHzZVpWhY38oEoPyaNfz3azzbwovBV5FXTG
/PCCpAc5z1Fyswx2SjT11tHSPFj14ghK9VMxLBjtvLD7rxk3LgBGAaZm/uhm4OUQZW+zHuzJhtMn
2pR1eydohd4l31Bd59wM1JLv08cFDHV4msaHu5oZwlklIaU/Cr8CLAXX+pkJnYAvGQmq8vllypka
ac/7SOo1oK8ldsrBeCRSfpxFoDXPx2ig5Koh3/w11MsdTIdrIZ5lQdAoLJHWV28EpgVjvdGHsjGl
huDOVZmLZqQiQisUjUC8k/aZNb4s6oFbrzIX6W30lsVHheDxTPVMuqD/0DOD7hEv0eqR+qYWf9hi
3QHN82VxIknSHwc5wnEc8DxiG+5KAMq3RWO13SzO3Zjwn1cgG9M0QOkt21aECmJtDf89+sAdMCgd
JKf3yMLYG0yMdeOYec4Zvov7jsx0oGgRTu+Luy7x8qCqg+XQmNrmcrFNSHc+AsxzAg+J04MZXZBX
Fi6CYlj7pPM38UOHo5ECYd1aYlT9U7brwAC0eicIPqc6GAzl5Eq324y57ZO0MDACMAX4bRYDfEMW
5fXh8qmWT68O1Q7YC2rNukGMqHth5hAR+eYUrRrw9X2j6g4HhE6SBY954UwpnmfpJNYVBEjavwgR
B5VAuAGRYSCr1KRR9bFGWyNhy4DKAkx49y8vDVcTbR+aI/1QyzMc/7hkQ8pOwktqUNBMbj8TEABv
NDEYDlRIK/72UmAeWzAylJYS+iV5WUwpDRRa+z57TU7wzlPx8QWLB/UKV84JXUfMWf+oI5CUTkAw
8tYPyRgWgcTdDjhAB9P38CMgLWj3BW/R9LhR5F3dHxi7BnO9rAHVa9TLeeD5MNfojs3ge6U7v6iR
24cKC1kVHJ/xNc36RM1SfEkV3jc+YeE/7wWMYr4BYLofBMsZzpHSHnSQ2mACprKrcugGrqB0afX2
7SqZbbqSK2DjzfmphlNF0WLB++oXqCsu49u8luVTvgOlLHfTHPv22ogdnuLktCBn037wBipxVhRz
XCmKnd8d1idpwy8s/jnXTWhJ5zszIfu1jf1/JvPN9y1U3WKAHmK+5L42auVHzT6sRiVDn2VvjQpK
/oHVFb82uWZndTCm0tzmaFBefGw3q3++E/8PUN4XppAPqgG+z/zfQuyM0xbtuEjFdEyyQ7MeloMh
Ms7/ft6OpZukYWTp4Ob+GnMfGyT0PYh5yamspHu+9CNo5AnrPvhsqTN2ttzeyTG1envpO5FBoSeQ
tHVTSJ00ZxWo9gIrXxlidbQBm9kDAmY7yRsk26uumNm96bV6aa9RnI7PUxZuVjydmCS78VQfZ9rY
YuTotkNjo/p+9wZswuh/hE/aQNoLuQjpBJz7MepKVzvsR8Cii0Chv/EnUeDJQL2tT0yxQEp2K1Cu
unIu/iiOjyHFZfrHTZSYbDTR31b8aGmRdwi41uUE0htwWu8CQV7KWVmi91Qy57e+gnvAefbRAM36
4c0Ah2SsSW4M3qggCGeJ1FwU9tvr2WlFXa8/H/J9RHsKou+qScTg/8oJKpKokXl2k1JXURzaT4V8
e7zo+C4tBeH3FnPRhHoCJmY3AL0WVilYd4iYC2RE6c7WX1hVly7Yd4deQmth7Nhdi466pDpFSTUR
j1rEzNpXGltVCG9HeRMp9oVyw76J/MTL7v61aX9i4ll7JO851PF3NILzzjxROeG8HmdBGEBpsi+q
kDsuXXlv0sk3F3Z2mjLYy/5b+9UqA8E86HOdEvk5BaKR4c3cj67yYok4VDgCX8SaIhIjCnxJokDj
jwGKvE/g9gTUJ0Kkqy8bnYiLZ+rkFWfiYGPBh3Wpii+lxupeiYn/I0gvXsbJYWsL7NfxzyqgoSD/
c6OCP71M+peQFyP/sNP53T2/luywKh5NqstyG/DjdgR+ihw+yJn25AJ1PoxCDgY/cWK0/rW0ieDq
SqMVPtVJYvyfSKhS3nNbv8gqluSi85lb63mBtVpeVan3Q8RQtUIL7fVATZkO2eJS8NdFvjkDbRT5
a8Nu/N+aFhxhQ3Gx+TQp5H1KALBl6OTQshjzOLUfddA1gOkxuswK0Xkwz1DygzkLibr1c/5Q70d+
1PrMwHJORn6uR7z9UT7y50NIMJ3sFqlF7b3vmWwwqZb8xt/r/Zz1914Bh90R613Vo9WW9LV+irgN
uw+ursjEW7sdjnj9EjSLDL33H/TwS9WhEF+ijkKFKVQOde9NOoOBYYxevfIhCcEsUKFEafPgo7dE
XuSc0DHhDpMM9gBj63Z3WNsuzEdNsEO02LHVw3VyIm5DDuPsO6mLflwNEo9UjPAn0qEgHmdUlPwS
8Q4UONdpK4pNiDSfc7pMdAcLui6K6xvQSbzKdogR8zKJ4gGsVq81bUDGVa5jUxvVSffBm/BNA8nZ
k1S6Pp883MxfPpqMbn4C32PG0caczFn586t5AD0azIR9k4UgFCQeb7ibO2mrLdDBRUlERQ590YXM
VlzMY+1RRdpW3p186yRcLqLspfuPSVPleAGJsGYbz8RgFxBYYshhCTO/EQLGTl86xlatxShDW31S
Nf/rvhRixiuWXtZA2e96ZlfhOQ2ktdMWBn2XLSLWOKSSqYk/MK1zVA9Wu0T/+WEKTfpguQ9/JKjy
jAbjIRG4MkG8pyGdYnrh2yX3eRhrACevPj3VF0Z6vaO78g35949B2itaCFJ6TLrbUcmpUdlutJia
U8le83dslMH1cRU8MO9hudZTVL9n2Ew7XNnnocyNvx98VuHx5ctn1U8bj93rkMBl81IBBH8QDuTR
qGyhP6o0o0OTfnGnRn4bHTrdl0D6OcI9+GuLH3JfrqR1C0KLftPoZIYr2OzHa2TjYJ5yTh5JiiGO
sW+mShpldjr1T6FSzidDDHGRINxSfd4T1wrn8Zq1+XCkAYkTKK0AKvnpyWBRUpTFNS2M857G061E
w4xKdgtnCiUMiimGhsRvoSzp5dvRN7NECfNgIiFMmR81CKQVVzo3DJUjeQK9d6HigYNvmbQzh+Hq
v81xmgJd4EIIZ4fUmv7JiDXVxdb0ciFUXIhJ6P6ko0gieC/YVtutQ0VjSjjck6OlsOgeiWC0Htww
Ur7294SpQqyg8MPOi3+WPzMwdBwaVsTWAWA1n9kvmhCm+Zp1YVPHTtlkrr9tbglXTX1DJQWX16jh
+Yxnf/qOqRwZAnj5M3zs6bKLv7yQc0cn9+f4KHwsNnpMYcDd/d8EKAdicBS5k/egVZ5l/JRVyLSo
bd0q2v8WJlMI/gABGpUf9u2uUL5lteznPbTAKH4EJ6O1hNqJkqyXJ7yDA+vO/8cihRGPm+GuiMaN
8Dv31GVqFU9+2V6RKv6tqXcGSDN/mandL6zcB8zvdPlrZQb2koO5sv4aCgLQC0PhJ9pIEDjoFqaN
2M98K/wEnlwSIqoyXcK2DomD4QwNuyB7SRs35uOLj6cvoxjYN65BjSaHVue+jq4UlRiuWnb1gRrT
w1vEggCfbGnUjPg2FTUShcCSQDVz6/7Irq/NpFgylEp9Pzx9mDnrwmL6udD9nT4+wGgwa/hzRK6B
RRfbFZCPOZIhiZif45NV7h5D48BxxCk4w/jm99FgQgIB5XXrfUa0MNIQKmS9LSLOONzbNU4FdS3V
jMEnZPRbsIV7xGAH/y53DEeSjNZBuUxW6yvK/7QTEI9CCY4Dg37sQ54Uv8/tQ8vH5b9X5h9wBG9N
ogRjUA5Tq9RSapJn/1UdRhTAd6sTMH9+8igw3EMnbSD/fbOBD6ini6qx3nJQF0LtgZTSvbEfCBSz
Ir0BLzgO5PtDYeZazmy2wRDsrZmpPDN6gFx9uHs8TOl8tlFUksa2qT0CBoQPL9UFla+a4M6jsLo5
mTlfccNPu+DTBazCnPs5+2+jpNm/LNtce2jk/f3nmyxRJ0UFg0oK2327pL2j3eEMvMmo2dmsDnHP
MqVSIPAP5uNYexl/rwz1g4v0YwMTkf/+cDZR6Ps3Pof5UQV7D76+qZrtc1ZbyfVvVwlLkEBsHM2e
B2ZdlXjg1EtE3VDj98zSC14wUCx1FSkk7VysQq9rV/2FaRxdp6vVt+O3FeCcXa7++SAohcl73lEx
FdQEZtApEH80mh+nxIWoVXfDGmHipSH2iH3O/QMOYHLioOlfEfkObWZkZnrJwcsjBhDSvl7lY0iJ
H4M6KLwBPWBJiZNus7uk9KZ002nt8vmroacEJVxlpAjgSqBkRUc+V4mpv5tRJXipx5UqiGyA6tku
206cR2UE+H9Ro9+pzgSyAaY3d+q1K9ng8B+1WupQiFbJZx0hzfoAs+OPjZ4HOvuxMeje6CkvCNj+
S7v4YtF3J7TiDgMMa/VQZRbFMi1TbfIkgzhK37W7UBdMYxHevOGJ4WoGSvu4HXKWhLUHRxcEZnWp
ZaXhNyzC/q62DHrwf56zt1I7zXwXsxPDCCgIObcHv9nMegkkr6mmm87EOb8OPmXMcz3hhXXLs1Ph
Lsk2251sLogM592tWtzDA4/G/hykUi1AtAhGQluHUoXhRQEsvv8blkHNDnO70tV7EiCGzRVDO0TC
PcybegdM8RnrrRladvVBbNpXPza9+QIqxL30mwKO2uo0ETY17+5/k/9FSATltt5ZnOfFuaB5YLIP
UbTlT4MZI2/tkYwc7y0lLPjQQI1MFscqe+V/L630K3lWtHTGjy24cN9tZ+vBy460BFvu1e8d2fMT
cpK5DEGBRJl8K0o4EHm7S59JJzj6/+X6rDBhWyZcZkvVOTLGxqR6hXSlz/HzJQBKN1TfPLOGJBKu
+QrP9pGIPBRbbAiPvKbMogSx0ocYBWLUlxu82Yvg/WbYifglE7XInj7Z3NkvZrtEjLB8fHm5DxWt
E5yuxmwCpC27C/PxCCRtPm8hrAYuLNd+O0kTZOofrt0VjIjGG/fTkz2ZJYGdqrvKVeUzDk+9hZ9y
3ZGK+oOBdMBQQ4T0ASTJEeYacu8rjF0DLae6RxIt1/L57iQ6jzxmTfpuzzC1YLPCocgDQ/h8WdTl
J/DAAnbaOd+szklIQr8Rwaarkc4c0noEI7viRBdUCj4B0c87KUV68S7hwm/qIbEAoWc8UYjzj3EL
cbFfcoGsiVtwFkfs+hU/H+/MiZrmeHuQM1eYur6K27DptJXjgMkOhgr+PY8UEHOjdn8JypsLlLbX
t2esZK0pjiuOPs/Bw0EnDPlML9pgt3NgSbJpxK+lpvFruTzkoQR00vgDVY72Fz/AwkCwYM3B+Ez8
amars1YCD3Omz8/H1f335MvqUnmQbPtqlm6NVNbpaDc1pV8ohxDxit51ilcccSRzRvOJXawiqq+5
cwAnsCbOgMTdwh+is+n48UKgAwCywRlWq2sl8WQRmg/isMeJkDCHd9S9ZEyq6IJq48047mCcimU3
LZAlZK0xp1nILAVSw8iaySXHt7VWinFeRPslalu4IzQZ2RA2kqJAJ3vG8PaX3pFOCmbVCqNZ5mwB
pzYHGAIz/qIGT4fcv8gIbUpIUkU6XAJlpHjDDmOtrDinXqB1JMF1coeehl6i2y+Gv/CflrXh83/b
oWwd2sM12frW240JNJtI3+96s9xQ3qTfdWofio5hL/vHaC0l3DAEmWPriyESwvgsVSphBMjRc9zf
WH4O3OfSZWxbXkVNq3lAGAtSayM3LM6ONWlBgN48HC2ljukQQNHtmzqsWFYjr/hH1dvNwpx2D+43
4g3+HCI9smXBvkYs39UIo0/yKchzL/k4+yhxuz7OkQOTJbVGZcp3Jk7P0GJ35/30S55GEaRYMBHq
53men61Ad9S2jSFQ+ms1KXMWYmIyXUW8Y7f6iWxyr9PfCSgj4XSAs46Q92m/5comXEFxqz9Oy2mk
srQVIRdOrYnj7/y9GUjdPEG5/120vRidxhu8znNpstGYz5XC77PRfJeX3PI/2/IE6cV2OCmdlJJ2
vBzbjZtP7NTI+DWfbGGBn2hQtY9oLAw/Ea3MXnOXHdT29JGDOmsrtsC9l8TO+o+bm04YwlZDbiYM
GY/Z6mzKvJrbxNup9Tezpx3LInRNCuNX1RsoSYBKeMAIWAp0pndovjXgzNIQvjk0SSj5OLuNn09B
yCtxPfeku1lPWhp9ZV7crpYIUZX8F2qTzrKfhNIOPKcj/3tMBtZvSHbfLmsiwFHadDw6LI45geG8
Qumkw1/py4t1t0d0cN7MLcU0dnZ7Hrkxu+X1TIwgkSiN6/JmKV4LbpC/KMJH4r8QT6uNWlp0iyoi
mwkDRvnWF35E2HywGLszL5Ue+MRB/yrWl7eTfILor7H/hUEixirAqaW90z7XNZKYhVQFQxrcmSD5
Cxdpsa++ecQhd9m1Ku3xzDKPui6dyWdi54RcBiC/h71o98nOvvBZV+eaTR24DiuRAbiZ1fRsf0nK
BwGglIdLybFJzpm3ZMhuw4NIwklCQ7oIbBaaHl426NMGAeqhQXOIogOzdu0aomWua7IdFOfoXFb2
fHUDq55uYBbt9j5b215YcnFvJ0uOJwIBf31IRon9LZ1C5c5TEbb4VdKYTPVIZcjrqMLTi2axJ1cr
MYvz/u2KhQjX9N6uh7uik7KfF8tw4vzFncEkO9Q7T4o3iwzZPyZmHuwjWe9Nhyvx49Yk79LiHMK8
wzF9ygiWCz++WwsQcv2tQoR3CGYEp/PJznFRHDTMTQ+tQi4/qf3IGOr/uWoN41zCg/ppvCi6sk2i
tpooUiaq+LDtJymTkS4F6R4TqEb7vQQebjjxHAqkuDrrPrBclKnEWQ9j/od+80s3Kn1H1Oz8CYZD
QtaBBEdIgT7Wvg0dEJ9VlxMa8OiuYBUCT0HBifxT8yPEKVuTFR9avuHkQAVgY+xDsI4NS6z2kD3b
UOitTljwOdSG/nkD0WraC+A3teu2sGLYSjoxBu5wNxNcPx/lgtfCWC0YipxVONB0SPl2lHNy4tv/
lk7YMAKh21c7YC0rmNLgDFhi0kUQq4se96+LCdmUhJAWv1bD+RHsseXEUO+Y4cDzMefVpHCMxkAV
IPKPHkrw80taKFDFnVBxJRcPdjTqnFMgh5ozBwCGPAr4UmcD6G5lQdmCks6uhinhuf4cA2EFNqzo
gkydltaEOzaF9TpFB7n5pYG6oqAsdu8encAP1SaieUUfG+cc964dypewakhmld3f1hKQt8rJGCzO
roqui49M2vDVgpuX78kBe2wDLlHX0+JJtdOhOXE5FQ/9Dei1KYEFB0oGTbcVDejA5/VD1j3i0Up8
Gl0v6DM2DxjNM5nBmJbvnm3nrHAyN8OjuwOP5jpxZ9hECrOQAY+HiceBMWySTQn4cBeLCA+Sl5uO
v3oU+aCr1RKoR0p41IbqhwkOTrkVi3hKkCq/DyrUhvjgyvabocJNLi3olTAUBw4QygxzxakFOnHN
FfzRimeUjs4JbU4vBWEogq8O/A++VkP2MqGWBARxMOcvcNUx4nwXQPAJmmjPA3wy3vzERRaOOGzm
/QaIwGIh6acgeLlVu4bCs18BXkoXgCpw8RFpC5SpJq26VZycvYR/K5JRG2gb1mSFFTwxP+KY9aoO
btjuWQ55Tft4m0CA+HJ2or7x7Tb/3ON9BJlf7dV6FnKHE6y5mku2XWJdoRd1cNe/OrDLdsIUgHjY
NEAov3stfAvWJjFYxRZwBQNFQofgIMzjVxKY+3Unde9rZ2BTkZbFkVSHue+GSNbXBvC6fwHpJ7Q0
FaACVhEZA2ngUVBALoneFDfiCRifg0iv7yrLLSpaFbdY1CeaOhF6LYjk2crHotkyVLHadv75B8+9
Tu3X9Q6+yr7cQdd+JjRjZV+S/YTdS+2j7lifLFjkX0TPwco42Jy6SDmYpCJdW+MQH+kZvs+0/z2F
7Ebj8/RvDL22QOZVBg4Prt6xwQ1x96L2mGGIO2us2EPneSQjWJYLyPtru2O823ybn75WhwD6fQLQ
DDcTuNAtl8p0je3a+EZUtYVhCZMN17AvkL/PN0reX2A9Sprs6IzBoTbL0O2i5s/zMB7m8RsSsCBC
ZVLPAqW/4QxAuj/VsbtxJ4+5FvsL/5nbyLMyfSDM0rBaVD/F0/8znkg/7O73aBcBJK86JqACxhlm
3/OKqkPCTxWC5daNpVltNKewjiseuo8SXl9d27TOK4wr7ytQz18fukQ388pJmCOGsKbQ+z/th6XM
ze2bx1TU0EUxTt/tsTsbUk8s/SaPHwPJnhNuyg453AKQ4L3tCyg9zqrYNSEqyHSBbfMxy5qtWG1r
BqXHuTs0XhEo0kloldp+GQZCBjGwzFK2XzcgnqjmoIGQwsO4E5ZN0OOCPIAFuUUzHqZWOK3NLYQA
9XGBImUc9YUqNxxFPaqcWR0QVwFwytaZ50BwBsALI29/wJGsvD/AiXKw4ijKrz7/wy8703Iv/0iL
zcCGRPzAn2AnTKTewYcO+vbvNhl24x89m2O5GRIktp8CLgmPw9aIZrQNZSk3U76UMGdWEFyQuvsy
I1H166Yw338c3RNWIiuBOdKGiiGJ4CKhUb7yi9acpbuu5YRp0cK1EDVeb07ZCCVBAK6DZrKjQqIp
iahpv7rQ9HNWeY975Ujnnh46+x87B41TIUJEhGfjRIrHd+CL1FmexKNmocJATWU5P//OWkdZHaeo
LSr+dF7BhUkfG/ZZOdt/aTSbZCZiNIEt6uydFVlKyaF9BAfhFM/kKOVkWniifPCZwAUAq45dQgFr
sw7lBPrqlfTXUr7CE44noGwT3pe7Zdqv8ZPnnc1XewLkPSi22xbGkIM1rOcN1MOuCNLEGHigxidT
dG/JiSIixT38xf3DFXRiGHGwTFRNfNBcjlpFlNH3ZXJUCvQO3n53/P7+MWhMx+eqi8tEWU9VRxhX
xfxGsgcUKBKLc2VVsorbreAkRa3F2peByV9BKVu1wYE1lRAFRR3PYB1IBtniB9ikKC6DrsGJHPIu
CpLUGPvt0X4fIdrDLAWqLxVvCA0gsdowPDQisvU/YBqSQxFjQzbdjICrkckE9hywlEXmoBuDV7MU
MTxhaFwjulpRcZlahzGLR1SwJklDBhie2KB/zKn9R8Y9knGowfsLgYXsWDhuLIDf/LvLABxx1Roq
/0dSXxWwzSLZKtcwZQVECkjDHw2aSR8qLtoDkDqa3+pAk96YoiRDL/z6LO1EDfHEToGZI/iWhrpw
V8CgYiZEbOJrlsGKOI3tv+DtK06oKdqnKBRT9S7wdfwg7djs+sxXgVTKNTSlt4SK6rhaUfsq8V4D
+9hP+K4oZbueX/e0ltKccxL6yB4u/fNM8qhvSN1mWAylHTTuedHP712CcPM1SaxDaMvBSUsb2cMu
gmUkkSp03XfZkw4X8JqAE/kdetmPSSp1yyuSOcePQClJU6VU0mgM5dpiN+kojtmYlAY0xMh4IhBv
EZZPGeHTkD6yQu13gycKDW3SMrKLhTHBVDj4bSktikk76DNhufklrtCqx+Bx5L4+SKCsNTyKQYNJ
XuoblWLLFkBhc1yJN8OoPNWxOB9NIC8UROvxLdnLZoLYj6QjHz+gHHIWfipPzlBML4a7exum5Cm5
YRBaIgLFWEPYjiQSRyJVTvVVd4LMCGURmTgono0Ran4mXcEsvc2Q/dCZzDx+T/loqaN5dnTH3qdB
0SYKPNVK/OhPGKtJdrRCWRfMjbc9YH6C5o09txRC8DIz6x94iWFDp1nDm4kiYJnCMlfK4ya9QfRI
WSl35VoUmJdZGjuTIXftN4ioZu91uM5fKXutFgB4ijUZU9CQoWP+fFt1gb7GQtZKOYbKNqfaQDeL
lmgScxOb2KzERwSaSAxYFHEt+FdmvMCpVlpGXuWlT3lcJHwbRRASGHDOlEyg27rWv0KGTvEKLu90
Rpr58d2R85xt/aMom2dvnqyWleRVFC/vsVTNksGFp091kMmgENqS2mHW9ofCRvx5Cx1KcWLbHcHL
i0lKHjqE43UZahL0U6kWWJmvG8Fw01ZqWP9dduWEvL6Cg8qr2m2lhwr/DYmz/pJMSFWqfit0DL/y
o8V61zzTe5GxhHbSeRkE3FMeC3uBachuLB0MIBX8Yyrz4Ez8/A/b4sC88r3U6eQeHgJ2uz04IX8j
ie/sgTPN2tImzu6SSb9m24Yi4nA0nrZuGbGA59G9qLOQo7vnms/6POF2VQIObj6JG5m+TD/9mVzt
GVR/Yca8uQ/U01wLFGk3iTFLI4rbkAoAo0o762wwSTfG/nFQUugszhOeQcLYkI3OKYg53TFoEWcy
3kUVHmgGOwChbdkcgbmF7+lfc2ooCUP/vuIeurd+TUZ3RrAOxdEdGwDKCZiZU+eTeJ1D5zpm8ZC1
3mzW1sq9YTQHJNKevXs+08fkanqUzxvfQ/JMOJ0GTYJyQ26ieCSHuD7BSBFfm8sHRXzJZtpTd7OP
UqD/KdLszAGEBGKPnZqt/T1DaqpRVjXFEcg+43QuUGrd4VuCjNXHsBAhAGp9t0QJy2UZTq7ZALZH
8rw6Hf/pD72il7cbN3Y+tzec2ZqDW6dsRMbBwoRVnhDqelebKBIRcK1DgbN/rEfwaJBY03SY0bhc
Nvddi1RkIFoSkAcF3rNEIxw/PocI4tXNk4alTnft20g1PBJtX1SK6SUiW5MwO8pw4g/XAC1/WZgE
Lr4tC6dRP0mnkaVpaLrEk663OWIzl/Fae6HNrtOe5IqJtQ4Wd3IkJjYDn6/Tgpy3zZDcUXfdu3Sl
DgpHEt33MMthgPtqLpL4QCdl4iGkSEKmyj7NFdjACLhohhSFMs+PxPl/cmVK0MNsf+PIF4+oLZ4Y
/lP7oeajQImMmaR7njj5Q3x+QFZXDBbW0dOmxAccIt3+gz+GrEz0INF93gda/88JI36rJDUo2bYU
1yAJ8Tb6rrTZNDoOfYa7cMB0rXrw906Y2OsPtPdnBNgxmjtKYmS1xWWVFyZuyxNOcHyEbX6fExSY
+v7b334O1I5QijfUYit1qx3vD2b3WOi9/kkLW3TizPMxr35tMzC+hjRmT0I7WR4sgCRIDtbliscd
SVEYKKcY9Jh31F5rmEpQ1FHXY4ryjrDATFSRSvDpTsN48r80zBl4CygDnheKKcFd0LXZGBFVxVP6
FfYSlebYONrjD6Rgy2LC9R0zJXf/whb7DmCg+hCr6aSXXKhKN8OxS8WgoQHXSWfjhx98iZvOdGrt
nRCdbC3O0z+qFUH7kghoWyDNS3XBW7wqxnbuFBsOP6PGVHJMxtnaiTABJCJ17VVxwtBUhuymvc4t
oMFcwCBFqmA13uKa0Hc9K4kF4ZivFMuNqFBlJ7ePyulj1Tsvbt3QmCbJ6gu8Mj/xPwJPVk/YIHsv
CVAAZhI3ae/PLeEnf0m80xF7h3MlsdqxksihKwkUtHVHYTOdbcMsRShvSZU9NNRZ/+GPSemLMFee
aVhRgkxiTRv8iJvirDLOo9rr62yAmtRk6fQsSenVtZHrgIY0kornSNGeb5zbLjXjX/6QEiec1Z1A
GVG571vZ+m5XxJ+OhClClU69WjpE57A8j7anHMI9S6zNvvJRDF3GBNUWXrjdtlSlquB33aVUFFkT
eioGhc3ctqH3PW5/saGA6W4AqEhxOXeyr8bddVAjK2QdwVRYXgQ6rr01YkAmDnEn4p50nQV7yftF
ba7g62A4C9nD0z67IRlVVS292iYWARN6dfGIuu1exlvwhbPq8d7dd1XljJZQRIlFglBKCIgRWfSy
vLGOI2kvB5RAg8L7i8CbExvBabIaYa5aYYZ4ZX29YyJB4b/0PgdzGVeXYY4ej2ejgVwjdQQlcn8m
bTvLcREyxLTFIPkxbbU5DKIosKWPoQwJOwhPANs9jM2l0E/WqYBnw2zMzxZu+7yXYlLc+QUbQLWn
mUvRSAoIuQvTEzVM+7o9KwvNktT1PJhvEOdpRUyuXB2e04JwgQOTsoZZBE82ZcEjeLrBCUU8yh8U
eIzuExF6sbiq6WwjXB7ywbmyqkmj+5d3LSqG/MkOVK7f84XEMdbVm02UrsEWyEvWCzshShpvEm0W
oedVwHb4K4MN1F9zR0j5uuCnLonO5eEs54MqaUE+Bhbs+9Y1j0jU/4PEW+2BvcFs/x5b62RFb0km
EXXeHusDLLJRZTx6Oq9IFh9PmUJpISyVnwXKzdMQC18OoO3GfsEWHde5J9/xicybRI3LiwijeyUX
ExhgXmqQZYXD9gKepnZTGA/nRTw5DgEBVS/dOtrQW/XWmHmR7kqUwp8+xaPmcqpWyjCm2P1QIUg6
Nta8WrNtIKhYqfp9H6oxvDT5cDv/BjDRmJsplyBNqYCQTLMZr5MmEZDtsZF2dRh9Atdx8eF65TAc
g7LUjVyM1H2KXkmamfLgJ5TNOfdjZ5se94CUWNW882ML+1mjR+YWVLfNEsTRgsZ7R3NpDtOzBR2Z
H1S9ExOwgAsv+B+b/nDcStbY1pbQdZb1mkhsFDU8TzP7kx3UHcvAzkYjEKU+GMH+IaBec8ZlFpGE
VItbT+vqfbi2AFHxbtaLNYhvpunCseVw8D2UfDptOzErg1NUg/eBDOkcM3UwVnhN+Hse+64WHGBf
GvFAD8Cn23045iA1PMAV4C/ZN8eAL3Ax+E9CEbRBNEjpe/fxcLadnU5Wq4YzIR+iqJ8OEbhAoeS7
eT5Pkl8D3DjmvGs56Fizha1ELj93kzTPU6x+7xB85x+Fs7ojQIbNAxorvs5TetOLUvM/NDb+Gjkt
0GK5WtzSDekyuvvusB8HDvkbA+vs6dnF/5tYU9ktj3ImVMHY1Jj0QRW9uoqQwhfm+CwfyUj+93a/
GlvEPynjjB/42bqjQ/GCusHy1nh9lfpDLT0KQzMj8Cx9O/q8NHj7hwwolqKEf5gCemp3BOflSP/X
XGxHce4jrPLeKkOeIOxOMgbjASnPlOFuDx3qAdYUv+kcGRJ0evYg6MOHelONgUFSgRf2Bb5QqRt7
ZnsqxfN/gWqFvYOkDBC67H1jkF0pjomBTDMBb1442L2eakRY47VIhTogDjV4Zu49f3N4ZUq2etxy
2f/8+josw82iuIV4PA7EpQ2VcXrPj2y5ffNlWcZyzF3b8o45WFr+/TZVnf0xYto4H1JsNO+M4VM1
0gh6L75UAt4RiB4oS5ssfeqY16Z7hvgxMdUbXB1N19xozzd+8UMWigTx0hKzwHg0/JrmQEjRl7UX
kuOtUlxGIeWq51z8ns5E/kscgBfbZfU05OGvHw4ezk8WYvLi2z1u5KzfGeHzLbbMdZrJ8EmDWtuM
R2jwC5Qhg/md9BnhYKNMGi3DXejpTIZpUANWjzWEQk33hL1RX36nfuyLAG8s0LIvHpLxa6OaWwEm
NtpU2OZnJsfPuhN43JigwMIQyAq/tPPA17BA7z8PfbP4RSmvt/s4Vm9ocVAL6/00eX7a28NEy1Gq
uQnktx9MPjCT+y8s6lPu4EsJ5Pj1Mab4XU4ECDI12uzscJYOv6vLfBgJuAHyuSjd21wQ4NrzQ0/E
XdjvDr0go4LZGq0I32OwlIU9Bdxc4RYsi2DQtafJF05QHp7dTPCpa5VXctdmwfmpGPXjN7w3aOMz
bobVgh/EFONTfNlbgWHX6Z3K7Ait9f3pJ4W3S/p7oaV9NZdYw5/S41p4Ytg0YdqOxA1gSL5e+Uiy
83C6QU22D1F31qlNepwVojWPFHcbrjlcO/pkhrdkUIyWNdFAnAjZaEMqUibXEFes21MqXgiQl8ko
HQwwDQsujKKokbWPA50vXoXSPNy8fl0PTcqVQGwCHEGmHiEeG7arhdU9LYHAj9co3sbgndBrkZga
u1VyVc4CXLF5IJosiB8Y9DK6iZwbl0XhqeVM/u2d5njvePNiXAQshA6ntY5VmM4Mj/L9xo11mtJe
qfoJbNIi78gJhT2FQNy+x2OV8tIOe3PjFqJoG7Dd5T4/CjBKQWZxEZrnd6oy/in3EwnZDOxy0UWh
5JVfmtkCiRfOd+SDu5SrtA4FzjtOaabQl/xlo+IIoA50vQxk/Yos93ZTRVi2+GKGVfxShA+bPXt7
gnk8bwzMLx3rpw9EuJqjZ97wdwAaH0nRqHGClztOYN1oSgNCdyjxtcAZosiiISW9UrEYfUQKWyJs
SfhC4W/pKGhEjxPuW2YN3C/PkBB1kjlhgUAjC74CYkiQSjhXGjUAlnNuysLjq3K1XkdCFjVNjlFQ
ty+OZcq5RNfQ0P2iz3zB9loxg8t3wHAMiF28i0QMiJ5HC6/zlUjkNTIdfA9mHHnXoDdpX2vNjoAC
l1cG8vc5MvR8nS7yDYUWxATBO6LSE81kvh2o87Tj2EhRTnB0d2FEh9ba0RJ/+akrTHzgx22MaxqE
EDXSgzosu65/xIFOlhL6dsguuuvSwxtLtiTOVcOpKjbXSAavdfu6MpZFSvhwl0pjBJYTXJ9Vqy4s
aHBIWXij/5uDs9JDFEb17LzCMphXrHNOv9x4eW+9d/7wzfVj9aFbNZPZgP1ZPb8EStGb5nHl3oqY
kQnaILz7ESuAhAbUooXn4FH4KSBKnXG52Xz0CJLpSBkYJwbjXoHdTaGjzx0FNztbvznNz+NqQYLz
Us0P0Nm2e2j5l6y+0Xu3HojghS/N4cegwt1QKlvgBq8WppsLjPqUxiHdhOGIZWvPWnObUV3KbRG6
y6QtxUwHWcqCNeJJyPtpvaqcG4/mtIpVch89DX02iuG79bXlO1yXPp0QDer34me6B/IxNpzM9RM9
96d0Fz25GYaO9KEIe9hZNGJPcs3jnLOkHACjBlvdcXrZFUXp358rLCppp0olCH+30h5zPv+7gLim
0tDxXOEQWtoChDR7bVRyQCHsCEuifYEbXHDxekJu4DsPP6W7IJA35fH7KPGRUaFU4+ZevH+5/E3A
wMBaMgDzKW8Qdge8d413/QqF6SPP+JnVwNoozn27+RfSecGExqLIJBMbHJQSuXmJOpwK3LIhv8/D
UJQRYmTdx+C9kyJZNY5G4skl+F5/Q4Z4Sa8LMmqBX1EB5i/o19em0Pkskdsej+iUxn42WE8Csg7P
ua59ZyXXTIDrs01ciNc3MVZNa/YQuo57s1tWiMneyYi5/YBU/utkOrrG1hKY29/tZr0a2/FMkKQi
6HBrvLVuJT5vTNyGeBiFo4TsSsHuWCMFn/++OuGxi6YNiKp2qpJYaly2jnkUmhFZhpdt0zypnsuR
WkTEw40xGurpj1ZSOCBZfG71Eueb2LsCIrHiJirYaxguV+7f4+Uyrla/5NjsOS1M/KpgxUCpTToP
R5TK7VVsoGSyWHVgkHq/SUHgJg6I9oxPrwNnrowzv9krrt3AHc5XF/qkCewgRU7TaEAbrlUzr2Ho
WVU8qbe9T3uyaUxWVvYeqpw0qn1iMbnxPGRR8IzmAkk2gjW1sLJW+hmtAKzg5cepd1fAoNnMyz3/
yUs1pFONj/Ml1sUnTxVhezz2r3z5ySG1xMaZA3fS0Hjc2rRc41CAe8PHY4PIByPq4+nudfdbxJsG
ARBReehKaJdc/8u8iVST04MGj2RzMh5bF8glXB/XeJPG2XFlTDPiW1xNEME4GhSRCxA1SvWM7A94
B6T4MzeKpRf6ERoFEK3PQFMYw3rshlOsYxnwM+8p8O0JE1/FHGvheyzy4saajnwcW3dI2/Uob+In
MVXk5Dd5fAaMw6fRX42kwWFzFAhtDIDJKvRyYgtwtPrBpDk1uyGC3BMjIoa9QtF77ivMzqSroh5e
QesmZwmmEuaDDe7hS7kkaTgmsfA4tiI/s6WQ75d9/yi8RW3LN3b/htegNYGtnMRzwzu1WAKLyAI2
DLO3Zh2BrBPXptWOfprkhR2+jGAw2ovqt4vAjb86uhOm5XP6RfgX8ju1W0dv0Egxf/3GRdWCsczH
a8dRdmU5yr5HQxjqYEMgBojjt5PwX+BLA7SRB69jwIZeXdM7Y+xpLp1iha1yiX8wJ+G1bjUOSuku
lCesCVpY4YK0G7UAGgbzIcec1wfq1luT2wMW44zSYFT4gkVLSgwDVXC836Q1cwf+msDzaA3dO8yR
XC/lxGdtkHVkzocJpN29YNOLA4XtZHdpnw3RhDunTQoZ+Li/UyKUKqb8srVpvP1T9HuWarcUPdPV
jyJJL1WYiLFPddGsbeBTMm39BLOap9/jZf8jzv33SAGIxiNm+IteGLUbEdQ5rLHszpZZi8ooZNjO
E1LPauHJ1TCG1OTwLM6wyFbabxaD85M6o0y/z8zWvk33I8aFOX0Crdm4SEdqFXA0Iro00OvzyxAO
5r+5O5ff2+yIpwSYuCAYRzIO8W0ZlrBo7DdDF+FuJNc1jTaTHw22cStFhlx9e595aTLJ1wdUwyYA
VvTplHoz/G1mWHXC7pVb1EGFPS2cvXLr8CjNRR+T/vIVgybp6jo+JchV2bImIx2PiA8g4fDMhHN5
jNpye2iGTJKmlqAh2Q06heJj5iFwjU8OZhhm/puRQ0Tu829/3RSFU7RrbKHL4sUdoDVudJOIvpSs
cYL1FoDQgfvmBK7B84ZyuV9v+O3EW6RXosi9NnGpyRVUHMIIHxnUunrV1g8sYUe46OzWp+hWpLfL
t9Y998sT3YKMFbUl7KGXNBg4kQUnLuYVoFzLPX4rAiylzpCspmbfysy+jXm6Oj+26MXvaWhySJLZ
Jm7+Nr4i5jRDQMPRw/dTnIbQVim5slwcA0xh1iB/3vkfigcVpp47iVi/1XVUmdfFOFxc7VAe1X1N
vZcuiOy7vHkBwYZ1UbYhOaBnQDIIQxcklPmR0svnXsL76humT0eI5wWfcQVJ6hn5oEDIByBY/Eun
csAj0mVbhqPneOpARdGoKrqswkhdvhzRObfMv2vLCGuge9ag1MiVcJ6/gyK9KtWZ/gEbEFjGG9vX
hknyOC4M3mA5mafJJ3nodS/6eyeTsl+B/Lzrjjj0OcmVYvEB3bFOC5oAhwExrBDKzwWGRDm8JtLO
71NWkoZzaKPO4xdVYBizLvgTeTvHGc4U+YphGU3095cqc1haaR0/oJW8YCaJI2V7qwdAsBX1xiVA
j5M8bqsTFBqrUbc9TzJRUm1c+23uPS8ZKxX1ethshxTEVk1yFc3TEeI28hauXJmeBe4+o//FAE0O
1LlCCfGJFrBQ1uG+6yat/Uefktol3g//asLn/Us74yubENK/staw50ORtD9taSGyfjEcqt0RBXmZ
fJV8xPxIpbU3Epg9x2mdWiGMnVc2+2k/PB16ABxHHvMvTkOQdZRZi9muYf2qUmS4p0lvEmly26UC
6GdKMFAQu5V2wcdeWvevXhSD0Qy5JNqTl9mssHrk6e2WOSy+A9pNSOXFJ35B4J4giLikHufPQmeo
ti7/24dvtx8T1NEyzmcYs3pogeDUYVLF+aD8NOW+arsvI+VFx+r7vvV4O2OJXCd59Mffk7MFHXfm
GYC1d74Qyo3xyMjpUhDgE+Z6v0EWkU09kk5kYYIbdImVGld7FVJOyQPzvgIZqqlpR2eKPm336FP1
APCPF0IVOo4Mi2jGYtfoZOg8EJVfhfib9QB28FdvZdv1hLDVmd1GEm5aOxoFhZ23hNNZMnvSubqe
gZJsm6aHp6h2lSuod1k9QKHwvD8tdwaUcg/Z2ltwAF9pcZ/lSopWuvgkxihoHDstvU7YJT1yINTx
Y0IzF0mGgrs1hiFK59D0zrTT3PzOVxqfyqd6totkI9BYFI013VIiRITxjEuCpVZ8SCWXx9yAxdO5
oelvfQKQXG61EC8EbQMncBf115xTx9dgHky1kI7bpIQOzS7UOyKEiqZnVdsHwqzo3C+JYFBOXm4h
nB/l81+cJ5VQwhuY0u7YX+R1wM1lJWtkBEMcZmkeOMyTS6EVGia4LLA8nLmLBQfFgevfHUegG39U
clUprmmZCF3UU3bQMY0ikUPkRnJ6v/AkIf9mtd7gROy9G0hK4Is3gV9LdSjIHlWS1sRKyz6OfImT
EoPXpKjBzB2tMdtwrBwrkscaTUrT/pyGQlK/F0lujjrm7w61VcDxFZGyNoM+xHTSjXpLj3yiIrcu
WzoffV9ehXLEDcy6z3Gq1zuvdXaQrWnFca/mMu39LR/XdliRN+M13HG2mJwKohgsB6WtcQRkIXiw
hdVHqsxpjVB3p2C5IuM7auBiWMPI9Hsc1WOgnTl4x4WahhnVp/cPkWWKIfuCJb4q+KFUiBpeI3Gh
/FdjMlKMexZdaOg6lMqLxpYeCjyksuNIc8dyl6VuVrihO9K/TzCoxLfXuFg3L+HVwXva0uCAcO6i
+t6eyHqmEfsxAMt9DSyx8VTy/epupj6zb53I7bzGqQqvBo2AJ4aB37KZhsoLt/zWzxaKCiSGqXqA
6IfnKbKumaKU8+oJG61WYzGoIJcS7ONvgEsiicIXGEB54LqBg+gFgwaTB+k7/l0k6TG0LPJ1/FeH
6Ko2+CEots29u92D9yiFinBZQlxs+brU5weovNJ/ke/WapQ8yyVKZ5IR5mgak4mE8TMRHzsxL0en
t84kvPLkBjH2qN7SBrqxrDzspd2iv/uh1R2RnOcXX8LBfZsL5o+WAKPr/n6uUTm8w4zx4zq5WLI7
xcl9KsSckhrnAKW1fUxjR2hMcjstN5dXfmbOUKK0CguMm4y9f0YnlXchuIGs2NE83SE0s+9NU5PY
pQrBljEZu4ycJJVYygLajNSYI+cL8MiXbQP7CKORfFbSNgGr6gurlRHUd7MfzzXu8AnJcEVklDRG
snSfSVwlZDZgiHv6+1UwXiWxeGerclcW1Z4+h44C4dMbdyY4Q/1XGfGxFQIICpA7VP5K44dY84H7
46o07x/3Cvtf+7PFGWodI5DsYXHKgigWrtuVXn99BWG5dpGW1Rne1gIqurCZGompVSKqMSay/pza
H1McpQiMHuzRm7mNzL0ru0/a4yLRseqQdJymIABL23Dt8aykElUmyyDESgSeeXGwd86A/CTa1n2Z
DDJD0pPOAAG80eDlVKVSDLXxY2JaGwrXt6hjXCq8b+NjmRMUts/RQDzWLFNThdEz/+NkHTpZfrA5
NJVgYU2wq4M3Aa14YJHjRMzUggG6d9zEEZ8GIiAst8dfVwAQ4KLVNVwKnU0JVQp6J8NME1drGKqF
u++sXMP0xPDFG9f4iCYDBBc90SdSf7j4jDI/XF+DzdLsChK8TKHGDyKKbOZqCz8HLuGr46zq4ZmF
IiLyi9BjOPrkYRioG3La2a5DUfWzKOcBCdGrU2Qjoaj7WsAUAtWqpxfYBqf1U63I14XlXJnLCsQ2
xRmaP59SDohylV0A7ExKMXTxMRnZXn9WsoC/uUt4juh4Tp7iEircqwgjgaFqTp9NnibwFfaFtX3Z
wZDs09t7D2MafX/YSYoQOnswIQE6O+F5GvbJQ/UM/tcAgp23k9awy4N406uzn+K3+VDxWtVedVp2
sNvfO/7dCv2pYhsASjw2VZ61G27Pg5y3+Oc4YtYtFbtZ+L0sf5I5fdknXTU4qR81944/5cLMa6OO
jhhhRWigUWM1YLl3VyOqhNNB+MGwtEclZ4WwDtKFen1ux3AGFdnfbkmi2XA/Emv3CL3oESyvqahH
t7a4gjfxuy0VgYnpFWeddQFvlSY/8Gd1/i5s71euTBykze/b4WBJZwVSgldNmiV0GMU89Tozb4XO
ikqKI2GnnWkatxoJ1uE0jpvYCSnER9GiiZdS4+/BpLxkBKHW6zY5EYkETqHbv22hYOdt8YBn61uR
qPFrsi/LJJQsxXG9JO0wNaZcdbjqoQf2vXIQz2ri2LtvSgtmevwYKqgzacF73327+1b0EtOUrB1q
Q1sInToAJ/UAdm/HAnAF38BZn37AnR/J7HjeWv+vT+pefYKj4zmllGlEG30tEdX2LNCb6UMHvJmB
7HX31/Nu0961aXSht1cKVL4K7bQgl0fhnqyQSiBGfTKUDTBnTY9a8yBhYgYiDT0J7U/EgLVL4haT
qcRfkXE++9SFo3eLdh8h8olmezy/8mKJqQrKk3gifLmX2Jt1ejMaw7sDm4+dsVz2xwJtsP9cE69m
oq7FGkOQGCnMoMSCQGCjhnn7a/Ik9lVihPxPi6ESiM14sFFpXkck7BSiI8/VqQ5ABPH7RnKW8H+Z
H7gU413QbayWzEDlo9iKd/JTA6QPQi4mkHfpSM/RRoDXL1eH4CrVo+Dt5zRLKPcjP9kozSOMPAZ0
m+5bT5tIS00WzuFrF5dpp0xOkbwtdbBO0nOMH3gzZAPDEivA8PUxCdad0iNOpYiW0LwmoJ/jSV7I
rCtJWba9UWJOPYUi4M0zWw/5LDmjVMWc6JfSF7MX7yiSBrwQiRXvnsT74LyDJCYlWZej40D4UiSt
inw/2WHVMRl5WZQ1k2jCIydLhhDCqH+cDguap8KgsKTryuMgFKl7dzSMgdueeH8LB4SW0J2uMw+q
eKfx2Fv4rQ0G1xKW7WF9NXwomlPCFPCvOhNUaWnDnxN3DEY+qHW0Avl9Ztr3xxDN92BlCznc/5c8
61TliW7NF+GZReP40MNGpY2ymSrAZZmLXIDruHC/daSXJR0o74G5TAIJgnl1OyjLxjLw+xEnxyV1
SqJnp9j4mf0VpeAPs/NwhzluvK1o85OpU80SjjMWWI16HKqw0D8gA3mQHN4WqICJFCd9VqY7v5Qx
1hKDVRqhsI/hddP8/jpoKCON1ocqLpis8vbvQwNina1MM8w6XPumBlGazo3OX4BDllIKPDNWvdrE
ttPces+n9/5HOV2J4dsoIvVHCtxnC/UBHa66pYwEuDIwVRg6qQksOBfIE+tmExfGz/ZTIBd3mCtQ
fgD5Lq0nDAYNAziGCchJTzP1ZRwhGqbnN0huXLB/G2Ny5erZqwhCUEehJLJbG3iujcrSbUiuKcbA
3vEGCXK7a42Wmfa4Zhu1+SgZc4l32jsedKJ/H6KN9ZfiD4oHJqI6Z5VeO9X7atgeYdAd7+ID1G5d
1ymbklw3rM7ZXBfz07yKiZs5ZR02caRkCOAVqoLU21ul4YQEJ8Bbl8/E27gCHe5ldc7a5tD2ihgN
xiWsdyglDJRO76rCk8b32ktV/A4b2EjTLBB4nLl2H97BMh/qEHLym+YAEnqdsVyu7f4N8GnA+2+j
+2iNNfJ77VxUYY5+Jx+DlGFidnsOzL6T9m8JXEIMFMh1iqtVYj1kwOv0hZPfDY/K7qTB0X0YsdHk
PdvLzO/qoU6we6WS/KUnZGRC03RyBZm28CFi34fhMP+LtumXwXI9bSLoEoDgHyHn1Of/enAR5z6S
aO3WdPdm4QE+rIQknf2aN8hezYBk08Z0OHz6xGEIl4x05bQsFusM5wgQTLbCNQejCX+Gbu6p6yvT
hUL+EYs92yUwyyYu6iqjPfMmv48eZNB0Zerpa4kpw8Kzw5FGWFwOiyvHnlX+bdCQDvNYN61l2YJG
0lbUmq4e7lYjqIeeyP+Bd7AIM7PiXhxXMYi2bFodg2kN+Wd4pmLp3oDfuxZoaftRBjA3pPhJN7Gh
4RfNyp/v5nL61B3X7vFoUxdxPmDCL0LQ1sHMZVvm3/iqR0HvzJ/poQ2Ln2X3akzCzvTTHU7yHHvP
tN53EnlPCjQo9L6pomVIzWp6N6IoUghfL+XJEPtvQxZ16d9EAuGNCmuWWs0DZB/eqxB4VRalgaAF
3Gr3gdSEOKlkB61sBDjwfs2vLhVOOShJ9ATVGW8i9l37kIYj/ruV40KukCFJSAkgFHfdm3LtYmLI
b8j+nEUzas/z9ZlOZqVUVZRj+nA4SmKa37/Up4sUxs0URQ5JHvUZwatJmMAEA9V2Ay9UivGWlxGu
KNxyK9ybslXZYj4RWk1AT1FBxVGxc03FeUeY2DlcN+6d0shyhrPGt0dmKvSOqbvMLm7eIxlHKF1e
Z8BW4gSlB91GP3ouhwLP/kbSwJz4/zhsK4FKjlKWlcyPeqIhcfvrp2prdIBTJj+LZQ2QWrMYGfnl
7K2+sujK3/LToTsHiarQLgVX04mlgTAL/NCm8e1FylUvlkomf5YJ33vNH7LjCyryexGaDJ3UPI5W
yWJWwpnFx/NPyZI+fQlXRm2Ok6Yr8f5RI02duXFpUtBT4c0ovm95yiwPZ0i30x0xuuk+RWbMoX+a
6E904LPfRTg3nFkK7e+6O6RqKrCFrKDPNHA86TnafQ6m2vh3p87r+E4qNipXgpm5eLBizpDyJ67e
BYVWD8kDDJh+zxVEM9POUEePUY0ar8oAzpKG0kBOj3Syiyp3lrVe2Z8yD9EaNNT3NjC2ypTzhJle
B7AWuobiaXyI7k/nB0x+KGSG5zPUv31YBBXTy4oJSqtjomxKQkZ8VNVQ0tIHiMHTDZNFDh5LRm1t
7LfUyNjTus7yzxUvALcRV0HRVmiM2Zgvg9j4t0SGdpsnDji2avxDAD8PlEQ8vkWcQ28hJQ2aRB3m
b5KTs8T3bz96/YTd1SWwLhR03UsLzJyFFpE4FZ0p97QpX8RJEhDgXG8U7K0Sef3D+0/RmVWAo34/
3NYDNdBybfLPGFYfpTQavn1UeRD0M+dAZyfRLNWX9LYFXYVs1+yZad2BWK/pHFTEzW30Ecj6ZqP3
mxTTTOXkFUJIPoYSsUH8at0bmDqSO2az3Y/PX93eCPsALqXbCHCWPw2blDFP4ONFIflblo3eg3ub
oCuJac8AXZYmBLMg7/z5KunPo0/XvSklZaSI7H/F2xq5OB1lbhNy6+7eogoiBTP835kcV/rcUTdX
bXtRCPzbQ2CzKWV+5w+d0tgC4GJyXHwsHyVHcCdptHJFAyaq9shp0Rk/lj6xDEGYY9SPnyq9Rx9K
1XD67oHK5RTKRxAXrfV1+F7/KFC0VJ85Inrr3yplLFFXomxki90SdXvxDo343+5AoHFfqMhr1jbB
co7jkZhIEvEJrDpcZD/0jgtGylSxlVMyVOMiWY1Q9NyUvgiqlL5xsHVhNkN6azye/Gekzg2cMKiJ
0zdqpq2Ape98Y+GJjUHYeLDctBuLc+rHXOnY2NCYkEEK4FuwYTXZbCacNK15dFNwRJAxbgHdUxRX
149I7hn6ilVmc0s1o9MPeS5yOqH7P0x2pxHIoQ62MWnoNlV8/T94C796zC9GISo6ms4/UDTvJjpB
QgrQPmH6oImCFjPzH7P2gc2KmN2xlWZjSCZ19vqB3Ntk4eFjVe4itFxdQVw85DtZLrAbrbzUheK8
xu3wkOOg49FYSS0Dw/thI/7clG5Xilv+F2grnVVelgL6jArV2pAzWKy2ns72gPkrvvLw78lxU3wt
B6lUnMRYXnu1AtArnJRklnJLnpc9bjDDLlM1lPOHVk1lrnsqd/zTduuQjnobyRaWE+XbChWawqAh
b/98GC3gKyQZ37QC0azr43s7gxbCzK1lSy9M9/Ls8D2AxeMQIF4GNJX7n9u5v2O4RTL1lGRrfV9l
jEdTLJFZHjt7KEZPJakLHG1vPeZzDgHZlW2CFCPb+cvCYLQMW4PC0BferqDuFpQ6/qdbm82Mnsw0
u9pbeyoyQ59aGseWvR9Bp6F845fgmMELmvtC2BLeeXxHiqI9Sek2tlW64MQfahrBt40BrLMlcWT7
gjvdpi45pMWrVQ89wV/FoeYO3NB3F6sKdusfTyG9/+BxRajWSC4LtG7Abu4F/Nl+1Xc8U+m3uve0
Zzz6T7zPhqukMq/DEVsWttx5URwMNorh4e4qNKMumh2QIGTxahAK7+JwKKXCCrJ+phosGMvvdSgl
gQFVLTZ7sfmFynaf5hNm34IsKDlShd9rwX96D6mPSX5OTOXapoQhc2AvK7idfduTJ1oUz47O20ZO
UwkJyNOV4CSOZGfVCaBs9Z8td6m/Rx6emumrwfcvlpT+c8p7lrcpO33COt/U/dUfY2YR5ZZWK9pj
CyGS3zKb84ccHje/4s/4XS7Zb4rPrQaMI5+oCmey10i6vdRSWDFSKF3a/87XbNXNvsmsU4ALWaDN
BHYCP4eB3/TWA2pXVsPTRGFmSlYnaVm7MA3e6TV/un9KH9mo0S6za4ORv0MvHlAjNEKejxT3blJV
XtU3xWubHq3wm25y6e1pELWyo3geMoNgC2RpbsXPgp3s9StCAq5c/8NxdtMoLG7PuCvpEvXawwYG
XbB+U5G7IG6/V39fdWzuIoWfAaamutlisfQjzcNwUFwN3lTk7O2H1XrsO+pxHp2Tbe9PgozrODXb
CEId+Fe77Z04yc9pQde02FsDVn6xZGf7P26kyhA7ikwJUQups3g1knUDiR2ZJk53jLFDh7qh6fA+
bU5ZxzhT1hTJuVdeXqwlMCgp25mFVNG/xPl73jsQs0l6QbXV8ZSPD1SHD+MSZwXSzLXMa11wH9bc
mAEu3V/1oKfP6uhdLpC4tOH7hpAJnwynDOpfP0VKLapDMq9R21xXgPnqvlV/NyuvWcdtwz8DaMS6
rw5trn8Nehfb/1LfyXAd++zD9Q8NeDqsRjZAEzOGRn7ssPmY0J1y6pylZzC8Lg8VRc8o2+Ezfbj1
rpiNl0RUjp9a8npdIKOcGEZBVQ3e4K0FzQE5nHOi217hqiWSp5zTQJja5rEqYtpAmkF26CfQtU7Z
PFKCYrDktBzrIEPnRtUiLBcI4reNOpV2oxEEVN/iKBcIxCLTm0aGoRZlF4jcHy6K+SV60mEmMSr8
HkwujAaBn4iy5putHEDhvTYk0++gy8sY7+/o3fvF8ObcBE4Vb593S4V4oiv3dbCX9//0kwKqx/av
nnNoqyDazf5+TmnIZaXqzPiWpP16CBg0JI1hR7hsxr7NYPEBiAQudzhpizA1voBCy38DzHmYVcw1
5GRXNkb+qRtpItOxhhIwb/xFgHHlGuiR+HZY6j2phm9+fFrw+HZv+3/pT32+MNy/RYNa6XVaR/IX
htuSQZWv+LF38nlFINfKyzwYX3aYW4mfpesfI3eOipNLvjWSdj04z/54SbrVifmD9HKvOrN2cQaw
kuf3YIS24g/Uj5bClV2/OVMtgk2UuM91M3w3AYoZsYndLsdN+JjpkW+LRbfYUmgxGJNk2GVrJaCt
MkgbPaHsK6tC1aJG74hy85qjG4hY5BvVPHFnyZs6Ru9OkwTKhjzJ9nQzSSjVAOBZgon+iPc/sKc4
2+5ETYmoyA+3k2J8tILHiQ+MBiUbz4ETtYH+qA8j5TYdMEjE8wiMGW7uG9ZWTfjFcA6mTChClhNr
uNtDKoZkC/r4CTRtepG3JUd/Kimf4UNUGTKmsqZy+ngyyESQgYMA/OxsJm3LKSK+eyN8xG7q9/X1
LVMX316zbnhLD5u1mctyiN4NWWLoYnydEFkeSsLVI4xMTU3grOKHeUKJvDZPz6YU5v20PooCfJgU
P1bBFGZJUoYAZmlRFqFKdwksEURCz1FWM/89eaw/YpDkuN8oQTqCVGTbRsT3PEgaO8L76JUAs2qB
KDx0aD1axxTtkQrulIN1XZwcLMAGTavImCNTMI0eIIErExgdLaPHLzCU4CUg12cmhSc2azD5ztnT
2x4PmUSxfEUi+RvKnT087lj1hXXS/boBCTEIprc3/TH+aqvHTJiqBqSMZl2b6dck8iIQb2D8m0ac
fgtHhJsRHd+2MDGqMqyvNTx6XoIxoOWfzOfwznLnQ6NmaH4syzJxRNAbsmGYXPCCrI+I4cPEN09a
Y9LzoRlalmq6HQzHOfi34qQfbyxV7ymhkxd+z8WDN2XEnf3kObE8J8LX63nHiAf3go8krkSxS6DS
apVpEDtkjZlcce3kiwAcXgmRyHVWL/G+LbZOjGRCQ/nmeJwedm4cEk6k+zljCisKz3bXjl0yWJVT
11cBcL0nFMLC6wDZ/DGTCXLiN/0sfFjv3252XmAn8FqNRFSmh3ppdUCYbCdie0uFzTzg90feJcGL
CICltFXACvTdym+DrG2wrtb8dN7sjHgEOO568YQD22SZl/zGiMZ6Zg1YL5D2KblVYjYYQW72ZrXU
Rug6sHcb/9XIdelJ4MCXwzl/v6MhxLfdaNLzEBIfMxYZV+F5744u0Bc2ZxuJmTGV26QKo/8w7q3y
v+RjnoTjQiZebgfRririX9O+A0eid2Pi69XfI6ADzLziRCwLEIum4l8631A8uyL8ayUiKhOfZbQ2
rFtfoa73/PaT+qsePRnG/0+Pmn6+cRFqLlVd9DJhAXxIPmrJQmTBSKWTBROU7ekoyGopWk7YVYKL
ZFQTtHeFIzlbqhHEWDWnYgvTI4DhFQ107Nwtk/oHe+y+NpYyKq/lCdn2HYudMQ6byvsaW0Ul1DLK
EWJ9Onms8NMLuu84KiCZ1t6t7QTBHgPe1W/llwDe/Q+mKISO0H5s2rmV++/JlVXNi33jpQbm8bLh
WP5HQHDRTtjQnRccOC+DoWuAUiNlT/KK+0AiWc9Tnnfp3Zl/su55D+VPVU08LTEXlmg6pok5iLdb
+33aw1OgX58Tc0AP5lXiZ9oO3U1Q97gcZHjJ6s9dmDTyHrJGZ/zqJLuMl6aRdGrqFnjK/w44GBsC
nnODnlOcWy8+ELt8F6kYnwt13/ktYOaRjrmDchUCAZoLXCfVs2PWPnq8x7CFrhr3KmGLK9uUNTe4
IbMPi7dFwvUK3UY1sQH0MyxnQ4eiKSZb7d8BTZLZBeo1GNgLYCbFwFRRaV5wRVOaFeIVHIQQLlQH
cSE7ygRlsz753cQZk24mI7BoBZ+tPOogEoEMxqR8Je+oP2e8FOU28hiAOulqiXpdjSTc4F+3aF4u
p03LKzZ4rH44Zh/l65VCjaYm6mNcDLL4WECp6Owhgr3aeKXL36UJYoUP9wgI/cnQNocc8nldifQr
omMiNhCgavUktn0g7oNUUhBtQL0dmp9o3Xv+RQwAxytkm5U/jxqvi5qntEd1FpKKBkAqJKdOH5Qs
DFXzq1FAjQc4F3FGthLFnlb5fo4OkIbR4nh+66BBA3StXilsa3Vm8QJ0J4UnK+W3MtrIkm2DGJ71
qom1RpF3C7l5ZnAm8ILKktL/i4rTQYnAAnrPly9oUr3Y1Q7CsXwTCKspm9+NhZEOmkwNCeKSTH6o
btJgNWbNLLQTOUNGw3aHpdLVhoFrh9jn3No4KWTjsPZvdyDHHwgT0IHuZcYoeBmR0HR25oIdlH2B
LDAYNiAxwsuITT48bvpF+wDLWPmG0Qb/yf8BrjL47EZMQS/7LSSmOyXRObGo+XmTqZsqpi6E2ppU
4bnWTwvDTNgjWyyHAn3HOD76M8toH/nEvkvLpqBGsBoIY86x55YuTzL4TW65ve/DeNR4PbdYEWC8
ej+04OySLvAlmRehbqz5PGlnS1UHKJcqHQKsAjnCT2rRmKsejE7eUy0pwO4jqr0xKt/Ai5KM8SdY
z8fa64tmPpPz+/o7F6cDVMrZhfbrNMwSRUnxlrl4eSZPqJqPNE75ZXBKEFDz+v52ploOyHExiZJO
XHjYiif3N/+7CCEdeqeRPxSz0NHtNNtL12RwbH+9O3Nme18KAgCR/BO60lWOGsyJA3gsoHRoHUOT
wxDyyNgyUGkWkh5WLyDlqfr+MNrkn32+L8EnOJtac/Cc6+jvXnDqyPMIyIR7feTz52zH+3sy2kjf
L9Dl/Nnr03RsuEe5YT+gxEQbLsJ2AjduU9BpKSR+TZcVrmO5FaJ+pQ7iJ63WFRADooEnt3jCnS4j
aAumQiZsVdkieLokymGxQmPKlAVhteMPuEZWkDLk3fDRqjcP3BSj/aHPXgNt+hPy3nXYOM20Q7H7
io/WWGIfiJTHGKQbBvCCBcoSfN/cGFCBh155sw+hrzw0KrsCgr5JreRM5k3fsTitS6pN1qH5HguE
OfJVYEbsFQ6M/IhmXDaIYhX1IghD8Nxdwsw7sH0vd4owAb3cLYjPJQ9go3wjBthnikf9TunHCq47
sf+1FpYzfPJqos9U1JodR4AgRF8qlVjrlk9lwZTaAR+MjbXJjc0OR1f3JrcKlLDctohMEoKSz1TV
2IU+vg+b3M/hWyd/oRRJtgKL6rhT8CFkhb89Nlg9qTclB1pg+JWEoefY2s6wQqiSs9G0zdo+lIPr
RpWt5TuFJqiy/RFF7ryBfeU8+SXRNht1YdLCcKFQC1AhsNkwejfMM0mGQbJyYyz4SVAJvSxroH/O
Kc/43CW3aNSutx/5gZRcBjqi+Ex9ExDEbgKXI9Pkkf7DqUelJevkvEDG2R3GvWOxTE+euq2gd9Fe
4YkvAIEfCeSwuzfXBoobER/CFTGcvQRoNoHCS21QAIaIaOdiqc7dtDwA7ZI0atxG/YpVQUIp4/ZN
WxuP6DMTtiy4WFaoOnsACdQjATphCVL0kjeoCT2UZuI7c/RfskDWBPcMzRzM0XIhgtupNkzO576n
aBjDyKYNLZzbSD23FiKoGtNsbh6Q+8m+KsIzUkpVOW5S6t1TPO0JGPUSv4IecsyyzTg9SCVb1vSR
I7iZIIA5MkXIE7IAKdYcSyrkYl1Mcz2dOjsjLIa1XpO/iYLkQIQZ+8ApdP15o0YDhWfbnUYCeAS6
G7fviX0lEHY0qPNmO1ZXO0ZX6BI9p2/aHV2WSxxOOfA2PR326zGnnI0VouUUb4Jv4Ri3k2bIqaT2
h1xEnglas2DqKdEuSQcn2iZUBeo2wXVdTgbG0bXwON9872QM1c7UMrOykCLa2+RgQrJVNXiZ2qJ+
R+YsJcVhpOiglLOrV0JKNRiYskq0L1+ZdSeOXxwcab+tTr5JcvF8Sj6+c9KRVXAo5+g51t9Cxxjz
n5wuSjQKYvr23J5EoOgr5g5AZhfFridJ+HVKZoTz+V0fgJINI3X8UTTDt65j32yWf77SYU0CysXh
WT8W1DAAxQh8ILHsVPldIU7v6WYkAwvhvmkOuMnRMjDaISucdRWNR1R0sF20fSQ9FgNZhb66uwH/
2it6WzBAZMLc9QDs/em2Eiz6I/+0UrytF0+1njngOrRAzclZcar2ttFPfHA7HAWtAXyVttxUzQK+
kxY8nwl6k0IlMNZqe80/YdxD/I/lEAGE2TBelgDHryZlFSslDG9PG8yKoNUQ7ou5Wwt0UghCAnHW
ZyWK4LXHtvDQj2aGsHMr7koZyY8Fx0IcbI8eP4x1rmIcTgGZ5ovm2fgNUbvQMViUJ7E6U5QPeI7i
0xzHKi8NhlQRGTC18HOlQK+m8mwvbeDtXo/Lko2qKCuNzbF22Ksi1Xsum8bgw5T7YlnltWvoNNuV
9Gvxhc6LSOhRwIeRoumQPqNSly0S9Z6dYucON4D+JO1RzejtQ9nYvX6UV2c1yPtDh92HGm6wUOuZ
MJA6BpF+RPvPTmZ1ADrzuKgXnRsPLU0cOK+SWWqoshfYd77mPYsFVUotOXHOb2ky5o6pheeM7lYV
ggclRBZN7SxEcgrJQetiBJ4SXsmmX+Vy0zEqMEYci3ZOP5Ffw3xjbkD7Ah5zAEURiB/Kz4BF/bvj
37gSsYkjYY3Tk+GjF43lFfPISJAcw26LOCoAxnTvt5L8vfmIBRZ2UWgB2aJ+5MyRlM225UxpEXEc
cX17IJ3gDR7WHBugo7+d5EcMBKo4G0K0K53TRZ+b5/t9Dei0rVz4J8gG5GXVvaMbB/begad4oc0Z
xEig4BJnZR6pLG8CGlZ4IcqqMywH3Km/XYErv98jpvnB0TjHwWjlkOXHy4E5oYYtUUbXHiASillL
R3KXcSj4IYK0uJBlscgP/0owFjKIlw1MU52gBaoJdeRj9t0he/eMgagysPjess9a0hRgA15NmdCE
EVP/PDwEC9/FvrRAs18bh+oWVXa+A56dopo15BexpOm9THMwjB+uz/h4GAMpHm7FvKmWTXxQXgxI
f+DmMquuZ1zCClENXKhXdPcIoEhW9Pg7r178nsdUMJ+EDKsQia1Vm4z1jd16FGsy6pHcT/hlqX2D
02da3Dn8sCJCCBZkxqhnN8T9nrOU1URUdg/RzFpcMulmj1PAHkhQGC2kQwq4eKjZLIbRs0/xXX0+
+TfO+6DA1b2pveFtQKEjqZmEyv5javlHJhZ2paO0ImjugDDVv8bOIV1hOFObDZVgOAsg7tfF26Wy
TExuoiK4kQ720hX7eCvF7bSWuWJo086v4RI/HWvBgIG7+p0lEjnynenff9zQu/59WMOjHyz6r/x2
dDTxL9csLubVxi/PRleduOPz2DIWtKqTsGdq/tUXY+MshGk2lEBOhdkbVrPztBg28v0lHg9WBqUV
LsMEtBTOwG2YLeGCIDAVfmRq+iGLTvyopuckCz5vvSos00o5xqJyrJWBGAFDocEASTVMnXbiEWC2
9FmXDSzqdRJeqZ3R8QqSK+AB4ftBzEYxgTyJ/YGgSoCZSOZvqP93TkUYFO6H7VsBd61FLo575O2M
sKnbrsoStW5JsY2Uhj75q38wZ5JJQ+1mRRSeEBznIhKpILfiNBr3GurYvOqksKTHq9BmJ9qXalPx
l/ELRbwmUvsqYkrRTSf+YJZFhgew8LcYCJtlpukfQoxVgRMspU39N2JeQMUGKyvFCz0nfElbrGEV
tabOJHllT2bpSNwXPMpzuWLEJLFKwXC0aJPlRAl8oqEMGTuSPMBt5RSJdz2CE8vhPgGQCywrrbqs
jpGFAPqoRZ7BVOqCHP29bBWUZ27X6UCdkWX0vZvUdnV8lmvFDFhLs7NX/GILqIrJbEhWZiYXA+YX
lW1qtD6iG9MXjoHWps+xuO41IgMEDlEbugiIwnw49cftQZp66cEiz4bX12PbLQ7Z4pJuSkS2ncbk
tXVVTh3dCekv68SWiNL+iQZQnPUstHCbNWjLMZrUHvlS9HwUsKp3+qvYl4UqNFJMuxbJN/tSrmXF
rZzxpocgPbDASHuohsZVQg1BvJcva3T2mmgLRTZaeRnWqkyJOP4P0d9gjLMtHN32iFLIMiHuDA0v
4C1M6yggBMZKwds3nf4rbzjKZwNnPb94SbGRNgyage9AXNg8DIRXXewZcXolqwgcHxMwl5gJSLh9
XZzyP4jZjnhFrOJ6LOjifTmKo9qPetQMbmGRQY/4e0/+ijlsrr7HyQR3gNRMJoJU3N+Dur7APeh1
W6J1JGVB9k5hMUgTJPx3jVDSl0BwtcQmORIniq2XkOydkeYIXBsfHyELOh88Qju/yb+NFQ9NCBr2
FPnOM8KXt2mRPR1P/xWoKL9HojyFpP1JVq1WOqtEXJ0P+w1NbMz8EDeKHzKf4YEzsPBpft3AtyaH
BQ2mpLS16uBGM9ucUHMNn6Dc5W6UN3ZW3eCpS6N6Sfn2XKFM7Js8LkTssXmGDi/05QKbj/gt+8Dr
d6uuLka/5mcepAD09QRaYlSIJ25gfnuuTfnyGrNyvYfulEQRUuMI4M7fnSFh8KR/jaNFxuiGvSXe
ulcpl9mIR14ItaxnlvCOz2Kvl3bliyhCkqFaUqR0xIo++KnmGU7J3SkaIj/K2Rkk5k15zdpgYaMC
E61FElR4byEfYv3IilTTamUrXS5bvKZjGQdrgJpSgSi+73uBRrL65pNzbvwu0gCLp+vLt5ATVED/
iNVUw2DCPdR2AqpDCyMG6P1b/HHul8xjmIjfhwgQeUEWYgR8SEe6VSkz+oMkM1b+ZyzRhZkAuis/
ED6pevSWMjJGtw+SYDy/fOZiKziKKB4cARZfa+LSY0A6hayr/9wYVY3r+/j6uJanw76qotNMS5Fs
R6Zo+CSG+IH4BJiGu/NatK+BqtJ4TSg31FQtoyN7okqkob/mZt0oW1GQVv8JDXaPdca9D0NU7AOR
D/whqeFOsdu53Fi0daCPxkYI30693SeyYU7cIIEMTqpU+OhJ/EtAxY+kwXpNSkUes39gxfXuECrk
je6gPIGuwVkzEBcSOkf2d55VLTVTXhhwjpO9QDRHj3AlhQY/0eD/Tez9G4GJaHYuAMDs9nefWceK
bWVVXcYPm+1pZu9Hpj59zy0/cBVkxOf4MV9spDvnaSLaWbByeZQS7Ro8WPlyLgLCHp4gdvCqzzcO
jzVa6ZOLgV/dVrFBFUeRudkuTnhTx1pAsfhiyYjmoLFyhVnOMo9GkmpbQ4zgyZNGYLDgh8/6g6kL
8bIPVtiMYwi3FfEjZdu5q8qwXvKj85Xo/OJUmUcXreBy8EOz70jE+8QlE4u8MpwHlOR8PMn6lzIK
YHhp5AhiBIb7M9hcmEai+tD62GXJVDXm0vZbpPdii8Q5BLGYJntfpd328fsVwgmFbqXkRJrgYF23
i2TMK1G9D+3dBWSF8NwIovSOx9nVUUapMxRP6GSFT8np6ahyMhamiYVVavY0nc9MN0lczQaGOwYe
IJBCEHBGzSHG5CVBHJA6k/ZVIz3TLtaDM/PvUqbsMnGJuoHaDb3eWSIKJzAwspiINOcKG8pCtanb
/GdOO0yrea2/pIeHwcKYd+wAk2WBarffczV/de1t/JHRymrTmB9JzrRojvn1o9paZFRbaXyrZ+Rh
GS3SRNky0ryvmVHyREKnMS5syRSRWWZhVEtj+A/jsO6aJVVk5X20LFCY5TRryEOPNTz4DgZd5VaE
i3FW/VrucWGnm4ZEW9apLxcICLDNBXOq72wi2rEI9Qo5K+31GcGDzrCFdDho2qpzYDtUMg8SNsr9
KZeiTf9ZYeAjzEdm6fy9CMB1CcaNu0yOmySQoV4tzNC9w8k9HZgBEyiHz7QXPFoaACKfVfxe8RFd
xP1kwVfJFixk+pd46IQaxq1g63ONdRsZG2nR7FcVRHaJE0nsRfEX/JZ9AzeSEQoLlhA/PPbeeBx1
do7WrDI8TZnV0+6sBqxBXzG+32bSHvduUO27t99TrYkEamAzc0cIn2vXikdVU2KLuqaN/SGX9vt5
lm/IV0kgBLGkjGOizDGwW/GfsUz+D3XMB42zFM4kBCHKiuy9zn5dGO0bsFaOM9+wzcmwf/h6E3hg
Xm/bquuHwBXh6PI8x7lM7UeP1+8bg9Ri3n1yhhJnwqYgj/XAtVjcdIfIEFVxw+1IQoAoOSvBNHPD
Q0lrr6+k7xrfmBOuCP1zqJ/iwJC9mswqKMWMy3sVI9NpkdjEBvs5KcyNELcXr8XdBjg9AkIp5BNB
yTRRLU0OkKs4CnvxwQv2OIvTvk533loMZYWEEG14ctec2FME2BFSLLC6vSpmm57sd3c5Bc87OhGH
DTmOLO0bPMXfQtZGWiKAhotnZPgIJl6G5HZWdpD+bF6F7U8B6Ci23RtVj/tzCs9/c3vyzzfSn3Rj
Ae+ZmRDS/YpbwlRy2pPI84XFiGnZ6N/vZ3MkbrFw/dUduQlAoTkbDiLGQBHphOOYnfBr6kPvtrIN
XM3iZjh+joX3szLYze8vRKmro/8I2uAZILyh1f5RONL44pkCbVhHlRGXLp6lvOZuEPcHh+Oqh1UQ
OsxnxEe1B+aAPI3EvaUvb1bdlLgTzy1LrdPoTVNhfhsNZ5cEVZk/l6PLNB7zxDZpzczAXGoJBMrI
f3tVSVtp6GbgumcXUluwXhx2mg7U56ApkaGqm9JTgfyRSfSOB7+z9k3rVp4CDzD4MYAoMKlmnlPQ
pasdG1zni1NyOnPALKyfCT1wGsQVCZdp6mvHS+huENUlTgDimSTjF6PFTpDAsOE+GN9j/aieGLAO
DZ5Y0MHstL4y7d/ThArrkSsa5ug5BGgTnxlj0IdNRC768cEQzx3rqs49aQ36ufAXucHV9bjxvusy
ouWtiBNLmAj1+Yfx7gcOKONZsah1R1VsObEjkZL9tEPI7ONUqRbYhB1HMdUEL3Nxim4jSTpf0cOs
AD2ysreWpfCiwUOtG6ecETVxLTwuGbY1wJirJKUybsQQ4rGhq4eMP9qq77Oq1pD+9yZl45CVX9D7
CfCozG+jevbFflYnzGZU2W+bG/MQ4NxDX0R/3s53WhpjBFDXVQvp7b1ODiUauv/Hg0kTdDG3Crga
DcY9jJuU8djY4C75EKKZZMRJbHlf43IcL7LrqsKpKHKeKHvE0em4fV2P48/MMyW4BBX3+x31/waA
tNO2xExU5ejWSLVS/tJmRQDYHP4bPJn25DDNfJ4Op7RTK0ymh9Be7/JoLWu00GYgFl+PZpfgPxLZ
sniO25igA/5ymH8pwcv6kG0bq+8h9bSueawgNaXiCcEX8We0fyjipEdS713OJlBPYKf6QCChK/OT
H+5txf/aXXEdyf2V+D9sjiBRpE7q2WLq8Y49XgSbXnpcIiQYtSI6mDdcZrbf2/7pvGCmsmalSn0u
14U3R23SpeWJxG5W3KhEQwsbZPutJQ0+IwovUC28fHobK4dtc/i4lk5FdcOHTQyE6KJ2I29pDSsB
UteJHkHClpsUso+DbvGFE8KFPXuLrHGhdzv0WBczfry1aO6Tjz8P3uBZ5+3C4mV17oRciwiT6yBx
2LZoAMkgFB9XfpagNSpSiGF1olk+SVly8OMMUXyzDx9DIbzpLOek4we3Zd5ivcyKDD6mV1gsf8zA
VEXRVBvXXVtfeRuPcnw/bCuz+LkKxJNv5q94ek3J2SAdVQfkasLsLhvYLs1QFPyhRUWZcEwfYSbN
dJhfvCZ9DDczm0D55RIF7UOoLheF0BHw+RHIVJrx0rDfTL1Yz4oy/2V1wobp8Cuazp+Kqc0zS0Yv
nsggn0gz91E8LGLceLP3IiGGpu0/vJZRjI4OjjZZSuCdXM2cuMEIfzbIFxCxgydX5a3CkGcrjOzN
A3yJkg0fPjLqth+ZZGnms8oYxhSnbHsQqhDc4M21yhNxN1JJgSSI4dALc/NxTgrpFH6y5DChEadC
QkWc32nN3meY+Fb4S59jcfQqkw1kPq8TCLtZHvwCCeLcSIr2nuV2D7XQBq714vlYIaNPQ/SWwZLW
OYGHtJ8yRIM+OQyrnZ+WtyNkkORsKGOIfNrPTU9qpCpX24qEuDhJsiUq+6ToA2PgUiP2766JVG3Y
e7bg/G7b8kdegm7+wyZmG9vxZTDuh2q0AhugaLSEwZtV/LvjIjVEqv4ksJLq6lw35B5b9QhGLwJo
PrMMpX2lL87/6IG3KJlIBOlxip2GiutAxjZCBAcoNrzvJZPAjbvkI/e3NH+SCff8zVjGmA+FCiMO
7eXmqLREHSIytQ9DI/XTwQn8VK3bXRQgsPZRf7H21DD2rJ9UrHYs3CyxQUciYHQ+Mlrm441iKd4O
pojkR3h+ff6QUqZwEvbGeitQLEVoSG+3OUbSRJtU/Qb4RDE+o7eiVQd60O+a6FF4bWIemGG8LLku
hzLy9ARPjRQeXpDC+4vdZ7aL6oR/y0fthVmmvHOSYMXX2wPZJREx50I1rcxiXJI28MEn2D1K0h5z
pgJK0C8+6oQ+YphWpfMf1k2Sj8B0mWEoLpX8L03kC48dZ3jWQwFKhALT3ySNT4z6tl+0ElADYhUQ
Oeya4Nz+I9kbitT7bhd/Dwlh5ZDGd+LRVCCjuRAIWjSMEB7pU9p0VRVaVda9m3vHtYZjvRpq4Dcq
moOT4zl+oTbXjQ794tt0TMua2mHR4O6TkYJCOUi1KrB/QF/BqeRiX9O0yyk9i0SPoXnE9B96DBMQ
yX+oLxOc5YpGlnuz6+L937d9MLW/KAX/PNS0neCk6JOMWNLuiU1xD8u5bacWVG3gWMYvHEL4XIIm
DH8294ET3kpPNvnFn/IhmdtKt1fqsB0HuvGpBPY32A2Ddc6NgC/78wfTEg/ylGp52Ox9Aa/BVdsP
pHuqBp7WvyicZzai3O7XfKrkRDJZoqrhtzD56Vh04B/09u3U1JrS3TA3RTRZ74fXJKyUlRDKeoa/
GCfWvHMhAQ+bAy2I/rKrMrqLke0qlwrxvbszlKoe6JrzmtpQjXbcycpo1mEDn+c3VUBn9diDYcUH
bCQFGU/gIHU4Jx6mKKZ0Qq/NUU5siaklagYSp955c40nM+SLRoAN7Klp1Z/+kmNjjztJ0WV+b65u
UNminvnXd7byKLuTTt5yFfrodZeomaIEW58A1uds4aOQ3fKQpFRrEP2lXZuaxc3LZ0JKqLyH83dx
JXb8oeFirYxsLcsXr6KBm3mKgRdpxUk6Fz7AQDzI1Xcl6ccU2TteJesx5z2crF8ULn0nq/DNISYS
kPGPLPmWh8r7jGgaLczrDDgpevhC1Pq0fAeG4wewIX+8BdiDgZk+kCahnIy1Tvk0L+ZaOjuwe6pD
3DEyaYBKo4t3xluzB8OwjhlAJJ0/gQPAmHSW58bIGCf2V6ks5zgfnEsWC/Rhgg25qHy32qFyF4or
kp9WDNpKIiGyk+mTf9cQnkkh3WlfbjTZFK3rSwRzFJtmNa1MyCv8kvw1ZYdz95ehefl53hrfsKPr
GfDhx6Uyppwib6Vd1YgZfLobIS9/BVgbnOWISH5blVkYimMbBMSq9kSbku0iveBICFuNGzAbj9JT
ojqxt0zQNz/woMnGbuqSfV2U6EFwcwWmBzVK134IFigy/WyPhf2Ms9Re4pgefzzJODmq9yf5dUee
cJMV7DnMZAwuj2tz+TVzPwzwRsRAIKPWB206FUg5o34F9BzSaXkTZflFRHZxYGBA5jwg46rFrQlB
LgXcKL9PLCczKv/YR4Q6qJ1LxmSQ8JHwVW3KgOdsLl6xdCa8wJHJrrtLR/BJvcKztqcPjTgLs/Ww
urZaCDJxgGuGMxGOWE2aaaBUCxIlG3pQxRq8lyqbq+2vCRYTJIrouRLCATJcdwky7tEWJfMrwjok
xQE9ku2WAqaeRw4JQHCdTdzUfaTCkL18s59kjUZSyADPXPZl/C2mnuW1VBi/6Y5Uwg52mLh6MZN5
WCOhVF3Nvv02sZGrdFwF0HMgiCSPkrNj/7P6v0P2XxY1NoFuypMYe5Iv3rDvpGwNlzqfIPqOyLEs
K8/RtK1EEyWJoSmVdf3HrKmbwH/yIf5oY2d8ANmjUzqzslh3JsCWFeIFMhWfpIFy7kQtuQ7G5erO
Jfr0HeR/k+Kr4EhJ4fVX0bjP70gXl+VStdYZmLlzYv92BQAmvs+GWIpt1178tuTYJQOmhix4lfPB
kqP2hWx+i7muUhfY8IrOiDRcpfisG+PpWMRkbxDThPp26tKQ6zunZBA8VNh9yLwX6p/nfxkFf2NM
Kp+pPgvnWhlA01oZU0y11i2TTn0wdLY9B9v53nho02Kxer7eqrnC+ZTOTW0bCAdKXPpB6SxMAtnb
c4kIF6ffxkVkUoiNejJwcMt5FhBNLPeAL/1agUL+pDOY6oakWQG+jGN20AISa0YqBqoxLkkN5xEJ
pmnOx67exjDm1iQBoTtU1gfZjTAGDk6yvUSGc9nOifQ2cSdNQUAAs2fswGfXZfAHl8SAVFxogl23
TbCt0u91yB7iaA6d6exULQmnU3aJBcVpYI47iaD0lDmxedrZ7NO+UM4bnLBzgWHY2s0HoAmZFI7k
qFAhVmo8xNva+9Qt0NQVEzKOnO/Dne0wkpQ7FFtL4QcbUGbK7V8DFFRQJnua95iQd25sBtk6LMPa
9JLLw4VswYScr2H5+JIIcPrSYrs0MFapnKWJs53av3gqfnV2Vpvhw3zLt/1Cp/GpIYgpbjptYQLQ
zrg9btGHFQsOpT2xeRZICOnnvZZrh8DXhGubRknrJtNOAHkhcs+yvNoMAUqJmrzmjd/M1lxOQX0K
maB595dfoRIMC1f2ALwsZL3HQtEpOmtq1Qv2iwxtatnFoDaM6hCC52IyTYJAyAt9Sv4S+cENKZ81
MMvrBPFHtYCAU1yyAyp8Jcip5NIYt/WgSddx2e1WSGWj6FwZyhx4rD1LVLcAjJ2dUF5/oRSb+NGR
WZJ7BcM1DqSY60hMtn1exRotP/Akptbg0P8I0y7r2k3mGxgD7IfQzvRpDnbCgq9g/4uCBIOglpW9
kRIL20/+524asUYeUTWE0qpuXaIkMvQ0qmNK5BboFMfUKrUfVkDYgLCFRSlPDctejLMiO1tk89gL
ibmVqj9ThNT5rbOruz5r0BYR3R2QSOklb8k5/1JRmGIBqIiO/6vPBgL6u0BwLJSEoH22JljAhiCy
RFYzWsjZdslPogr32/5N3vmVS7B+jMJXQUPxOSpGCIWopp36arRBabfZO2hsRXgjxze6udPd0cXD
JwepE7OeXie3jGJIXoeIP9/XLxCGgbIpthWV4IGxxYQ1KcKJNrohTDMvQVR6G1rWZrSrbgMGox17
RN16ywili3KUAOR/vESQRHKAUr2484ENYcICUmEz8OF2g5FtMkgPRCi1wd6LqizT5sPLOQCftlcM
g7JoAlcIUb/PSPTq0bZZGRuKGrlVRVugtrRLVq4bUmhw4dYFBkH140Jkg668Wy/jretXgT4U20G9
uYCRNBOK5P+UaNPoTWvt3UdqssdOcVV1OzGEOtgOQAcbozfa+y2xIugV6x0sW/aAE8T8vCNGAKNd
vlQ3IPW7FkTwy2xQZZ63CvlbMkNxBj7u2L28/4WZSjt8jFEFEZL+aVnso2IMKUCAyjzg808cIVQu
WmuslIDcQFi0oEtZGPk1D89rocobbZtRTts8K7ctcyAoTdYHyRBzpLcyf8enkPldNwv8p8vG/Q7C
hVXTIgYf7RfvRNZZzfAhe+kyK4Hp+W+RJwZdAleHiFTSJsVyCaEjFC5V4yPKUCDCNUdgyFPQA+va
pE3GTGMHzK6Zjfjfg+e0/2jN8OUTIbzsgTdM0DjPemPs4QE/vEYbpKCYAjlWcLxm2a+euEMiP6tv
VQ+aP+xGehwGi8EWfkkO8uF7zFZhj9q9lnbCS4k051xcFzFXOT6u4qKJyoYzZlDKaaL8QVwi6tDT
sG4goQOhFLIl28wiVXDtr7IL1boxWbcoEFN6IR5bp2+bEAk/qU+Udn6ALa2M7K/rhqxWtJIz2YLr
7YppjIlQEqQjNUuCWVNlKNvwDa18GuM3E8ForIXF+Ya3rgQqr+NZW/4inwjPwd6zH71Zt9Um6zDU
JijhZRH61lSOpB1z9KKSnf13GQh3F2rIO/WBeIH/N3ZsDdJ0CnRsmgRb7gMZdMvQJ8JiYNT3yJVQ
fXk0dlwp0dYlqUBuYJnlsT5rHgYGFDFGy9QvvGJRe+QW37Nf2YfonEgHD0XG4aOQjmYSjgdF6EZI
lsSbjpsCeV0ev8t+QHaLR2PPTn4nY5i7eHai2Covcrdgee6hWN5m9qK1mNbMyA6aJJbwzLM/uVp9
S5xKFEKHLYQs+yt01dxxJ//ywgMwTjiOxyy/GzGVo1yBSEq0EpOzulxBGpiJz6FPBE0Vh51P6Qfe
lU6gXUCRjspOOZOkT/iWNeGy1ff7BOy5XIl7GWT+dcbDat8La//qDACPeHCnRXptDtnN0oxmSasp
6/E/7YTtxz+rwlsYq+OiAFYuDNBPMQfCRkiVLtYnojodsuM8eMEP9LM1prkzYP7/xUwF3NMIhTM2
qM7bZZEJ6XwdaYUUZTclHUVcM0DR8iRsRDJTLFJF8rZWMBg7YHydzjGHMZ5+8/fvxMt0WIU1N2O+
qAxyZHjhOysO6fDBDYQCasH273uEDKdtJVtbhWTdeYP/p2qweklJmxvIuYo0XYFu5uHbvzZmd4Ey
KRNI0wptun5VYcVelIK/EQMHW0j+t4oDhfeUFuiu/U2VWvm8JqB5C6Z5GEo1i04osZghWcglXe+I
9aaHg9pJFxuOAzyJ2e8pF/8px/pzDp53UEMsVv4I2GeihJH2n3adsZhkJTwdJAz0snbQuSB85sc2
jYefU5Wym0aRWpCX60Q1zqRi9cyBzoV1/woEnPQCcDN34GfWQwB3PNTMLtbINRFyFkxF5FsS8+s6
urhIDoJYp1oiv/bGj/4I5bNBgjDp4+kw0HcGlVhRAuMBwHL3tawQSWQxp3ijDmXqZSuo46ukXWgY
B7hlcLsg6hVHP6dv5HQCJaiKSra5uvABnocgQr85mRu01RWlcB2WA0w28mt3v2pYcaN580AnBPY6
9siTGcWzx0OaSTRrtngQfu639fgDmlNPDH2xtfvst/wNC6bqolZuuRPsVHmFFmXGFgvQu4KLMKcI
zAH9dVvURTLG1a19tusBG98kaATqyftZcij6Vo8Y6Lra0QmlGkplhICZW0BWjFHS+j133j402hnH
K8RhzUKZmRCwBG7HhYdtEBGXq09Ggc0SArJTJkG6Y9sSI+uKuUrgxqkzDfMfsh8BsD2WUCJNM/r5
/acLDykfVHE0gA9Qs+3XSncr3pPzm2jXZjgcJst+7CXtqbS33JitRrDD99yV+4p4ya5UihAQJNtH
c987+2wlGpGVuAZ01UjWFxN+4xDuW6BFOJTwpBmwHZJ1qz1BMaKX+7vvU0bs0pZiDyjThmG/Rbik
Vn+BrmqqfpJU1lJ4Ne63ushQuGjVR4RgyTPE53+q24aGfSDNypRZ72mnVIj5/JrNkcuGmSzRY6Ut
krDbxa2HTAfbWu3srznPJ0hn4MezIyaP0lz4GyVqAerTt2UrAE3OUFvpZD5kAfszHrB0ugj1BLGi
SbLeFEMK3PmC8vT2RUVwIVCc6eYUFOotesuBLDazwo1EE/zKJkgwJE5CL4HUnY8doAJ7G638DxWk
Ex+JKce5JWGsCMC+N1fLEOoGYEtxJIwr+k0GCYSuAoYYwh4scT5cnluCmyy0GGY2kmMKX1PkiHaH
wsbA9bvPo4DxxXFO9KpP08Eclek6/flEv9Yo+nbpJPMsGUrNSecm3WeMmhXdr7Pek0Z+NDmgIWHi
6Rk8JNGAFN3yKI9dZq4XEPhY1AOIgfM/b5JU0nb/CTkE+Elbmged8nQPbHwFGstTV+eAtiv1ot0x
RLR3Kh12W/oFktppEmUnNfeN4AU16ewDeibUUO/IDs6055ehkfs0EI6DZAMS/LbqMoEbhyJmPS/N
NE6/qC30WMF9Xx88i8CYVnPYl9f/XjnQJc8sJxc40WgriH2RgVgHduYTsKT3LnXpM9kv5oAnv+Dq
dQRmapZh2Iysc3JZ84Uko83bkPwojIyS5fUzGxmVjkYmB7gzStcdymhcYJ/lGcSyOovktTuxW28E
shhga4XRe7FHlqy4O7B98gqtHLJ+lrsD49xsQIXy4VhaVPKDr9DQiaDXAt5Jyfc5w25IaG41qxmm
AfhpwEvBEZFduDF4qC7B+MIwgCt1rfoxXlsUvvlJNGOI2hHdStuw8rI95rBh/B4Z7l/4ciehp9GK
hXGi9f0eWiYHVg/Sg/B8GxXBtREiwWfDC8gQShuydz1tRElnNR4oz9jorUf8Uvb5IND4WPwk7tI/
6CLsz2PzzL9FrqlgjI8xahJjALgcQwpCysd4o+z5ClZnaUMsO5NIYBV97g3GCk/JSjPBbEaMyk0K
B5Bpd07lGoRVfDmWkDcqXTc2WbvJyttj1Zufa1K6Ez/3fO7LUjkraajcHPneVvyiPZeBj9y/8Iwi
zWLq6zfBTljohpk26VhAqMkmSzWIt/Wkl1qh7D9fW38ptnZvzr1o6nxS9S6Jc4/FIfEQ6+MiCI8s
0YSRCl/ck6VuLTqhrOZpVv/dBtAtamLrhTNm2dcYw+a8Fl8VwQyJXke/1vlE1d4tJ+ut1wOdtECJ
UpiigEAMCC/nN3AGZ7uc1M2uSxHut0/RAjcwLKz80R9QHVqV3dkbD/Gjc0whvKC/n8+a6NqFu5rm
HbbcJ3a5Ztpp2SQBdZEO82KBCSNh8YRMrXkgAZm8B32Y/6cIxJt35hiY67qisGX04fP1iF0BowJg
ymTOagVnBP7kuIX7XPMvmlPnd5kEh1REbwqG7gHnIMYkAsOF9mKTm+fNpXJCuAF5p7F2XGL1YpHR
RZdIgG5USrxqbT13Fm4LtPNE/IIOmpLyeIYMCICLS09bubQpHA896Axo9WPimKAOXaKJ2UPSGkhk
TM5Ve1ACnhJQAeGARAhtW1gFKAAtK/2v1xRa3vXh52tKRk3g5oAgFpj13+SyxUF/EYZkuzt/LI8I
ZI3L3p9RhDKDgfUMF2xHz3n7zoq31gsZgdcFvDfZ1v+nw0Y9Gy+eNVxy/K3SB/B/En4TdJUbct8r
NAlZxCoseuwx2dkfvTgwtAnvqLuuLk57EdTUqoTCneUr/uNGtcwVMeozdT5w1RnIjhRoxCoPLLNj
OOaRDUeULsWp4NaBL1hm3/q8LpEz48GKTW2m7XVwamzeUtqal2qqmzGMwwEby4dlPYindTONE5Ic
tQjKwyJXIY75kS46pVVR06vYm1uNT2fNMCe96EPGTlrZFy5HyjrOeoDFbUIRFz8px59VT7K+rtAb
tYW5ecQW2oimvaPZF5YNS/r2i4yTHIT8D13RtsBzPK1HvUqcGVv6xGH6Y8gc4x1JsLUmGTAzPN71
fxmos2dFGSOHKACUsSW01Oa25qXxIWrdJZhXqgCXLEms1lT0xOD2Auba+/Gb4n4jCT1UKSOfpgOm
Jig0g3ElSm28cihojf2fT3Qrt/vm5JU7ojosBFDE3RHbbnam9piMR6ZU6b2oDkRJzA7She2xQcr6
pdEell3XquF8JCCBZHo2jNwQWShNJiIYBy3jQkTOfMncc6+TaahJAanPC3R9vIsl9cQGD0544Mlw
gBwCgUkLogjgD2hO5LslP9yjNO+37DgT9lH+/xsbyo6ahwo3gxGARTkw74QFkLzxou1moAmxwUHs
Y60w6rHMqRxqkOKIdkwLiAV5SZEKIoiMs9JExXZVfUo8VRnilNjGtE319Q4CcRW0z13hu8zBOSUt
YtExPdFtekgPfc/f0FhpHSIGN9+J0d1XN44gwkSi7JqDVvV5iY7nARoMLdiUYcENbYS4z6Wan8At
S0wtVJXSEwnPDz4wmoaKguRj0dxYISCEcXgosYBlXxGHMUap6g2FSuuYahmC0KImjM0bFnNMapv0
hYXaqMxPwYT7HnT268L2bhgT/UQ/hIdzjYL5grpsu+zA6v8byh3Mp8EUHVFBX6a+CIc1neYHUKex
m+YJEY5PMkuXU42IvUccUUMKY2MJDW0PhVa+49b4KCkp4igGYFzhTFcIWtqrRFm8HANThP8wQlsX
Xroith9KRlrafCFLhpCTLD/RvF8ciV9HfU3hhJTcW/weYXIa/PnkK8SmY1I5N8IlKO/a6obMh+oq
GlGQxtEewWMIER7JJhAREn2ndJ+4zzHhYUHNKLztku3WWLNm17oqWgcRb10W1GnM3Ko6rn6coE3f
NfgNLXqXkl6C6ZBgcEhY7+8b18wIxQQwdLIL3604rmlbQBp2e3RWRNJrYeeqbL3OLq6z1pAnBvmG
hlu1EECJzEj/pOwpG14qOII0bVGRt6JkNHMITWSwwcnkVBoItAiS64aUdrbzWzq60zl8OCkkjAzr
BAS+MccT/LleLrDCpetoejcUOe+FpEFdpgZLUpF9AjOGz0VI+kNlr9BWuR6Hc1gBVbD8T+KsGF4b
fCFopnwUJ9jTtDFDLtXLRXec6MB8yLazo2cZtu9VSccnOJEuuO95t+ELILIR+dO95EhbeFJfQTwB
SfcocN19/NqJnMJ5ki05qx6CxetFkuozI6rBWrbr+3OmVmPMSoVd4Yw5VmNth5lcSO6dMCyfeRCz
DBH1wp9y2PSpdpk1OW8369jguiwesIoh25xpIj2Fz2bQSrRapUrwgVF0qx5+HlaipajeJORn8wTn
qVbniCeXb9z9dVI4BV9he9M86zQIOuhVkBOcUz6K+ne5XakIpMbYqkMXe2VbzWd8fJTxnFRtvjaB
jAdyhlyy8Aao7N09MqDgiPkxUnEHioZXkAyc0MjmZxu4U8EETDHRXFD/ni2+dGv6oXDWJXpVfBwZ
5r1cd4RSjykbsaq2hsuyMSHz5oxrvGberzqO0uTgTuaouizHkPMcGiiQB2/vMHbTmLkoiLCzrgRf
UAW6pKNhwX1l8hyJFRekrP3yTK1zFjFyigcrwDBaYB4uQOxzNyFyeBtO7LP+iso2oQJibK2JGd1c
y4AZEmA3GjQB13RLt53LGFXh+xpk7oAiIfkZauCu4ZpcobmZvd+bVVn2S4IbsVO7tuAZxjC7Q4Zo
wiX9dPvFzydPqt//mI61/H8mdRy3oHBed9ZIXZWSbHou94H/u2i0WvUmIMB1StFA62TXMxQdjlVm
P3idZD54igx/QLyOUSlFyYgZpFAgU6kqDtVukjoBCJDE/RIQkyDnLGSZ7H3vqlzip8tFfnjFTuHG
qApqcry287f1x42yDIITV9KxodS7sanGBcXcbUC1KtEO399zzmr2dxvjxiWWRmfjYTpokyY0T7wT
JGiYMPikX2vYpGxpv1w1oKeegke4JcIM1PrgTQw5Ms6aEUs1oI/dJVc2/BL1MmVr79rHNHpQDAhB
dI99ejbqiS4zrys5WxSTEjCOtA3GZJajDsOdvUMepQMULST31of5imKU8ZF5z+AUVLQXpnC6hofj
lMPj8mhqw6nxSknJzIS397XxYNvnCvT16DcFTiJdEHApRVY7+o76TS8tUm+EKxvKBYYHQ+A9Evf8
7WiLmq010ucvkLbvYrwBrY5l+ProOr0WeaaEyQr/SFY/qCZw1EZc/tGQcMoZyexbtpl7Um+AQccf
duBV9DgIf4vRa0EJLYp2JubnYU6PbaQ6fUIUv6B48QTw0Os81/OQWLWYAGe/M37vmsT+7nklEDH+
gYCr+kgE/wBsCUpHWssG0k50P/s/me3Q9hlFZBpfCHhl0D2bu6PdQ6YHjhwLQrf2vRLCdGLx2Z54
sNfxrJTGTBsLo2b3yYBrgoGoWOqAWIZilh9E7vekcUVMl29EGHaXfQIv8Ho+8qepaIITJTqxIal7
7IwBXKwmCMrCcuvskGOP02Hob9S1sk4Mgnk0P6cImRt6JR3m2728vt3I2jUQ+hW3sfjD2YjaicUM
rce01YOU9SpTSv44mwUBNZRnyMmh2Hqf2rZMjt2MnBRWaiA9k+Dz7wblI1P0TqLQdMXSvrC52wvE
hCvz1YwvIpOBXSr6++QCqLjp5+b3fHPLizK4deksDvjG0GZT1sNAgSaQHrtAD+ovvzW5qgpdT+dZ
GxGd8L0TDvHWu7NqCOCXeKvwQaLnvxb7EvKqmprklxZcK/79UMsZ7C2ykllmNcdVFaWQVqKOzc6V
6uFB/5u+LoEvsOd5hWCoH10/+e7UDVFbq8qaSiL8CQsodugwgXRRFduxrei+UGByjeyml0JNu7DP
cFso6Ph8d9t58HswQPc/6kBHrq7ATH/FQlqiKeIPoxj6hv/7k04OvwSv1AanTiADw6OEf7B9tmUO
WIVHz6Ehaeu3xsZ5ELeAr9VrUEGTVJPFFK+/tY3OGUIkr9u/IMUDDY4efctHCA6jTJfmpL4YPuM/
Os502pCCKReCyul99cH5Ib+YX+uajrJ4aTDCnsOaKieKcuNuKC0w4fUu+XCPGTR3UhstLtn2AO1C
Y6ugmV7BgkixzHHvWS7KGAn9FWEmJFqkTWcoGLB66WXV7/T5QH9wxxn8zTcsz7cdqqdAcHbjqW//
vn4I3CmmjsiUcrp5Yhzh841XbIrKzQKeqYsbLLI/gXZ/rzImV+7hAp9HICrVZEE5jedHQT5FGqEr
Gevu5B2WvVaWrmgzLkuf4lsiZAWB5OyxiC73UmFr1LKCkJCqGL44bhJ1339M7KlfNQz5xxNf7x5r
mbWp/q4cG/9vI4OFmLjSgx1DJyUBgfQE2LCETvcXwE7kl4V6itIuPj/zfw/dIRr8cKijGQ31MKVL
nzosftv6aQ7m6Zksyu+AUIgM8S5pAFynSnmDbXTPSKPO4ReJllAREiwGMH9ldbr/U+IRBRTpn5q3
w9zFRTnt4NpA75g3sb8ehTp4QWmpAnVlCpjhv6irGNFA5H+XUu/2fmZ1cBM4hzN0SQ/k7ikZ1Tlf
WJic6FcedpukDd40Ug5Xs8QdV8RZ/1ebxo3urmvT/wpwcm6oXIeWC0gzwCyHSipOuS2tB+vZcj70
qObWtVLW2PnAYLjyYK3NmdWZpd8WKtZySYFCY2tjyTuuPYRV+mPjy/cB4S8XhlU5WoDqHn1rKXwb
0cfJVdFAhTVmUlHnBVO2UNAdVX4pZm1TJED6MaVPLggqRAp2/tE0AzQfpDDbVEfKzTI9JL/3dy41
I5dQ1t/nvpaKGSnHbQx2GWoPttROAjcl1Qe7zUStVBvlbsqFNUIoaYuhgdEmy9fzGIR83XqD3f1W
zOxLIRgvVT1YEpNlO0EdYFAaxK4Z7fyKYX2TQHpAVj7iDVmWcxnUg5OA3xKUdzeSaumC2UNyOiWj
7viYQELQc3GcnYTiTk84U4IiMXw1alDbFPTk+izCcWVzNVn/1SUQPU+bMAgmBPFSweexbWdrLOHT
azYbwLoAicB8TgPaI/H7jtUOPugw1q0dRGK5OzMVfgJv/q+AT8Wti9tpTxCMIkU/s6IlYAxvQJhh
5lWDFAMLE65KGfW561nVyb2CZLC8bkQuFmHwVidN4lrTyj2g7mVCEXHtGp583SGmCzeSjop3Tjrp
sHKQzGMagLpOMJphfsAWTH802/PPLyCrhyNvYZ+fuJsYEIzJ7sfoJkJdxRaiJyJf3U7A5BqXbFSu
kVgdMMzHLgQlTrmlnZFl4kSQiYt65uoWGRip1ICpthxFEecttisEpEZFqP430IGbGV8nrOCWPqCy
Jgs+qwP6+YZ2r37PF3kZdTioCvqt7M50RoTDrLG/HPa5Q2XGZNlKhMpzUknXkpFhAMjLwJhYMsyq
CeV5/u+MIJC/OBu35ox6l1hdFuuh0KnCyKSjp5tTHS+fHqTL1LLHU+wxW26a0V/Co5sTUiNx7jyy
jT/Lk6d1n06zr57MptjJUcNGbX0IFhWCRh9JmO647XLLNmkTITUrANGziDWAdQ1J5j6QHgiFzIEa
kHLFWWwtzmSyqaOpYvFL1KXCGUE2yrH+683FzIiSz5pSHR5XfP2byzVTrpOatc8hh2cJHTHXsRNJ
kkySqJuXd8oGIuXf4qOiWMYudjfmGxTrHUft8QpxZKc8SRIXrDE1gJDgtFi3jgVHth3cyL5H1muQ
9jUI0LARbSaUI/Dj2x9QOZdgVVGTc/pxUsXVf5E9rLjQk+JR86dUgCEXw7NS/w84U542kgs3DdVc
M6DFi4fx0hQCW2Xr/YX0rkZOXv/cemg3/FNwbwUTnx6qdLjeXmapO7DHwoaYqiOaoxpTClOACBBP
1VKsVxC13mH9RxNJxCb2JasKghFbLUJFKq6bWAUuhaUsa3mCZYy8RByiuZEOWVbl+rDImuw3a0lr
QvXevSC5hwo1spAvoFxVfU7bz9CeT1RXNRS1IMzFAWmprBliPzy+LVe863vD2iP6h0TpyIa6tUZO
xPBjD8U9DoTDmxS0jFtznLHZBhKaqfGu3R27q0xVQVE0mu2+kmmI+32GmOxz728VdgVoOvCE5Ikb
NogLDXChJE/+CTuNq7FTK6RwYFpKWYG7dV5Yt5NMOhvQbzMRXuX+2LPT/kV6UpzyHGFJQ4Lb6bXO
tiAtsv/iggiDcgu24ukN7LbOubNmMXRdy51cG92OIi1orEqQYQRxa+hTvOW4Vx6DlO+FBlvFEbZR
rPIIGjqdHRo225Mjo05x8ewAl9DRIFdvAWMd8c91KtOVGLj3OXWIqyRD8lpWjUW2rmPQtrVHa5g0
5p+znEXmYaHYJ5az/bHq8JRPzt0qphlHDIX/NJO14rZhmCsEOgmMar8T/1pHXwFNO4bIuPhVaXSB
vC2UsS8AIx9FJmYwOkUMs1wZ7SwsFF62Lp5mNX0cKk6qMwbazvyis6XR3BNkRMGu2IKtxgWCASWb
GD9uC/KAGx+CRu8EmBGyYnZCi7RBqWpzQ3LbGguMTXUtb/NQf67RnAcV6MzcOSx9GdRk183syHUi
afShvPRgk7HVb1w9fKSEiiv2A2O1KkTo+X4NDOvAoPQst22OxYZVaHOI5aniq3W3ZrBPtOVvRMh8
T1GG/6rnoouTGsKYnhRQfRbukTdUUuHBNREn5PauBdjI+t9U0vTag4zVwjsCadvb0mU8cX3jFP2z
Y1Hy22XShgEBOK6HZrB5lfm0bfOgZhHsNj9YNiD7U1WbUqvQm0Xgzgg9A5rGfVuEF4P0j6ztSRw6
LxN+kRwXSfW5kXI3XNDtlv+/re9WU95LEfpUm2ssFWzXOLEN4OyL+U98MSYLUyPuyWQf7qwbvEU0
wt710qlSQcetVg2qQ2SdToVnhxi+vN4bDusb0cAbSGJsRPLHZtfGffMtioUIkD6ADnoRTDmlgM6M
H58zgrPjCK6g//oeWM/w0XSBRtGuUyYSEkAfjgr0dCawqVOvfOxLQJHvj+V1RWQaVezf8dOl38dQ
6iqHZYwApX5snpiZO/S5yo8CX8JnvkEgcXCkAInYxbSJIFSMPhx0QDdDDlCtJTmk80j+avJu73CI
qN+dSZOF4LGYnptKIFkFO1lRNH2YFNV7/+B23bYbm6ECzcNtndM996kL0d18vxHRoaXwdELscm+C
cdH0cAlWXIOWy8TM4opYKN1FAPkkqrA7R2SfcgmFyikei1ivAMUkhQz0ItgKR71c9kMtv13CG8yr
6nrpUA9tley6T4+iFewhkICmYTU3nAbbishq+OcfgXqtxjlU3UAq/rwHxcbpRC80y8YWoCry2bqD
0BxMgtOQ6TNuRxSP4a6gQHKpM0V8wEBIHnNqQnjmeWF9duk194qy49HLv6C7j7wqbQk96nYF1C1J
LV53zPAjDrwutRkuqsm84XeNQGf/eE93DfS8mMsl8fpQOHS7ILrBe6WyB0hbmhEmCdEyS6hHQ0ge
0e2jW8rgQeDass8EsIlq8jofHBi6rxniO5qg6SRAm1sA1pc2nB4QcxoasqDcWe+Kx1WyHeqltc/w
TvdkpiANqwaOoOzQQ/A6j447v1I36hHQBEKFjHRpWgm+v9X2Rtg3HgQZT1YrV+XQdH2gA8U0L9Np
/ySACG31lhK6dGTC0OcfzLZ3T5UL1LNn/qtMzNbHjxQ76dN89ELtFzKBxli9wMEOwNiYK6as97Tj
LSu0HwoFIOzWcTfHiYz4HsXwxYJ1A/qAUE4NWI21y8U08nYR8stf8w7YCOicmUcuTDWS1NY9qYlS
yysKyDuTJ5353pOK7jGlFitMeMdtww7wx4TX9RU7m/MPfh2hTsuGywXch/EJYWvh0nyCROceYAZx
+ZysrxfWjUgVnll/2BT09FMKIb3JBRLLYt/rr17L7bHRJjMGM/ePTD1sG/CJN11OubTDJ0aU5C1k
Ft+wxWG4z6aUnaYck34RDrN79rYqQ0O+ZT6d7NePZrNllA2+2v5B7Ro7NAnViIU5R2YAJc829rXm
9I7u3Pzlz5AMRqfR9aFdgKWrJ3KWVP18Ijrg46Z49bpUMBgD13f+0OxEASXMm6OdoCxc7+drl5w6
CarvROJrCQ1Mt8PIhYUF9ZuGpnStLt/k6AypxFjPlIDpLHE1DvVXRp+Uzyi+oryLZLnXY2dal+A6
vrkA7YdkTfsISm5wC/NE2+2ql4z9VlOgO8vZPmIU9WK5pDIDZzLMNXIjYow8azUIcqCitp2FUPTX
SDipzzZ/G+QQeVzbqPrOcuqbDz09xCAWiDMA/W/9Y+PtOfUuu7qxozIpuGVx8c4scwxNcnxJJBjW
kX8l8QS5gMwSKbXvYNPs4RF82H9mVx4EzIvJnnCpbq0Qh00lrdbWhPNDWX44UpzJS714iy+kCYKu
dBxngRcFnqtDCPJNiwISTF1Mr4bHHrW6bpwNR47DzQkQWAZo/Dp18ZCkiP1Vpoz+yXanS6HQH3Ke
w23IpYBo5AM2nUmGWBHfAW8OFhC8QAsG8sc2CwtDMBcjhC85AgfbtL4tlV/F3vICb+P7UCy8l28z
YD79SRP8lhe7w4DzXexpCEaAt7HUBiKWJb68MuGbTVDrVE3Cxv8P4c4S5xsOpng454GknYUXlL7m
min05swnzFWuLivRocREgP0Khe+GJemaJko1ET3ZKjtaDr2C79NiT5OuKtaNXauPc+RQilSm8QXc
1l0JIDa9WIFUfODfeLe0hk+/k+ODJuz2pKXMqXuwNSfyjyHJzQ3AtJTmDXoIpo0TrhhQKbYon6AI
hMzZhx8R4nFGXAc4scHUeMyvOJ6hZNRxnb8qoXqXxpPi7JveCwQclQwzF3mWYA58z02O1fEM4VnE
vuXZSEIc26ncgrKIi65aO7YX8x3BzlmAX0S2ZJ5Msx7M+Vg9csFLjTmuzRNJzaxPyevRGWPF7EaR
FzS3FzOdS+chn32XBE+lZs+pjg5vSb9XRhWzL36luJecsOQcN+e+IN53OmBQRKiX/7L836jODxVV
dNhruP1h+Ob3gSaO0bFzjGs1d0AOj0Pb36xV2ijxw06Vk+QtYuvffQiqCTROZ0FUlnVPeYZ/AVEq
pWPPB/d/LJc+8/FkuyN+L55sWrQZm2xr/HTEjuGSHDSrvnRgif0QSFLxFe0e8eDU5s/N60c1Tv5E
61P0ueVzS+16NbEfVTWPUbCqEsgi82nUwxyA9yUAXdhVBc9k6PoGBXKAqWeUptbjSnyKHET1j+AD
2ikz9pUJNkqL8t/hbsbICWZLCVXgpY5//ipGu6f7cJqePbh4USoDusHYrM97NUFXcm3+hv5z04Gl
CnFN0UmnGHQ3cGCtxm9eCQ3CQYtBwLPQh7vWHisEXlrykqeU9tsc3d87vmmJVV0L3xQDVw5fcf+v
P5UEd8R3UppcymM35HNupnaCDl62/uiwXHBWtL7SgLg5kHPmSzvAOztVy0ckhF/5wb/U8p0ZwsRX
IAoh8BuqqSWjj4e2PrsHpoleJrU4XU5jKjEx1IvoBljVYi73rn6PSADWnTujZOtYaJsY8f41+3Of
TXYhF7i1F4uOqmLZTSBy/dJXgYIf5bGxWHFWqB+JdUJxI83g9QlZTb4CtmUBvByrjgjrZXp71vin
gmIqMlGJtsRcKAluaG/QxM7jlFgBPlDyrrVM7q2ziaf0TaCgRCWR4hN0F/u0NF8yk9fapfw88DRc
pohoTszM9rOlZgBwGnpXsXUj5FaqL2hABLB/smmR0RI+3pPaKCKHIzfIchmjecJ93tCwCMVLnaUS
vE0QGsdml/FyljMkymDMLU+HvjOaT3blHy+KE0hBL4IziIEoZKPbFyupH2VhkBHb39Asr7tLjeJh
YGgSuqmSYo47VNpUeGJAxAobd5g7qU+5vKdcy2OnzoCs7x9RoCMVX7GXyO0wc7T3CfQQSp49rhWq
7USMWec0POwR9RlBXNbuFZK8cbnqLcEg2roPw6vyoK2FRW/cC6r4I9iAnBiZUNUkdx1ULERsMYxx
n8ivcbqGl3DSNpNdRFMt50fzTXErLTQm7wXTZJohsjQ7UqVO9pZN8S6dpJtmS+iEGGzL3+orQ1xh
dpwLJ8EZKtXzWMEximPYF5nE//co8lJ83/JGRuZNT3EdSntoQ0dZleuomqAAnTMHeSM0D+SvC/FG
5/DX3aFGvpTAEnmh9qCZ528EOa/6tU6FmeYwtpTquOJdl9N4VSX7O1J0/cL+vgzlcGAU0G0q/E8X
jzIJ8PhCKXDM9CDQl/XwMqAL2rmv9JfJmQMdAU/+e2+v/S5dJ8at0WwvgOUpNrZfk+4bgH3pBWeL
ihvqQloxQ/SnbD5O9yKSyCxOndG/UjRBl4yWsdBW59Zan0Am+V8WMweDX3QtMhCm/jfeKFm7J6rN
/RGV7GhuJbciE23OPCbfzi1MDcmBJuoaIQMZL6UWX0RZyA3OfU5Hqo3dC+GgCi5JV7HzZUYaYEfd
6YCnCJ2A1++9LMBQLDRJCnsbea6fehu2qBxvAAkHMaZfSFS3FpF1RIss4HqqGUvQXcZC3bLOSi2F
Wr2mTGyjNrPbA7p+VUHB4DjhixjZhsLThkBzwbyyBSGyooksomJBOiiEE0W0oG3xIWqtnPyZK7XJ
CEVczGlTQ4O2BLmaLb3AAy6KtszB+oVmt1DZ/GuJyS/fxFQnB3k+v9AQBSKxxu9vMGiCZGR3hfvj
hrQCCiawgfx+BRQb8izxd38Xc4zm0LHyOjd0g3jvbaKPGKalbpA5T49YuSHjwnWx/hN3tYJ3jecH
d8EPBa1VgZnOK6ocRth6sY32s7fSEi0Vmmo2jANTOA5iifjw8r7i4/hvNo7x6b10Si/HEawRfL8s
J0xbbDrpbaV1gg4exjdmCszDxSKLJGMGrO1Pc+oiysrOlJ82z7kquSl2/szMV0rUpnZTXnGleVWF
qTpa6rCxg7tGcP93AKTRlyP1tkvDfvhYTjQA8z475ezi+v4bR2pDUQBf8aIm9SAnYk/8DLK+IDjs
ajs2L5u5uJCaa7fK2HCa2xgp5nlsO4jHTWK0Mkt5MEiPhIlsULfvNNSdIMINyNPyo/iEC9AG7o9G
n3miA2QoP+a+V63fn7YOsKdKRtsoI21JqKRVrDMBSAKsH9b/CtpZsoql1a8GYT7IWhaSyBklDtVJ
hsSD1pL2jaJNJQZgYJr+XOGJEyDXmZ/lL+XwFqwAQHVZ37OWq2lqbdpPsL4sRbOf7GJCAy4HOuCR
9F3zftAVD+P+HTLcko4Leyt6BJ1gHwR2hYRksUabkWNo0Q88omqEtdURnGqtBNacDgoIrmIWSBok
ho6eRZRE6+iGVIfiIisIzAuiBSYdsAtj2NDcVvvSgWtja/5Z92dqkyX9B5qKYHhCg4ImClLdwbhN
kO1kjHeNeCwn8DHdYMKTS9g9xkks30nmNWTFQ6cK1p9Y5TE+t15Q2MZ5u3jQ6mklaFVsVlpT0Rww
0Df9/J+TcgQ+9fIbJSVHmaPM7E83VYmcp6ot7OtNO8b8adCfvqBzl/InbxJH4xcjAPy1K9fcKVIw
FkQdEGYvdUYhEpcIjI38AttoERoM+pzfMopOx3UwtepGHSiJ2IfHjd44ci9cabQH/654kY4feyko
ohKNtgSXdWT2ic5WDCDpoZlhcBusyLbE8PT5FucvP5I1X0WETbDJ79IQ04B3bL3Ad2svq8enCJ7v
x6T/AjFy/P8abBFQcNarUu8LIMF2hm+5PSEWsDHNt3R38g3fM+BwVUCj9FOCFw29zUSIcKVY6Btw
ljwtiyiqiXc0ahdxVR1T34PeFQHL5XENT5tlFbGF9HSovUuMn6bfgjMKBxXPvHYBjGKrXNSXpLy3
y2Rtf9WdNhwCe4McR1yYiJO2rMV97d25FWoXS2m622PP6ESGZcd4C/rPUDQLfZwxKgqO+99QjyuT
pQKqVLWRYmHicDNmxeoA5zsN7rA04wRcmCDM2TU2T9txh1m3YgHI8w2G8OJM9CmdNKy/YvP+Nx0u
rA/DZP26DdH4HzY6v8ECxW9ke+1IVbYV+fkNZw3Y97LwSMTfp/JKQkILN5VHXdMc2JJF7FGSnrJL
yJXeu/xpSdcL9xlGIXHwn4dofEU2TyCH8ocDLjW+hreT59Lf17KB48gpZVEPdCwP7k1NULQCtiTR
Lq4AYA96lNJisELVetxFtrAu9q3zZos89TX66wPR2okWxePGrTBGWiHpB0zCuWXVik6OXCeCvS5N
gqTf3Yo66fBiUL8sH8z8TzMCW5N9I3OeSjH84aCSgjXcRHPxNX581m6qM4oMxexlgvKvUxCD81Q/
kYE673DyGNJZLMYRRHq/LgmQxugNhZN3i2xm4Yk/96VNQHrEmafj3ooPf3HxeDu/xbPVgLsyt7A9
KQWBxymBmD7KbpO2kNOI7L2NFcmMoyucfCYvYL6NYcwL3ZomVHdsY09o7FPU35vitWX2KDKvMZq2
SC+dlsL8HsSDP5OF8ilr1Wu8glFFqzhJcEyrrKeybNbLTU4mFW7I5sS9thK/2U82uePDlkubH+0b
ujCte2gL25s4C2dGIaz+Wpd3VUeab8d7uGhBzWcpBGPMvVmNTrKHchqXSImiwJ3Zg5CvgiWm1kNj
LbfgpYIcR+GFoB1AiEifX4euoUXnujkGzmkmNVgaRt0vZRmpHniGqKl0aIZQIJRWJ7btXAxv08Le
O4MSQy/uy4oSEJ2kjHWEISbnN89ATMckAtY+pgQR4AZyiouJGtBgTd0Zo5pxc4Wl+4Cb8u8C8RYq
HSXwnZtOSnACjUohEDpXb0vw8loGOjSkVrl95HJmEcLLWRjiHeA1ydl8PqHFb5RxW6xNbW3/b9He
57jmnaj5D53B97OunMS4hfOgAZ2iNJ5YgLjw6eY2+9g///ccSTQeIDYR4uJ5MPQigf5dYBc09L6v
Zbvcdvn+BC8iFdURnfLBIxPaUERMHsimddRNs12bf6MgyYhDjvgQt1pcIW1pZCV8sUhBqnDp0dmt
GT3xnE3kUHnT5Hw/5BkCy7NlTkeJOIJF9Qt898grGcdCjz1th6RksaI+/jjhJ9bdRIYFaHHD9oza
WItk0sO/MTPDq74mcAudonsOS3bLbKGJRXXGLsMHoTq0RCLU0TB3wtYE49QimZZgM+FD4o8d6/nk
KpOKLoPsUQByG4QGPlQ8QueoxdvQxWKKVD9ZQN2HyeJpkN4MQazoc/rwgifx+DLr1w1njMHXWLGy
vuoi9qF9UYupafOxAwmDnDXD7hKlx35rEUNvl/r75Frvj3bXwjC0r/HQS7bTO7fnAAhunLFFzSU0
pI4iMHb5X80qW9TMXvP0mHro3YCW6equGI/9XMibhGDEQes6kRgs9LhFIEczZhXm2XblbWUsgDPL
BGk5EwQtvEY0rcGyCU8CnBpaHso9cMXoaVP/oPsTeGdH71DS7w/g5j/a1nOGf+yCky2tZDVKgJl6
OSi/Fj1xgguMwsJMXoEal3xXkS6ZNmOS2VwZX7Ix6WXlfhTXXLetbbnvx+zOsGRL34SjXasyeqnL
SCFJRwr1W+N27sHTCOpdsYy0r8D7UowLyfrjkyBJ9s+YR9mNHqyM/qrlcHXUlMBixBm0glpXUd1W
HY9nQLXH+jTj+uqvBCJnfwGGUENfKF5+55VF6Kh2Tm4u4Xe8WRRqFGgJ6a6u5UrrgvdCvisIbtSR
quI04qkgWblAz+bW2Yd6fS7J2tkpTWTV616JOhATmNoS4JGx1mW9VeIuNjmkacc0FjIO5yLpBpyB
zPSUYSBRu8e1Bljwq5YwJHi5iF15fQPMsKxRKqvunfIn4+GZAoPbiNEl8FXaJwg462m27rUD9gl3
IzAuH82lqAjElDktddCT5P09JIKT5Ol6wnOYh//bUlxjzGHymN2h+f4BSasjFI6lFszO/muIRQJv
y5y9NCeHTw7KP+JaMXx/RE8OMKHyl5Q9iGo7i46+fBxvrjuQzzwLHAD0CQNcNJh52gDSuKTVL3om
vy5jNaNDw49A/Fcs2K4Sa87BJBFpKcjnO+scPSaxsxD4l+rYap4zTwCG/Qy1Nr7sXQE3bF5JI/Fv
xbKTn9XZVPIKmbEjkeAeR/Oqf4MdDD8foc/LdDqEDtEP3liRIodrjZ1gDJBHhrdTPalpPLsLAzGz
1Ds83hcbmiGyEhUq4CKv/tErV6J25mKLo2Zdkkp3D/G1DZ63Q03Us5iHpMvFyeUNBlRsm/14TW1u
vjPayCgiIwkD1aOHLWqwiF+7s84NvChKS6n52Py3AiHdJNEaD4rzVt4LalKa4TkwwCLrC3ZYK3Zw
VpR52mK0EpZTzjPe0x9CJqT06A8hXBZDU5uV2RyD0VwRL11pG6iYVnx3owXHY8ElR/K+Q8DXKElC
Zd6NR17FxPhvnHGRgIPn4mHh7d/BTWyq2yB1ZdOTvW2Ut1ZxKi8GXkCscI7OHFonn9obKnZh2I+p
YwF3Ns8upAx+e3gOIZzkqeAmhho/cKeq8VJoHsphpbDCWcXKUN1faXV5y71RKqZmhuPf+S9ZzLeu
91EuRBQo5ib6lj0kaRkvAqsFJyDERQxxEp+uRfuFur5LvPkF/hIHnMO4mDmw7lg5SpKnJI+9loL4
MIbHCpVpC6YsZ7hVxLAYHzpmmwL0pgJavwjH1rcVD9/qzFUwNwmr9eoXMyIO+ogdiRlKSkQ/SKT7
XIKvy5ki9RSj0hUxXe4GjY/x3jAW8PtjeyOTuFrNP7VR5YzFFS7NtbDsNCgpIlB1dmhC89voQw5g
ptNjKmJdUdFQpwnpCJiUoriNMwR/l5bFxRDzc52Tqi8uGHvtuNgJUU6yXE8kpSpJTRcdovFF00pZ
w+hgVAXii/rZmf8w0xlYfY3qQ0z3+XGjjP9lkAR9XowcN+DgAMMVMt0mOhtf5SJ5uoov5zog/32v
NNymOI6VgK2IGRCes8c/sPZiODwXu6Djy90eMmbdysIWZN5JUmQCOYBzauSw7BoyuT0ghDyc15qJ
y9WyrFOqdhqHwEQwwv96MGdFT9/GkD9rtQoCVM/QnFZRfodMs6Y+UYtw6dzeXRSMuMq+xtkNZWRZ
1nexIVSzWrShv5FsvTvwCHSfGCx47QL/0wpb4V3c3kkKWpU/PRDzah53txVxiY7W26Bqr3jLoKYl
RdqefTBLrZSWYUWbuM+4dXPpm/STJ8X/ctrTX/QKf+27zWmSCgl+OVGE79syDo+ZovtPk8MiaMBx
9r3TpUY3Tb7aXPtrDpvW3zW4Zpcc/T2S5/mnwZJo2Hbe12nhRuzAyr8xZdMYxCqRc76C34c7kdSq
SsACyppIOMGT7+8zHfVSCb9eEFbAVAKInokdymA9jAG14V52qLzXMvfbfNDQwWBKkWCHYtFW4S4R
yQbMaEUBnX3Y2AbSpsWOxtXpqya7r2uy3s3wst40evHPJixrU9SgHi4zVZigkEB00vUWuxeABgU/
yIIJN6fQUkSGxyuP3DifxforsUH/EU1kGA/Sq+ygBiU7x92ndRMB/Ni2BTzP8t3CHmFLehl09NWG
Hx7Eqa3TRsPAE+GOGOjMRxP4yPFOZo4abX88Fum2lsUWLTRlcItqpNGXSJJImMA5Ok7xC9ZG3gt9
S4UKXE07XfgracpkOTPdEnyOdID+4D3OXelJSu5NPN2vr767Ke8Th5y7sO0x+TxYCTeDVlMGeC8Q
i0M1aoea8/Q1TqwOLgoY80Y6gCXx4TYl/NQOmM+FNaZKqh8PBKKttMO17nGmSIP+Iw9LvyP19aYy
sIsovMMRcjmjJRu2xkD7h5XnBmWvNR+qPFBZ+QvTobtR6vkhcURESz++TXvxvg/BsXQnnIh+JMpK
5Wdi8ZBDVg5ZGbI17cHKZ4mQGflawCZ+MHoJb4gvNLjd0y4OfhV1UZk6HwU6l5zGPhUh550/V+B7
7OutA2CQr+ZcNG6MdIWJUoGhgmxhBaLzLDs/Qa06Agxw042w+Um4+jAZXr4zIZML4sjjWhc2bWGv
fqi0WbedD70wBNV66ghX4xvUa6wWy+7X5aDLMVGZ48D3cIwANXrLewchk23hDKBucAa2Ru9WAvnj
+mmyK8GKzBFtlITZnQtDwljYQIwhrkZGTta9jwUFttnvPkni+SLaE9mPfexUQn+G6sCdGsBgdRvs
yeHR/YGyaFB/sK4xcgb2db4xK1ZMqoT5JvqmDUi/cgyfZFYHhxbW1bx7iWwF8lIMW3iyX8bWkQjN
O0tEwsnOKo7JdrKzos34ZkPKxk7rjoiYWi7OEHa81zft9LJScG0NBsumDFHjAd+YVSmcmPrLpwdx
DPI/uF2hfS5atXWKJohp+5/xWdbg+eZXx+XD0vsK/wKCKCk45Dp4GKbhCHYqEh9t1lHdHu9IxfWv
omkUDotNokcVgFwW4b27pm7gU6AJk3L0AKQDE1tjyXMIFuQXXkat4filrmx6v7YlMcmtEVSE4pFv
UNq7g21QXYjyGvCE438RFp7Xa/fBJNw6hWuVdjNIAB571vuSsgVrBQfozDw2ekE9U7+Tm/W08w4l
FgiyozLkamF/33yQ6njuIoKigc/R/8nCG1vtBQ68xCORUt8T1UMSd10xSwnq4yHpwwIyXjIHSlFi
pWguxp+sxwkN4+7U1/VgCeqfI0E/wGIXbxPxudQfJv5p6x7xC4jLn2Oc+O1S9uUdYjBBRPnKZAAg
hKI8CHeZjl1xy82ES0dLg9Z1pdbtdplW8mkXpu3TLq186ToJ/EJgCS9NyMe0NFqKBroky5xqZEXT
9ru8yTFt7zDGf5fQ+A7b4SbBb54rRuEiux4n3FDNdzika3jJGI+ZMMy4ysJEhU/1wg8dy5U/BFr1
1YXUIljXhSOXIL5SfqdrmOqEEhlethzAk2mnRyftNvqemh6Kwa0vCiAizgP+TAyMgHr4O2OsXbI3
BSNBl6sAe5XRs0Ot9R8PLUzFPI9Ej6re6QJbHvse9teZTS4EN5hoQtt/5DpFDAyEJKkzQ7XjHNAG
NWr3k5HrtPPA3tTN6Q7LRwYOzG0Ps4zx+TaDGbWzs400+wvyyGBFchOcMwfnqiNkZd4Hq+C1sh9p
23o02XumPJTtnRrh1vP6tPwgdhcKpLL37uWc4z3Zm9TGkpB5ckYjZ1+fOUsb4bmOku5v50A4CUHW
KPy4XtgBxli8Rqjhvrm9DgGpDnpP282A1NUbcQGaYvBRc+gHyBEooelO3V3AfcV1vmcOJGhE13nG
ZHD6q/XXYhRlxX1psIi0iVYM15yK47emXe3GLgRJSNlKRen6WlcMO8CAv7YW0KIqQu5i6w5jU/NP
yOJ1nP0ATjP3YBYzT5cmYsssWSNT5KSbQOxme9axgRmBfszqxMZCjR3TJ3SF8/qkV/PNgRywbrUQ
IYKAZ08wjZknitUfvjxTQsEKRElAOEDyMzzf3JWDqhqua9FV8uBJsGaeYGzJHtAWvVbOX88c6uSr
kerCbEAO/1C/p0rabzNBxLBwr2d0sMK/XwiYUttX54cACKOpOosCviyiV91b8FPoLt9U0RHbTsmh
ne0komwJIyDNUOsDO4S7OuEUN+L76YQ8WBgiDLQfgNoAI/L9UofQhkl/sR47+4BQb8kBEp5ywBs3
/mr21ytD9ymj5hi6Ya8AEd2/PMBfTRUUoOiND0MY1vcmG+c/QZ0qXaeEIYVhzfswNhwotinx2W/B
mJ4DNO0GvzvKWaaDqJVy7T37j4TDkP0xCLODJfJW3VrtzxxNESYtL3599T3kY5PAEhSwcAjoF1UI
LFUxqyKv/3aIyInJxowrVID9r3EVBGq5K+foGx6X1SARrcH71Lr8VeMrxc6yiLeo02F+ufbg5xnI
GCQpfpN+QehrWen0ydywGOclzS4hbKOIbE4Lw6zovnaz5cm6fyJCmsUU9ABNS038sgEmjibM6Usg
NV7VO9EoHPIesr8BInMaM9nxSrDP2MO0ORdCPOCAKvF3bPwu+/wL58fd9STleyIPh4T4FBCHJEhV
hhDfV/mu38GjN+1SViz0O0UWTV5mVh5VprtdDZR1tG5Y0umfAiMWMbB2KshPDthdRYKQxvAHh+RH
0cHgsNqCpL5O3PuRZlo3wJRMHlbvwTqtB81sGtgtO0n1KL68x9+xsDJU365qMfsK93JPjEo+C0qc
3qnAFMf3ibybrDOavztdx284Yx0PlaBkrAAQZ1p7rdmLKK5nCYb7BHt6kQonubNJu320Zu7ZvRjA
reVKI3AF/VcL2Obb/fFkbp8GnNl0exNEGbrWc07/pgqBYY9vzAafibfywSR8MQ8oO3aw/2ZUmCiy
V6bHYV4UzgwtKFxq3Ge+zSqZNIbZdmvRmX7z4uJbT/7W53YJBrw9Tuk9mtDf3y93vfXyu31b5axP
unzwpNgCqIFv44N4IX+t/CpJhSrIK7uCbVkwRVVZoV+x5Nt1mdJ9sLkizjoFghqO+ZnYpZraq8Ag
ZDhZorrHk8KGXYXdkPNuPYad2W45FNaBXOaumysKuhyB4L24aqE2+VqWphHPtXm2UxA1jOAWs7Y6
pX1s/2tfzvw+87BiK6BwYApTjBpXx19cL8Av0sqtbxsGzh4dn2gWaJTzbJbRJ1c8jjHFI8vBWaIj
NEbJ+EULLA3rGSAUtSYgkrS4Q+CUr0aZr7yebeOh5RO1VNOA01qnrFYIMDeNdzgOZ4rfuwVSHMcG
JubqFmXygQZKQOnUQAJirNCk1vPMXhjq6fnMLreZApnPE2G7TuQWdJIY63srX/euja64Gpf9PBfK
AptBkifw81xsdxc5hyR5qll0L9Xtl5WykR7NpusnXt39AUrDAxqeY1ZCEHRzRw/njKnCjbwurs9+
b/sLL0xfJbSUyyk/8tBQH5JlMfj6Y0YTEcXAx+VlcyHNzENur3VlCvK/gzBnKMCpJgJXpjCYXdBo
KinDgCe283bbEw61EhT+xKBWiUwTwxJgd9538I5TEMZvZ56gb2ykCbNIS8468KTej/wqG7pUgPU0
/mr423MeyshKWH4UKEuRCMT2iVje7kUgfIZblzpLVY+kvCF415TYKDINx3dPzL66ePtf0Wh6XDvQ
zf6WtM7Ac4qX3h681iTK8K6huMC1zRIhyG2BUqf4KpMUfC3LBynvxfUi4nxsJVIU+4P9xkm8Kh+z
2Blph75+aDCgDrcw4utLhXT3z64tkSXW7rLVWthjz5gVUH84JOof27SJxu9R8uD2H3saUTz2XSKO
t963zDSRyz076rYUe/SJkcWRufQ+XlFRcb45sc3pg4USFXp4Ew/9IjeyBugWwjy/ZEJ0uxWakoLn
2yWgL+F7DYwOxm0vGlajpKoxc5cEHVk3J4DI0eKP+hTjRWjItXP7x58hDtDo0Q/qNlhyFNgNw1Se
n+wKe/CPi+MUzJDZhyA63kzqPP19ihc0IoX+p4Ty+7Tw+wBPy54yT81/Xbde7FIOcHdJNAL/xcVe
8Vo8M0NcCu8Of1MFb90ZNoJ3wzgtFb79yvJ0yN1vxfiV8qRrHxz72mzY4I6pisPiZCvZhXKNmxB2
yP/7NdaYOPt9pk+a9Tj2gPBmSgXoZDijlUcaH/iAT/Fqk5AP+61puhQtcdnBXLBxOpUFStVqaFX0
XXeEYUjX1S2WzacKv5XOrwMCU4yQsP7pn3KNO/e6XO/A83GikvKBdZWT1JCve2jOD18FXr8mjotX
kwHSZZj3JlkzGXD8XZxIAtK4stYxpIhL1xeNcvXZD28YWUUegqcJCV3S6mb69wWmj+FP7nmnhr6c
4MT9j1L01XY6Of+Q8XJQ36ZWX5LXQSVbhALRSoxFSINYo6caoh38OUd1nRVLEEp8Ztp6HDrIGAGc
KA/GQVhAv3flmtaYBA6gZQ71g2u2FaPcL9U47aVLIofTKtYbxdlOV6/PZCgxxgLb4LpYk/Gs7072
kvRimsIXaXTnkupwIofIWmolIzypA4Rq79UUzyY4T16a9LqDG5/NwhMeqWXM2ad9MjYL2gxskUPN
M9mjUYaNI3a3326wwNp7/Ih0P9UCyjtD9uLPfNF0YHByPF1ChGarCoO+Ib7CbSMefdHfOpMsGR5v
sPz92Py7rDPCXlzTBU3kEL/5nGiL6XiVIkvgSYCzwjZ6+SWBreuRd6urBIvZ2fuHdYBgFcKZWmrP
c4X+cmegPSxf9jrCQGeusjOcvKbiEmSGlu5hrOjE0f0beK2SnXmm4Av09KH7AOtErR+U1cVidL4z
Gnt56diePTP0b4HfnSRBKQM3RFlwKVCZ8P0iewzQq4AhbWkBxH7fbMuQTzKMC/ZvEmw3Suxi+sIK
XJuOAT3By8BH/4mcxSvfeEbOwMrHsn1He/HvKw+GyehTz+Q5a/fMz7PgNBLnZt6Bjki8sLlxuxXp
UJhQecOEnKcEBxDzB0EexGrGenEjTRjt0+bEZz07+5QPCxUxPiylq04LRRu8qrYvlXQiY4WOumH2
sUKK5N2Xivg7UOc2zdW/w/6RpTyQnnMZiBq20zr06zeFOcBovrSjZpJV1UYlMnP+LnuGvW3a0euV
A3ESA29BF42OPl5HQPEN1CUYrecPCWEjIrk58OHqt+AxxU687v/s8upsazkNxv6AS7spTmNdbnBM
V6ma2T54WauTCnPnZNbLuBTCDHWvxFqhb9PrAIwZxq0h76vBcSBtNxZV2Q3BaP56jwis5++fe8p6
VweikuYKJ5iZyNKyxBSyEhZPFzLeG3fte231GlyGEZeM+Fw66fINokGRz1jR/EsvhLaMr4z0aPCG
RnmP+pu9Nw2kwk9iwIeXTy3z0M355OMQU5KHrdPv8waEx2c3pka3ckx7FQgxm9CB0IkqSMwHrjet
1XGPiCpcpc/LT1GbCVCww3MLYI+Njj+5gXc+1Ejd8Rydve/O8drl7HrvALswsLVTzP+OExctl1xU
KAJV/5pRXS9Qizwk2ZOwLCWYkfMr4iSBI99L/UL5jCDNP6wbUfN9JojmJL6OqmT5kEr6K/GUTYTa
20XIdGrTqg88HucJMRsLWk5h5Vz++PkU65jMywJXKjN2bzS5poWVqUijEVXXnLZFSPDJp795YrWY
49uXGt044En5h6cUwp6hJgtiPndaZ67KMco2LUQ9E+Q31al93kUWJ2H+ShCxA16aWSxVyLCLGYNR
NKJ2K6ypoCQBBNWAk/WqzJ88iam+wKHcXLbIX+nb8TSIMX5Ho7kZ+lD8nP5Og9whvIv/U5v3D/cQ
48GrrCWwvBr96KBM4eoH1jv93hwiyuiVAXVdUCKSK/VSTfUmjwVmz0IrG+TEYeHF+R1+XemPbKgd
jLBhaLjaGOQ4GhnTDUw7XJcQdHQX1dl/kGoyw4Epr8HF5xVEOQnEmlZYgbxjP/HjHY4Lp4etamt4
ndXirnYccm775hfFkAF6OrhHcxTCDqu8NLGE0m2EZSL/XECNVx/plE5SnHI6DjmkC09ot1D9dsfk
2x8+GJ5GyPQ9Of2IsiATEmiERouKhtKprPFpOkmqkFFwhUGLhXqJ1NmnY+PwA89QOUU8fLPgB4ZZ
gMT2RwghnfoRuE2lJ0GnsJj/a8YdJ9OsuPxe+gz7h8pwrQriWD89pJ+tRFI27zrhnDigNuVgJxUM
Dyg+86mfmGRjdzougQHyphofT4ZZw/G0MAJ3tUfutHe0iotZKzjOn6Z0BW26uvVmUFLQ82jaEk6+
cQfQGNrWQzUWebHXaWk95r6B6DzS/jX0CqaY5wc9AwkqglnkekOPI2fZ3levKMtJ+nhmY+KGCMRu
WiAtOVwLLVPGsWXLFJX/NoDpI0OsyLuVFSWj7WduOHM0UhCUBZ87aysimBu8zVUzKT9PZf47g5y8
GteasRVImPa/DK3/sGf10mkDjoU5U/0lznIhpLSkcDa30nixi5n30yq3oIeQUQPkZv+YarMG+lfT
wdh4+X9kYxiT9XFXPkSoKPzszyqiIuiNS3XJPnCG3awhHPZMcrv6ah0/0TX6DMrBcSirDtyc0TCw
u8SLLU191KSNfMST4D8TXy3P7CVPSOdTnrhM7yBeWm3xORbOcnO15EC1ndJFa4q6rTla3o9pvJPI
o23I3/xc74WvmKPa9qbiyhOGZ/5aNhlQqFfzS1XmH5lj7lgnrpyFWFs2cSj0xQ9tEnv9Kz5bEBJ4
5F0LnpPoDtcI70Td4ArAqXyDTO1XuEOnjc11VvOW8kUXf5dcclr3W0tN8Rlzv6M1IXTMep9d3FjH
gkitoNsp4m+WwLGffWW6YTKxe4iXDsMuNIioOmC73f1oaKyzGCAx4WIX461pv9iJ23BKu6ykwq56
HkODUXmqQyHSNeynx0B13rcAlZZnhR1AyyyugI0iXkt618VNIwCDw1btrXV9cnImj96NGGN+IfBD
45x7rIYQYlZ9o6PG0mw/kD2l/A5BgavNmz2zHXLBQTVMszZ/mDr8ZvMAHEt0hqV2XFREoreYDIPt
i16k7Y7/yPYnv5jfQeb3AsV7X3qpK4VJlpU8LPPP/dxiZwQTpiyy/vEqEmG5NptGGc/iFTSHCsCH
aZ6PjR89Ux3NLJTzfdaW2vA6YPpejzL2aMmwsT7QHZJ922yAK9vi6Bg0mGJ7jaF/jXLBvowocgcb
eW2A82iRNTIeP/OJCfv1QZ6Qky8Lp0h77jcL2PcdcivbYDJDAxDyRY0OT915uIZ73cK8+T/Zm8EK
jtkbHbP1GFnVdlWDlbUTuAuWzdC6u2kpniDBWbnAuxMUxzZfy0uShNheVPx3a+fsowikkF3/Oo4D
bJIdthDHP2qHFnAvEWe5plGlu/NawUXBA5NFAaiVKSiZskdipfCJuyxkhlv31qUg0YC5Z9UGGzk6
8elGh5VQ1AHCcXUZ3qsGsodt4GdNwTe7IsCM3ELiH6U6lT3DGq69GPbvzfxc1JdAVGLPy7n6itKg
x4YCInDr6FHQHtCf8+Ze6icb5lxCe16boZtHFSMyubavYR7vpkB8T0ZPQQi7QCERVQNRnnI3dgOU
OCs3QMVxeTbQcgNPsX0jTV2SVnz3ozSEmFWbtELu3ClkZ8LRDMegn2gUPdHNqx+Ry0Im0MjW1lvo
jQ9Ja/M/3qnhMM3BEKKyfFw3oiDE+iQGIwXSxqbvinYBXgfObIo1cvUxDJACmPJ9wPRIwhH2UrdH
e/Zhe7NHD9byLzQPZVkhIS2RCzoSp2/DNumlLJVs6utINYhqw3L/B/aDZS4EZ6PeWA8jyJK07CXY
mlkVe1DhxK6eHMQaKDrTDT3xYdNDQJr3tmSzWpYsOwBLzUJPPKc3ywyXVuMDFHQdsQvgGAeWwPj2
VR8ir+blzLbMg7rq6j33sOwMXF12Wi/wNVzTjmobB6KHieLvAkMSfBkQ17a2PhIDdYdMaQiNkXWW
pT5jBaGvhmpfx1IAp3kIxu9+j2gMkaPk2tx47AYehODiaXBuctQ01kIyH0snQpNThQ0AjmjU9cVa
qsGZw7vgnG04ycOn5pmfMNq3bUrw9qrA8zV1ieZfNRBmoI4qQphjaUyoACTOV9HoVZG6thSeShRv
9zG3b9AvFz0O4CAy8sfU+W+h7bE+Gr+ru9cdhAsBI/salgmZHSroLTDEj6L4Ujb/Lqc6lgv8T6os
7m/NTHUCWKyWRUi8tGOoX7epbB/d12ZagULSumgK8nP4do9coOTeiJg0WhZk/VPiDNJCAe9w5OOs
NH0YqerD0I+AeEp1nmEoXj0YZTaDh4Pm91UycfF91ws/oUltaTb0+uUoefHqBDMP5AsioOZHPBHs
z5+Lff9un17C3viIxnbIc1zt6JoJIsgS6nZO/pYYqWtLM3qAqwPHLhUG+TX1EnQhGVzR55mLqFb8
sue96dIvO1I4zY3k7MkM37PzE2gRPbdbvrEturnLUIVd06u5wKii/ekiEdX1H7iL1Fub8M6SAYQ5
/cg2fIL1owwGDfHuJhsQiXH4xKVq2KM938z8D+eucxZVL21VzwtVUIEkRHZD4nErKy3g4kxc87qT
O5hiCwdjjIfc+2V5/bPq/aH40h3TMtI8hT5LfGMFCyJvxLeTkUxkQ8rvkZoUkpn7MrbnrMgtY5jI
ktn51FixEI8i2gXu0oeDNcAkRJuwwabQAIK2fn3n1kKXtoiWFeay7GNOPoijgWzPGOk6PRBgTDqu
eUVTE1u0ze0lfTJZZ/PFXd9maYwOLp4Md6WQbaGipeI2EzEoL9qTgNvzTcAn0ZIoOdcL+CIjHHZ0
UZRsJKX9ranpyaJ8Z3coGDjHSuEr1sZiBTnCi0tGIzXji1TY+Y85hFcZB4I49IXgqsHlmt7xLid1
vmqHytHoC9AlmN19uNlPPapS8pFchN/LrdJiarCpcA0MgWFbHKh23h9pMUVJ7ZiI/rftGE/uy49S
UJrt3maX9qKdGe8wTlSl9uL/vGfjgDS5gS256C6ePVufBIO6pm+Y6/Vte/AVlU+XwbVvtII14m5U
qvFWJta2Fag7NpxXZzfLqeaE3qEP1qsMwBZoJoEyQpPxZ9seeLp07MG/JLUoa0oQwCU+9bdrhO6B
7d/bqZfmX1YjXuDpGm9lQjRo0jeLWsqdIm6xvsrONIaKvSGAWvr/3sjG9zNALphlREM+xBm6devR
yf2Xk7XhxZivFn+gPUkdssZhVmTd5+sUymw8wdvePxcOTGAbjXijamQ1m4cDn42O3VcDB6NpNWls
DRgOfRDgGfPddX1Y/PmgLhsckqVIs2AQVTnWUR4jVTajip8feAPh6S0BvHncnnKQ+OaDQ97EMKEA
wFHWZcVxYSO2BatYfadTv/LPAvgof8qPK1GiNPEpLdcEV0IVZLPugiI40N5XSrp3TJNhCBzfKsKB
kfQRShdp88bzy3J+H96n4uAlx9gFCMzvQJHDhiptqKmevYJ/hgvnFkhNiqCqk7mNc1k4uFXsOfs6
BYCMJs/YHCleOqpfdDbsHjcXzik2JgehSFJMchHKzO/N5FTpaq4uadvLTlijmXkWg7T1fbJpAkBo
8n0ffjUJ+bbypwqmi5BZaCtC5JbzZr7CjU4RKVPf6BQU/5zJiePPdck5U9bqqaxBy9iQqqPOF3od
x75dLWS5uEX5qspgQcXpGQ1JE5h8AKsZMHoVts7PPMMEN1dae37ZDh76Owtt6lPUnrFvkS8mUk1h
KW2bDvJZZrpcSlzWkq+Y/KXL2DqoAG/v7LxyTbSU+uBzRX7T9sl3n1RnhJdjTmtaj0ZUi0L4akUh
Zym4JkzyejEB7vhV9OWRctuVFrx8SMamGu1cQbiHhbPvLyg6mh0VZ5cjzfLxKazPuL3mGFIz/Bfv
Opf1xKExvznVzHcIU2qxTtvHIYFbjanSnIKOhzYbIC8RtyYGUrStr1YZyfHlWT7+mtMf8kalxwiI
KOqIBBg+dIRHouS5yQ810InXeNA4R7TdcOuVoSxDOKUy0N+Ju2qK1Ir/6+H2so1600nbinMK8KM2
Cs8+Ff3HqIfcLC+c2GRc46CAsEMbDe2UYQ3YPqDO7fRKvGMSubsIgDHwa7n2l112ydquD8bCVAVo
6wwbT1m3yETcEw2mar2tyUC3I9wmEx9qvN53ri2Ypeu5MwGWr6fkzRfvvOcE3XR3c4tWW5mZWFWq
1Vv3KoMo92LtkpFgp/Hi3dsF2QN8LKBirGpz32inbfOl+VdZxHB5JAs7hEzZWo+i1WUk9zSbum5o
L70PWtk8o33uNDwCUnQWhIqsSHC6wvFpNDfugpGW/JZvVobexr9GRj2oTeMekw2HB7Ky2vlFL8PD
o5bXMLwK+3PVezNept2L+yoYhTD98X7FqSBZuJ7S8SYmky7ljjybjj/fC20oltBvydAA4bJYmAKk
WANJwT9K0w5WcV5j006jdKKocJ5B4DTLxpb6ZkS1/PlE5VXxDflM7xz0GUyrmxWL+5fR4cHO3s0l
oZDbDd/o+8R9t95zG/Clz5TbCrJfs1sm7/i3P1blXOnuZ0IOLbG5GYFwIZGacTuL53CIt53Jh3dE
Tb55QrTu5ZrVJWOT+t+ykez7SNBOQAWZ+iUa3tn0kfiAW21He33G5wpiZAakaf7F/3I4p8XrLwO4
a/Qjhf57xK+rI9Y5/77itUTnIOAvA/3WRTzV0u2LIxh/7NRtJgG3x79JGhn1XGHTBFTDs6VjUYTJ
nbGEyO+zmL57WXjq7ZxS+5MXn0IyQ7Aq53EghLThIjxrycFD/ISgmCzap1Kdbjc1V0PGNL3f+gMc
g4WNrnNROSAVtJvO7dZovytPtth9bsMpQhQMG3+7G6scQyZ6qCxPbbl6MCQGXWv3d3KZHHQ+nMPA
+mS+6WIyYKWdhx9H9N14dYjVGaAdPUgbjuZmYquFSXT01fmFxKZ5+Q9lxEEC6PNzTkrFvo7sYvhd
X4gGM2uufJRotctm88kJapecVwtaRQ0ii88M1vg7hEn5NnNVXMHYUFir2SLxGlex6ORpodz5UZSH
nsrNndQMG2VxTKI30staMIhuBLKK5uL0K0arDtaBxGHW2Mi1LdOz2iWWOOsfgTp37JRfmU4TmWwq
UtS3+4RiZ6AeKOq8BS69R+WofVeGEfWcM40pobmtORrzzui2jV4KSBseHml/uogbyAbNiuuLk04n
onKxqgCIF5fn6athJHzTDcGXXUCOzGwlJ5EkjHt1//c0MSZt8HaUlAGDR494wdreZW3umk1JVMJT
1kLiQU4XqpkDw6sNnLhN1GxGzZ5mYvJ2OFsES2S1z0TWBwDXUyshdGHoMdqIgD0/+LSOIipoX4Jy
v+QYohgF/4qGpuEZ08Kmp4OAwczf8c/OlevEI0rRrRig1dw4rLZO08cfnjkCf1cnUdxyNVw9ecY3
s3gECQVhhV6Cf8Bf5Hnj+8j9Zk0i28hpITtJRwtfK0q04AWFpH439yEVKE5B34ln0kzo0XQLdm3Q
gHYrihlzj7GWuXt4Qva372oZTQMxucr7UrzBzQLXne95Lw1NcetoCa7bMHsvZJ27EyWKpbFwdrxo
DSizwrRyl+JqLhf9ab/aopAXk/WtvYziyEJCEhpNAq4xe15E0TqyWL6stod6znksimqMEK/P3S7t
yj4eforLTv0ZV/g+mBOb24zjyGnK1ix9bUFkD//xSEjKirLVtv0tKSiA30s9NacmQYpKhjaObRTS
LMafPO4JyxOooholL4UlswZA54HMTA/xSJTJzQq2R52DEHo7DkvCf+6x7NPTFSOoSEoPT9cyzRpE
hStyjQnOjRNeWWJTeQNohbZ695hqUvCt3obTrNLOXzAFYP7NCUCrMMeuZ0biAF3bNM6NkcQ3Bxo+
hi5Np9m7tGCxkLtixhibfwH3iuV0RVtR0pTthfTpLJgZIYy77+7cLDkHMMd8zI1CjTmVk9Jy1uCm
d1PpJiVyj1uzb1ieGWb7xri0VpdUctYLJYf3BQ0+0vYpbeYPZsJ2BjBD99GOcdWO5I+AzvEHPTnp
xs7P9IHSqqSrn6s++5hyWBnvZWxkrfpBqknqn/QJXyOgAt7oSmt7x3uU6/0sJpIWnhFATdESeG0C
rgSfLhzC6B5Amr0WvcPmhapzQuarBIYw9um3s10A7GVBeD5MpazaO1mNGtmLyivSNN6BFO7FJlYk
UtFovAaapvC3CRcZtbctJrjtg/21Pt7GRsHHQoYYoMo9M9U6e9MRiFCo+OODjgSZqYwnIn2bvdEo
lgcXsNhjQGagTYv4I1AWPY39HmnDzJYIJhLpSIaDercvJxRDRr6Y/KPRkl5apjq4E/QitKRCHxeq
uUfqdSTlHHYYRsl6CG5qSwd76A81qevhtOJOpzWaGAci0ReUwJQ96h8lom/a3iT2xGB55flX1ZVz
L6IhgJSdrDJiF0WaN7KnSJWDjkeP9KrGz2UvBGMeKSgk0m8cXpCZIaEYErr7hQB5NXRxIBtWV7ad
scrzw6hDFggZ6CiywWVeU0tTfWLP//PVyLa3LluZerOpl2iO1yb8OCh4Y6lnt/2eHaE1Lw/Jg6b5
n/Rc2mX/zEksctSUTnMUNempSBIZuWQWzH0UBNVULAT4i+b18Ib/f3iI+b7E9WRJooMPG3huof+u
4J7p/pzPR1HSlaXTMvasa6bo9AM1RxlDwajBJk8bGMEFIRC8cspNjcqziQCPtrjPsKHIZyYTeqJV
7TNs1Yl4C5VKpUa+Pv6PxGRxcowC3UlDNURmoKP218g9WwZaqeONspcKVw/dh8ZLel0kaBRN2ia2
SK5o/Cyuq3QILBJFyvnvbUZx7vkSHPFi0Ek+5tZZTRgmkKgNHawDoAnEHiIc65Zqtm78xBesSlHl
s8+VaE/RiSAs4W5On1qiqmm1ngdyKJN8yOuvQKqOGPV7Q+41UgXTv2EuJkwISh9Q6QBLKamnkOjP
DKfTrGwvymipYc7Ow7++gjm0fTH21PEVJORs5wekK+b1ymC/KTn34vzLKTY7lYKadQq9hr1ru5JD
o3VchTFCuqp6lOWQGCJOAJeyTEqS3yk4duJRB9xYjRW40PviJbfQTw7fbAM+6x2R0nE4LUBEc4cZ
iniqatMGPQeiMt9z1dWXb2AZ6HoiOvmNz5TCFUCSkJD5hEj39+8TUmweWqleMevWFfKL1JqcAn/I
e2qVLZmMbleo5e8j3+hkQHBgDl8Ko6FAuPgPMkSJ5F20FFeseZEciHxB5t/+yFdkry+1JC3mFiZH
4NmxxuxAkZMr32BBR1gbAC2jp/s2teQkZ2b7Mul11MktGH7ryCCHChxTV551vJe75VStzKIxBzRJ
R8w7h+QEp3dF3w+AVXRtWN5TgI7jKySSFK0bPGMBWJfTOH5AVqq1y3nHJKqhfjqePon0lvOk/Dln
cMxaAaYWFKz94pWVgAhog0jC2ASMQhxO2SihONN8g/SbROepQ38sIEFaZv/lR4jkSfKcyuBZuOt4
FX7ZJ6Ns4/Kcvp5HrgYQ3T4DeHFGLlTy4EtaAK2dmzvMejK1g+Djcjy6EFTQNA+SpJsJ71Tr+5G+
z46iDGgVC56SOp6Mrc9MYeZuL5+XXW1bh6UHuwNzPy7YCq8TsWmIedVmHofn9HyS4vSe1tzUoTFD
FFWe2MW/+OOofhD4XBZEgfitQgujeQjQvvv6K2CvB8+moAagpZQGTyXmDzyDXSiWx71Qon+lKlrT
LSHUxEDbx/zwABF8x0avta8fGtqG8VUM4Ujh0uQawlGqXjq6izgIg/KZJ/pi/MNky9i5cj9AURmO
Rj9o0JPCF7VdHc3YSvzdUFT5z1fwDUrylGFPdSzSaYO/cXMhLZ3CHux2NIy7FBvaXsY3VvgW9WgR
zIItdsaz0aw0no4dyBWw5xesk/67ek0NFZWZxFazCDpWPFWMuGUBJiS3K7craSrLj8JHiRIDV1PH
GKrGP2nrMB1/Je6MMjwoqwhGq/V5VIUWO08WNcxQLVemsxkLj61O3FLmZq0VUlnsnyOHKyjdLtGq
FQkV+U7DyolSB7hPFGhPsajk1EiPTXhJBQmXlWkPfbscivG8n1iEdex+7rhYPCYlyuTOHBLeypa2
bShS8Erzl5DtS6RMUXia0TJcegKZFRr1MiTsgak+k+xxLUUhle3QKXJNUewDImasknA294B7iaaM
zN8DTAcyxHbt3X5/E3Q+xZqfUULBOeGQtsay5U5OtZNmH4dn8jnq2s9m9TL04IEBFWsQTCN+IYlM
yXcEPomieLuMs5pxDa0CFltgoNDHWEstRb7HRKo+bbdSz0L/1XMMHdwpckj6/Q48p2gDqU2u0+zV
ADGKPgsIhD0scswp6nBVRqq8jCe3uYxu7dUeZWHv8NVrWQWu+rVTc+mx50ht4ivixaGahhQaB4en
Ti/ydyCkQQEFwzSZrOLNJbzxXKN2dLpN0zdEle1BR8NjUZcOxYugxn/Hn8G/HsxGjKDazsOPhgj4
yWrO9Q03V2ESt985Icvs1IjZb5BSxxnodKbPs+XWgCWodWVfkHokmhkdRl0QP9usD3k0g3ptBOPC
Wr6st4AaLs4mPQqvXdCrQyBnjbWVGWhx0QB1eTa4F4L39K7Zw9s0oByLC5bn8AycfUvn0jKR9fhy
3QTJK/z9NYlOx62Dga9k15ZSvrGRaVCTXWnqpfd5wgPPhCBoK8BcutUrCsP428sErSgBOIlXMKWg
NGKuGyPR2NjduHExcpF1FtDAoZ0Fgcjv098kP8zPWp+kDJlIhb/aHLci42jqMNQLW+X1lnA3tmqA
iYhgTUtqpNJRrXhSTNbGHveD/U39w6u+l6UJMaYQDSpLyGTfkC7DhqZY8VEl4rOB2RIfCwEPv/FA
RZUDzNw5ZGuVisBc2hS7oHqv2uORlZOtBkuGK5XK+o5lvT7csz1QjxOJkNjerYCxyw49GExJ/Ph5
WRyO/nQjfXxHb8JEP/QuP3sZT3L/6iefKWCb0jbzFD7pXnjI+/IUTwZgNfhSbAolNUNmmjEchfEX
HlxJq1KEqRvYz6LkQujzR+qm0lfCVx7XwOf4JtAYiC67basdC4RNQMAGKdK7udM5oXcFMjuCUwU9
UbzDQAKGlydGdTTIQXno+FqgloJxsYXMBLkmI8mTfI42wyEoOsunbcfddlO3pOaQnnZHEdv2dc4B
ACvx+a5Sx5miWVWgRpYSOxkxr4twYKCwIt5SSSk6BbDIuE21iAZ53UJVFD8wMjRKQO4TVtD7MgqK
Dm4EXiANMiL6uJugvuTgH2EdZNIEC8PcB/LbBxQXCDy8lJxvYOfr+hC5+TIUqXh6tAZObWsB1d2n
aotUiz7Ez6sZ12cWuf4W/commCdZtJw59VU+R0XdQYG7EPlR33IktejzLQLS+rA1uhsDIe6nnzMt
WN5xp72u/oMuv5DrEgrCbYNKMJh/JY64LI1wkTGnqiv3uBCGJA7l7OwHw9kKL+8O1r7uwgX2aKbM
MitflVmFrHCNhRbtxbutWSLKzbjvpJdk0LQXR/iOsP8mqnSbYw6GbsmPSZ/sxbu/+tYdxpkkIhLW
vZ6W/0UaJAQirbrpLZNPmGWgLczL2RweL3c2iq8WIgDOmj1sbxwNSc+WrpbV9iJh0QUqM9DNmalH
MxA/WYKnkL8eJSCAv53LgE9Kh80fkfuVe1FfiqojP1bUHB4iTsSipZwzYP+0JrtKjGRFLEXUw/DK
/Vl4KGTIf0dxNaOWFeyS1+eA6qodzPEroyvXkK1ugH2mZvA4oJ4p0QhE7kIP6My7n7r2rAQuElkh
3jEG+hgqzfQGCYASDzpy5y85tHpyUcHftLQ/DNlq/WxYa6PvcZFBzZMssgrtWkajS5wBLIQZBwl9
2Q76Y1uKbRhTU4mLQ6Bsy1IxLGhYqLv9VG2uHyertp/NrOMuOVp5o0eHO4pmZq8eV0pr8m0hjeBu
w9/UVNLOYwKv270I960xjiYiTbXh/THsOWbZbt9kJaS4HczgxOBv7DH5C1rRUZa951MIBhTgFVoi
hSefCUx7ZNJHdhNVFsWg9xgi94nJFtNuF6anfKm/gjCn35cAwIpgtUxGhPFKzLqs5aHSQw+cBexW
d2r+Hq29eHIP0GXrS7w6bWN0Azi34Qtvh89ZP+4v3HmPY/1y/5r2NH1BKucvdrfQHmppZLsJ2GL1
WfdDDEBN6+8KIbYxrIHHdlsSivjNQGkvX6XdBlzeZXkeb8nv7rX5mX4Ow7oIzcFOWr8XZMu8M/jw
kS3FGMrwsWIG8v9AB+53ts7KFDeO4Uixw7w0TRWQHby8HnHQF93+/qoq+Y8QM7BuH3DSU7pzThAw
wODilRJLmzd4mzbSA8pkLdpWJMt2NK9dXzozvewEwXm2PuiAzDcG5/GZ66NWUJEnr9IlGJz4D93+
Zq619YQ6Zc6FDmPPzCy4I0xc+HHs9WHBRI3g+z7Z9C10NqfgkoS3d7ENa8KoE2vdnWUi26j26iQd
xcD4I2afRmWRtRxPTzFEfofWX2k+ezGs0TClWqvhFqYxJ6lTe9cbfDrFawnL/Hd7gQNk0zIAshEW
qHxjVF0rxsAXrkc8ZLEKoJhurjoBdPKBwnbOwsCfzdZ5vmLS0ACLy2Uj6nEQGIpesxAT2oSl20mQ
KzcFTdFabjomtZhKFMiYYIxknBhlGf1wiy3qZwgCEqoupWhLFu6ZKkvaRrbgyWTCs3l+w/v5Vr9K
1aKqBkfJSc1nMQizyjnnLgtpQERuHYzG9cLoaQNNKgqxemZpn+XqL+v9Y7WnVz4FjPkZtAyXhffU
jfmYpICEqclAQkWHc9Ko3IE8BA5MX4qFAvHz9+AmqHTcmh54PlXeK2VTvJwwJ1dFzHDYc3O45AYy
RVGUon2SXLeo3Ei6fGlFb3aXyrP8XQXdCMWx141fYJd7x/eb3PpoNT6rYVVlshBhD/x/hHgWa90x
zk6v3APxA3Gy8Zs6wOjM5Ia7uReV4dksw4gqN6wmKPAMyfgylwANvIdvE8plXF7CtPnQfX80xr7w
ynEvCVau7VSeQVKKV528X8SQQACGJ173lbgOUatOQfzNik2IACYYUG4DrVE5UbYfNWCkbb45n1sR
Ne1E2RAZPHPgBO4l2xlheSZ1tI5b1++4jA308u7KgGML8o3E0/2PPwtiIyFHX9hCE1ALzDmXlQLX
JWdxXZ5HdgajBSSnSONAzboS7i4FwMZ1SNKetKIHtLqjAedn87DVq3YIbiuZBjGNLUiOQFM5p69o
mLuYGoZgnBvCYZ73+HmSGNfbsQKd7l8AzzdlI4cEoOvXDKL8O1HFYeP3QUr6QJb9qtc9hkIV/zN3
Fngrm9FW0CgNlkhwg7k5qDo7e5knkiY6NGZoQktQts4BhWLodRtIiqSXuhBN9y3+aGLLAcZ4CqsM
auIgjK0IXejLY0RsMNg20AUrH50H6CQZDJcDICdffdYzTuXzhkVkMi2vJsbnjCJzscf2DVYUW+E9
QPgaWXK6cPrQCe1nuHf/2FUL3ATHbjJ/gkbaa2oKO/+gAGN8DFe4FxYBXeUFEa9rARdrMwfeMahQ
GcrGeONEpAf7DodZGwIrdFeqzpWY6uv79qzdsDP7SHB/Fwa04xRsKh7nwgQd9D+PQZTIS0JBswFi
sn47ufTMqgZPZ0RPN/huqDDSY0HZ/J76flviuYAkuVeuk1ekm31UGwXln1FN8RveuSaCSOHEfpM7
8c3XEG4AlTnWMPWeUAqZuTb1na7/z2wy3E151tlzp1GJmSXzB5N/wLU/Vb8iXz87NQAWlj7hjtCW
leFIDvm/LQcGTgT0Z4w62/q2tqTboRaINEe1bp986gvItSY4FJCdS0VWRJeS0jHrLaJ3+1RcTKQ0
Vfeh/f0Fg8FXwmLc3sUWqDKXmDQCO8To9jq2BkMHyjJbbQYE74hODs9GXr6dLRwCtmiCqjPzAlye
rXdbGBLJI2PeysXE0DCG+RHMrWcJ3G5RIwl5ndB8QMriyblZNUJFJ029Xqd6whNdRPgS+sLsN2q0
RPUMY3MGWQHhMMMtYthlP6jo+W2deGOOVSP2yqHJkOjahv+DGGyMVd0B3U9p+D2oNTS4IAMnO4Lb
Xq/aBJJyqxVUxDPsz0J8bAGz7sgr8BUA4MMDneUAe9YVIawY2qMunQSwH+t370g/9FEg3LtoDaeg
GlyrcaZZfzDhj/wgtuyp05afnllH+ytns157cSflyRJ6lXmzIrQzJtKQNyFJAb/S12Qc8HI+gxEE
xwkjrpbJ/jyYEnR+JOSWJng4hMsUwXFarDDR/AN6u3xMg75bLjzdr+hCKggRVl9nTWHANVzZ4uRq
+r6md1Srfw1YP5xix53xwzu47B9wsa/dRlthbQA11CIp/rRfs2niHj57+ER2chFZaMVyZLeDtocS
mzfJqzQgliaBHPpZPYFFbuue1Oj6E4c+Hhah6Cd0eI10cmjhIPZ3uRLXvYWr4vDnGcckPYowwoZG
b2HHkbg1WK5ZJo4IF0Gs1XQByisSVQPXjPmCDIJrO/BJ1fjtSQBciKGes1KdELTrXZovKpBGe9pE
uuR38JLFiCyW2nJBoxtisDkaEUa5qGmRxCJ5/BM2bF3mQcQ7WfWgbUhiw02YPaIVBbjj64B/I5Wt
B0lEBUXt7Ah5yeyrwMDi2bLDFs0MzXq6+/Y3Bj8VCTo27cRbDR1egrTjgditU6bmF07SCzRWZVp5
weAkX7BRFFxXDlDV+NI3Oy/GIx/Cpsum+WFmNmCtjGy+9zU8/CtR3XOlPI69S2aVER3WE2GQVTxX
5bvdGS4GM1Yb0iOLn63EfJ7umpJQOIG6mPd5hwXuiU2ivBznrWNefUYYhS7d1KoyNfW5vgSmQM9d
wRgmaFOjcaaoWADFYT/gKcwvxoCKDE7bjcrd+2ESeWuG891ZLIOpuh3gyrprbxIkMwPKgNYIZcT/
t8DKVVgFbYQDqJBuwGb2B7j68JrY0HodwFqycqujfi3tldiqeftzr/5QLukRbgWAY2CxgrhUnm+c
PlT4w5sNU3CmAjlqXKtoMDQKvo0oNK7pZcGA0bCNgYYEK3Zguhn1yIz11yTGqbUpvfktKZnwfR0Z
smIf+0ePlR3IdCZ0q81DARph1SeOhBzD+70lK11c/Oru9+sk7nG5O3913l552PhAPDIUVUNNMvAZ
XwIoKZN7qF1TY5CCNCcF+KZ+CINUh4e3rLTxy9fiZsf/5XwyLuzPufjHigav8S9IBDa+UyM2aekM
IqO7S8tOHuZHSBkC9/49lYMOkX6OmJze4GZdCd0EhatKwhGxkSTYOI0Wrf3nmvMyt5dX5YjQBCre
/UGFmmp/1NHstZE67AB/dwdbt3YZqObRj4wU4+EtidIiYzYpm0XWfPKpULEwBQTCO4Fy904RwXIR
oyCGbgvWSAXnFyW44ltCOM6NbUbTloToEB3WDALphSfCv3A6LqGsGVqiguoE1rNAVzr3APmqAQVi
AU8tNRhIIiEodyIGI5979YaPF7/ujg1X3txuK2A1/3iodOC+5oHhhCsi1t/9fwQl8r8epjCvbYtc
MmVkc8oT27LAYwPcru9EaPfT3/gKjOy2YkpLAPVe4p7Ss4wuE1kBgcFfkID8rUS9cKtJE+42AYuf
2cMWUVGAp2w8Vuo3AASYcw9CsjBEPa202UUXDt32SsPmTpt+2LbrHIVvKSZy9f2ukLXSHnCYoJ0S
0XIY2Oa5hDU/fiDbApTVQ1I0O3E3e4mYfcP0tk6+zMipdeNXhTGsApTTXcXWgh3bN6Cg99XpDzyg
9DfxYoCA0buEqV8++RU1+Pn7hF4tpw/CzY5DiTarUfC6an8SCGaEfY0k4bs0rnisEfR6r8SUuyg5
nfOcRmlaSuJdFdoxcxeL6ebpLQ+uqm6QBgUpIy+TUsd0o4wR+xd3iYdqZaH1EzC2iwyK0qtH4jBn
+8Djt5hfN5VeVK/RqRsD7dvrrY/J0MxkIs4Ivl73WT8Ki8jOgMh9vgzY0e2ao9rF0AS8/+PGnE7w
dBCMKDNpxx6BWYGrvegmTMiZGwx8pP38kVeL3crFFtqQ/2p7cpsTwQuKE1fy5322Ke5OdOGBhN1K
5jSBeqYD+KZ6XA+ICmLD3mwe3eQq7Hsc0Jn8MMM28jkGCGLGDwra1RFgvrzjWib+N/w2eRBP1ZK6
+3jXgU5pcBr59S4C+B6tDK7yLsWikPWvjk4a074qQmxsRVx5hzOahY8/PWKzYYLlI9svxWMoclC+
o1eLSk7hdRnuXfN57grId4ujfswnQLm/ot8iv3i8z2adV1m4n0AlmzHDuZn3alMXRem3bPxeEyNA
4RY+VESjUBCNW3V6sSSrsHsq96YlYcDU9WpiIqgYnvLnysp/xvHdXpprx2wXEGvYWKW89+PESUBk
qUbz5J/U1jnvB3G8Sq4OEpDBL0WkVreltshf90feemsZnGCwxQ5mAZa1pTgQaLfxnUYjxB9z1TSX
PixruOpHdN41Bv8QiNS5/hdGx6TY08Vu/1NSAt+rjqytggeE5+4LvP/Z7t49ay7yXnxaja0Mu6lH
/zkU6SXieyVCguaqAuonyrD8S3jzy6lGu0JrJl5ewKbiitMfbLX1lR0SuEH0k8qfmV6rRFDsYF8F
8895KqbIdIgVVLXDncL/rz2f/9S8WHy98hzu7dy1cls2LOAWt59oy+YuiD35mpwmzTvmH2LfGVN+
Vaot9biWRJg1lvnCHFsJ9nsJlPwbOE3H6Ca08BTybTG1LljUBvCkv/FZ1bGneLWXhuBMX7RWT5j3
bYLHS9Hp31RAJefRDIy7cEbS9OfLljSSvbH8BbDTfToN1kqsvh55uq1AtFqwdczVrlZ1FuTWYrAI
tpEuOal4MVUrzoFskHHG4p908TJrkTmsVbXoem/Auvw4fJTQ/92Pm7eXMbEplnQeyfX83up1o4Jj
lR0A2B6y6ZRWRkIMM3cahJFdbn195/FyLkGq+POFEb0UqrckdxTMAVd0DCSsdiky7Tbe3MBdZ4kU
KtiIat6OCljaRbNcMJ5Y/sWTl+YucYqqFf54wEgLWOtfuOqI/2IvTeFNbbLp+Pc2fHd7IbbktOer
rmMtzIYAgC5BLio+EjmfqpptJuFgYVHfytwFars5x6eiAn9vf13ODsjfp6y/yRzW6BXpsbVlIfzk
iMLj3iKjf25mMQ2gvVCiTIJduM3E0DGc0pAkqlQyRTsjh/owJsOW5BQS/NIBi36knxMQj8UUFAa8
cmYtzxQsEQArzM6AVUMtKaAFcifDs1DmOzffiYy5l7BerVPYd+ZZSzuNQ1h36U9hgZOHeQozV7WI
bw4J/kRxanMnuYTKPSV4v2T8IOIqdX4d1vQ5rGkN26aFInkjrX0VE1B98nYtRJ4Us0k9flJdsvIv
Cmi9NbFOB7RtSlJ/8TvhzZQnogWom2QRrifhAz8/qiK2UJbUla4a4iXSfjh2y2qqc0H5ue01Ky0U
sLhKaRZTLXL/QheT6vTtjja3CNSFq3+zCgw0ZrXGPGi3xqQ22Pt6BA8uebTN1nPV//nbCFOYM/h6
gs3dlKdVqT2jH6gksyd6ly6gVCoRg3sgMQ4DskHRHYTl1LsBj6SV5adR+/oGgpETdWjMbgO2A0Ec
geTfeGoDmHHtbXaGS0LxSdNLyNessvFKDjn4rNQbLAlE2jGkUV+V6qMxkPxTErk+XZOAbo/7UMBV
wodyE0ig3Bv1/6NATFageYrnVyh6ee0CZK2UoX0y5GCJW9G/nzVa9M8WcnSxneH7cQMRmJy0IPPS
8firLyf8uwLRb7XWnlYIJrrqWELjCW417YTLvcW4ahcHKNF3mXAVtR5dcIJkTYo1IaLKHJMdRqqe
+iIVQbRPw2RrjqTm74nx+G7G1Xnx1pryZ6zdmDQbyu+TbQ1ft3ah+8O6gyiub4IjB6s7HW6gEA6h
+qY0QRVlIaePye8V3pv5e1DlUKx2UjqJB52YLRQsmPr6wZaxMogWx9ILGQcUtR7tEc0ekzmdJycQ
E5o9LQzREAGxIAedePreF8P4il1ExK1h1wpwyc4bSfe4oKE0S7nyxjT9iakyVEV848ELyA8w/izj
aJjE2cyRFkVgOfy2wWDE64fJPwMKYa4WdkLccYSb/pqTLmmT1B2POXVZfOQl5xWcbk0gXFqlDT+s
7mFqWonbcXforCHTSSJKjmZBlZ3gFsY5xSPPedGzPKKa0Hi1FJust4XEFehFVjVzw7aQQCTGnhs4
IMehamTqM46+DfwjapT8pqmSD5IxGhdkpqYM/WukS8aNUv5nP4KjFsLCqnnEeFQJUhRgryJ4Xr06
z/YMMum19D6An37qvbcvdfKn7NTOvBfoLRrccdX2njkPTHDbc//1bBStdDPpyZiXhNl0/TkbHBaj
POA6Dfp1nrOCx6VhgvCCtuj9W804nLvh0YCDYHxjjqodySv5tFlCO1lToRYBYuPX9+eH0Jmow7iU
rN/5LCXKcwY3DoWWjpL8E5DE/C6wooXi5vRaxQ6CG3mFbk2fPJ81SO79yNKtBvY3NY9oKVLgUdBm
vb6UL5In7BrOT2cqoQ/h66HB5n5mMZXvkBOh3EHdIDU87eyEgQtfpycvND3xmM9LnabqC2TFjjSr
PtxCZtAyUHshaBLoOsKQ5lsj4+a7+WDik3SqQEBn/C+7JFRPque0dpYYZhpe5MFHFbtjd7wHv/HX
V0rxzvqw3/OMHE+vSVW1OtFpE0PHAAxw/3j40qcnTTvxriZ8D8oEMAPc5to8OOOBokLm0n4uvrtp
CON18YwcM4IeWDTarcAcyiXz+a2AYWgQdL8G1IJRct81wJgYC7rBQ5zJDWPSZM/iQo5Atw9Lw4GG
xQytS0tl4tdSfOclBLyUPFOSqW+HabCjypE4No29a0mD83GzxbCB8JYSViGySmY+h/jCbuyDxn9v
5v0Q/iiiyvPIBGOp/Jmmp16Tu4XYC44RCgrLU2TYqjcTa5WLaYdAK468keO6HvTrw/dou6KGSbnU
u/SLovXqNeGi4LZSn77othWAR9XFaoFNrhePEusDufR2IHpxY8NYCJJd7CuVN6KTXu9nPLJPSp32
aEJ7UYbLayjcvOpLTEnC9SfaJJzEpPt0rRWc7EPNvIEoU7VPYUx+bsTDUpRLmNXbZ/lcpzsvrgQ2
HAHQPQx45teeEJ8xVZ8Yuqi6H+ewVWs9n5ft1Z7mJT8TYYe18FscRsbTMQXP9LK4PLTOPOYSKdIi
QpSk3WZlb3I88R7n54SMd8vjqdIYjHZRvMc6hJduSMHIyJ1aAbStD40X/t336ul4dxEVtK6JOqlL
8GHra5bflqb/9hJJkOMPt+GY3Sw0RDDPCjSu3wpNSvTwZF2qdQCwy6zC1Xi8vfMDMf0FYhltQIbS
8fU1VnSIrcN0LNxIajqXefU+WEf6QMAhEvV1iXQD1nwhx3Je7KghwSq7649i52r1TvyE16O7oALj
dXXnYamDLEDTMvXPcKIqNp1Bgn3WSgUmJnWI972YnvYDkZhLCAFOsmRY+PBualBcUykbjJGAZx2x
eOaVCuEXPWIlYfQIS4poUMYc/ggU494R9eZ9rdkvTDqMopB8SE1V8niZybO+hV+ve2gkmCcCXWKm
M1FOer0+iLYXHq8gsRPvpxfIT55avphhzEH9GxY1B13y+DG9ExgBYjbIx4gO8AfIPkNker6FjHl+
ENijOV2YtxYKlEejfKIob+emiW6/VYxbfvMZdrkHR8U7H/ma+aede78/QNFWCnCJ/h9zJMH1lofn
cJfMaQScOS1toaS9ydNQY5prSFsQetdCU4vkykSKAqdfvG/8i0dvfSy9DVoJNdpaXdyZiET3sLyK
ui5T0BLMeE8uHqgmrQR5cfzCr/rEDV8SRQLQ9CXyOEY4K2WTqfPiF8QLBcXEevwevpQWtmqrimki
dIkArWWdfA+d8Wuc81xh77DCqFB/BzlpEUWNG1VZlfM5e9RbhQPBoELQpEvXZheZbVjnYsQVLnCC
TXySFACOSDocyoVPBsDXtyKDZ2KbzZtcaMjauHXrzcA0OlATkT940tAjdFIwLKNT8w/ld3NKfhT9
05pHt2q8kFPXQeqt02gFnIOHxWYv++NwSZxSN8dW0XdNoLggEf5pNW5WJU4T/+5A2JO/pH13x1l9
YfJA8zAJ72cFynNGRhv5FMCIMXKhe/WtAmqTEOBJB6sHuZTtm7TgqlW1dppRP4Y0naT82hJapC2U
pmr/7hhZeonT8muMmI761lACAJtYTrQZK4klO84xIAKU52QTn9Rl5OsPdkqrxW2B9TEDyaET68P9
0WkLwlBMPqsoE2rEHfQDseCK8i2mB1mB2nYaczY7bpHf0X2VrYKfs+jbew0wjD9B1KV3U1M/8Bh5
+X48WqV4ouiRSeaPuUpVcmMtsXGdldJoMFgYO6DS0pQb7HuUpFo6F0EGmBD7pKq++t6yn6IyFGa+
voBOKln6528i82QwSNX/34vbl23/tLt3XZQsQnl3gV5MYRi/oQ3HI/BiIcTBluQsrq1h53RYABSU
DmmUdEn9SstuH2TaQppc4MCHXbsFE4lXhNi899+UnsWPGGZB3aOczjBXOfSwmjXC3f0MtFD0kuK+
FRwPoEckRLwwTWQpfAcX8nBhkChgorrcexQ6a0RBs2TKqn+rcTb4xgXU9/0316/nw9KU/EwMLfa+
o1ZHlJ4jFSFzJiHMcbhDL4ywBprK6WIlOYqH24S0xwK620WjVaK9PUrbkhvNriJuKw0ZFu401Kfc
YKDrkhUNZXctdXVyPCMrFFZBuUr9M9Jk7E7qOjaA8IXeAv7Maw+acaHaVN0XTWrpoVaCeurw/NXV
O/5b0pY8RD5UstItYUhA/zbEhYIwG7leOhsU2eZUo7LzK3hXeVjSw2FtWdNU3YgPNiOUpTJneh1l
iJ028SqE4M52NxvO7vuaEjH4xTrvs6cHLwGKJ5mQmM6LXEwCWw+RnXA2RE6hBxp3RGHQ+QXUyGFr
2CDyY+CNFmPsPPJwRyrhUNLhX5J8MXvpYg51ZJzzFenqAQ2Xz2Bqgg13T1wyAy8WSFHDgCafPwkl
LJje2g6INYHpYV5Y48Ii/sP+/BGC7vtzekQ4LNMuPCQXcKTdwZr1ESn64z6JRujMkrpObgnJQW4w
JTiTiuwzFdL4qsN7b92LAQhClxrdeiUdtz47imVq0h1jQnx18WYMgsz3DIOOp1GbFoDPJkKmjGGo
qrTPDm+Bv9qUtnr0HLi5N3kZVANJ4myn5fz41kVamCpOm9m44BsoZj0xGtkRWDiV17/3BDAhDQiY
25r64d5edEGI21t8HpVPrBjjaoMg0XuqvZEGth4hPNAp9r2nuBbEsz41mOiuyvWeHLqZcsNK+B3/
5JurwOFYMHzeVWzvskLlGEjK2nhKNlX+PjuNKwA8lES101RsumaY2/e0HpObugQgmI4dHt38KvYD
AGTUJ8aap5buN71YxpQqkxhjz7YjC1+dT1mNzsn38a8AhiMG3G8YXp+U3jEtPu4D2EANCR1n3an9
mmfzhf3rbOZ9eSjUTMWfOb3jqzhAkpx+A2qqjq6D6Fe1CnVcwS7xnCqM9EP/HtfRmN2PBOQ93KdX
nPwaMbo2dt5zyeJnV7cCcTK5yeA27NhkjNH+dbbAlgcoKmSZMT/5dI7MFsr/5RhHKPlKZqtsWoRm
95AJWMSZKglQ/tNXnr8nGMHg26lECAe4Fxylh5MIxyzTJpVjcjvvslLCcfyctj6x5EZIKrRz2GeA
2oXZ4dCDiPx97oJn/0L7fnsXwTBpk4uJYbY1TfQrJAoVyGn/ajLdvahgE0PE38bXvSyRMLgHjq8b
4PYEvrhPn+UPuYZ4Cl1BsI63ga9EKN36gCO7zxDNbFrshyuDoSq2Kgr+seUe1jbpMQ9vCmrbIEV3
Kzs278SchpG9N0SXgHvG2VJ6N5DuU3a8pUMqd05rJ2Tzhcctj7DvL4mGKg0Ltdxc2U3u5oDVxNMA
047JbREOvP7XvOis1kUitVCDnAZfL9xnCBKQfuhxph/ef1hlDxQZdPSgQOhF4zekogYIa+zn+DuD
cqLXB1VUB+PjUHO1T6CSmKDv+J4qnmFI2zdHr/y2kOvs2jg/RSM3TBb6E6KI1eLr4fXVkLnTxzgu
qG7DmZpKrJ/Mfzt24p9yiPZEVve3OgkXU+O23clE523uX7KHNuIToA5zplmuFmX0O5v3o0MPnW/i
/+tNtIW+bL82fJbWQjVu2wc6Gww5PkuEgOm9axqjFHKWrYQkCVNi053LJ3hlXt0Ijz2vzoJn1KWO
Mbf22alYqYkIv7Yfhizk6pcX/qTQmLrmh9DzbDCFyOEYjSMGlVEVKTpIk/LWFvpsFlP70CGtJmYP
Iv4ie/atwbI8k/tAbOWH/m8QowvJds22gz5EwpAqD++WQE+4qEIwVS44Mkx7X0BpzGogmx7WLbis
NwXBTb96epl8nsY7yJNrsJaG23sC4C+AA6WabHYiDj/hqibX7lwuI8s0d6+nXNBwKjqnw1Tya8VI
TZP0gBT//GtHfydbDIw2PQXsh71nY/S1cDA+bv0CMRxPtzEUOyXmgVnj5thhp5kSFfSTloD5/KuC
vOjZkBZa0b/QVwBpNpAMNYQZSGxitM6s8BBj1XCadCh+a16GB4rp0Bv6M6ZACvwZkr3WkdqJlp0U
FgzYWf0VgU/MVSA9rnq17oYxUbV9p5OXs7WMSyOLm5rwCLwhmiI7PmaDsSmBaBWdVFVBFSLX0lB3
qGEqMBeQGE1z3A/XK8y4vr291pEJBGrkk+IuWs8txhvY72lekW7g6Io9u6Gta6UN7FugpiZn8qrm
KqbAbeMv+HQZUMoi5sbKvwTqbMaDF+RsjQiuQ2A6XZswI79yS+O0T/xxC5y50xSdiLQ8+lTFrTUy
9fDR6zW0fkR3xkj2o3rwJjCQ9RjJ73RAKAWDMs4L48maBMn7wZuw4iEqotK7OXlyOV7EKs0s+0+V
+AxNyb9WLgEcOCGtLc8Xc0ybMb49Ni0w56SzJyNdRyMCXJNYg8apGlbBt1Vow3NU/b9qAeYt6uv3
ZwzjH6ZveYXUrtiVmj0GOANrP6Whcoay3YLodFfXGVeNMOoDaHhv+7S5d2A4Ku0kN6KmVTn8tuzc
Sc21PbavhQ+GEBVYxL0kkPu7S1OOQYN+re8JmVlkULK28GkMfGpgh00yJtjtZl5pzNWPpA7WM7MC
Uck0hOrJQIVlxg9mnXW5Mp9JFxxWzKNMKmXyyTIjV4E2/K7GTmmB8bAC3BVmlzEnHoeDOXGccBRh
EFyn202rsU6W1whKQ1znvlSVtCoPd4/h+KXa0bJ13pUuzfXvTDaz5M3G+3KVYtVC18rzRdr9p2ls
u986tQpvKD8TtSWh2iy0btGxfg/YTifCHeDLB5jhHeJx2UTvFC+DQST2os0++ngKWdGLOgvnc3fL
3VbhMMo3aC4r1f6XgHvhto2NC6e6QBqjE0Q2/IfIQf6XLSQIMsQYiT0sI/GVIOjKXLtv6wPvzIym
Q1l3N4fQcYE1w4eOmaPgMQBvkKtEoxogy3/3GUpYNUoxDBsdC+AMEcdDnJslTUwtxeH4A7rCovtM
+9znMsnYXmun7cni4NRV0Swivj6Zkqjqpvv5Ga4GmVo2jSh/9iZm6z65ON7UAhGOq8BrvTUKyfa9
G2nszYz5oEEn5qUFMXYZnWh56+bR5DNliMA7aWO2pLbZpBXPtLZ75FGvvaT63oRH9J0ROdxtUFZm
IOdSwvperBW4mb/PldPYCZsDqjd0HFGT/XdL9ksApohHmgV0mGe7UtMz1PsxXniFDL5zi8sNljwl
ZANqildVLqeFSR27xH7/Dk/EjeZvGJrMb5I1ugZRTy2dREYMX964OcyNTcAqxn3Vordff+S3XDfi
w0NNs1ML1aULW3E7QQfGRdwnrNdyhDIxkLPS1ZzZ+rHGBQhcf9oAYp2/4pu/45kdHyKTWf8dSQUj
pvSokzZfWxSOvABL/9XpFS+rDit7Q65n4uKMCEnCyp10SVLS+iyANrBoDyKJwbuuokVbk0CWw0Ai
7Uk4SR+KpBZiPbPKhKIVXlsKp6oBMN8f7gpld7163EM4DbkJS/lzaUgOMn4jWx6z6QFAOQ65qFYn
rHG0oPPxjVwCgTCwYF5nJePNXoq1ruQjQZbpknoQ5D3vF10cX7xDxkGMNBlj4g2xc4pbNnGhYD4T
g6D7HkRXxVtFmgEbVFqvPBGvQ0Z+JquyAJJ2+7cVdradsJz56t/fhF9NZjykRWNBgl2mofrYzBU2
1DEdkvez4AV4LIcrqRkITu/9ObIi3pscp1UEC0hSap1rr6BM3ljvK9CPW+uIkHeN6KAMmPGBLMj8
nP/dxNaBFdjiX11hVnzyjenEgDZTVmtj/nHCnZ9JfcJYPAsJjTI6bEsdAE4SLAXVi3r4TUu18BrY
+VjUxHy6OyFs2BR2+nAhR75vdSteJL+C/lvAQHWnCLxXsosuaUlG+jD+UxXJiaZTKUE5NjY6/fwD
z3H6sww6oYvoBxOGKBOnbAH27GLzjgeBAAVhkACSwYKrs0MS8yDm19twILsdvoBHgoTD8Hr6fb3g
uaJgQkLAp1d5AaZozsPTSax8BrN++it+L13JKhaPB9Q/7wz+tKQ30avzyJixpEcoZo4V2LU8/yGn
+Awj9TxN70aT9mVIltircI2PQNAJfqK53kzjBoFIgzNSZx+u19J5MdWdNNF/TYnjHcLDllOUqlMc
QEc1tReIW0RR01lQAkunqprVdedTdyaFiktPwsECcb27zniKH35m1I1jlAt2MWSDMtXPeV1iCzoI
kVWft5oASYbjL0/F2gRSE4z5uyfhdzAMAMExXB+/QFyWhCBbwMPfXLCUEHxP29cATKniJ103TSHY
CdFeNeXwtNEftEbhBNO2bwP3F3qnMhF7oRDG0u7cWCEQ3LEQmwBm4N3wvDQ5pX4paHPD5bn3BwET
JvVOQXnzLx9dgCE5Ym6+NRPDV4iHtzh8KpaKNY4ZjxtJdPpdDqJwHHUiw9/wP4HOm/d7lp8kjmFd
bQXPX2WclO9WKyUstoCu8D7n8M3uqgTKENAp0HH20D689k6svBOWq6gr/cIHYP1OD6W+vt4zc865
i77AyZDFHg3Hs94H9tpyHZntA0JiP97WuZsclyiCwgOk0BHkqOvEuZw7PGokRRUc5WVVORBH33kV
XGA5wQnYUNCZmVi2C0lhTPWcb7j1NOgWoRNAfTzjelG2GZRPDTiDfAn0l6jrNnfyYWRDoC5Z8NqO
PdYpumtfmvOIYnaIzcvHRrQOhA8yBVQTMVwrnWh8wLTOzjqlcrWk7aJwumI1GGKMl0EbEE8SVvH0
eBP4Bf3ONsfppEwqMZ8E/7A1rMpPUc09/j4yYhwSHppfS00SMGT+JcP7zPZC0kSVL9/OpEEyJgYG
pPI0DtY//dgzQiR+cUKt+EAWscacPlzCLoaaeqJgIYLHC6J+evr5AfqOhWfbpTRh26gOwrbHZ3BM
hpmOD469kjg0n2+CZuQB6HZwzxWjvnlTNRPZ2/hfwWaYBKaZd6/hHwRTKfwH1MXrS6RqMDHQRFw3
f3tQ6H8jDAvEGbMg/JNDnStEHFw9MEwA1cO+n2h7ulipouHxI/J0qOsAenmSFPxqJwFVNMRvl4TL
Qn4KmrBSHvRpUM83X6IEmSaj/mK49JrKFNjvjMiGKPoeWZXuRi0qUKv9tcbzWa2P/yMPlaS9a7ML
VKOlXUsIiDED1eDsiEMEQswuAPgPXQb7bwchSLM47SQkbW0q/jsVJRln4o2ZhaxPJExuB0zjdCsU
713COnfX83yQqI8u1RFUHjR8MYg0qfPemNFgt38rokTdiVi6ogw6G2pY0J5uEAAxcF31MMS06EIZ
JtaSyAI32B0auVKclfKp5rAztG6gxYzDL+oCUavnqaXmZipXNkNtaB5msosmC6D1IvL8XP78jRom
wUJDPc/EJXU5Q0SYV2QwZNNONGe1Z7svAuM4MdShUrIku0OdJli0I8T3BeGQjrHRz4+7PVLa6Sd8
1CQsE/zx22foyOz43BSPXxu293WvGdR39CZM9V4pL3qGrz8WKL/yMcREZW02a5dYFXiwuubUohBH
atl0+WDEti5P/Vsy5UKPffqIR4mtd+XBEIb4cK0mqXQAZJyVLUhzcx99ztZhIws0VTApEw2dNqPY
nWGIoJYy0cwxpc2zJzwQmgpH79eX7AbWWFdlcu/MqYcwACkfbuGdslvflRQfkoSqUhXLkVc4vN2/
Ojq9vRG5Hvf/GYab2ybYE4eU+ylsvXvtHcQ7prlEZa638H/ifM6BZpI25qVtNg2uLUn5NYuPL4dP
7Steu67q5fCA2Nss3KiRvCWnYRiCq8QtcgwVHImOKuzUiKXPOdUsjh7A3SsotxKJyhCVrVdo1Ojl
s7iYqmCj+rBYMYdoAr15ylIa6xTA/XrOyAr3EZcchJPiEu9wg43mD+2hji2qu+HQBEg7NVzLjcNr
HBFTcGNEan5RzomqB/zr+Wu8CdnnKZcY7JQHsLTRP+wEkCYEGOmYhuzc0A3Uyi7Y2JmMjK5X//KD
5ikQQEutN1w/yCkrL4VNJyfpDwFyHflnklIlDdq7Cd3Nee8LUC9q9d2v/kyDhmGHp5UYsgxJaq1O
XTJk4aXHj6GGfRNeZzKSHi4XZfviKOD7sAvx0SzEQ6xLbEaFsJ8GoExMNJEa3XpzSyuoqQ85vduf
BVmv+6kKNugAxUvvmwblrwfjJOndWiFkvnbNev+CITL1WGB9jg/MmDrzGyiBICmb4IbU2cXUDocO
5G7opFvpfMr5l2/q8R+9+l7T7vxxt5Wjbb5QIJtYFnyztjDcRhjNPSjk0snQtOBYrn66m0Jw4ucF
E344cRd1Mtszg/PEqhOIEiujkxo+Bz7T9WC0rNftsSP10519xmSef+jDYbJKApOiI4PDooaQHNMD
7W0zsVjoKdx/GBu3iH6i4uHu6d5GUIsRg/ATWFEq/jN/Qc1hgjajLJJJGUkCSt5zpctWcgCaAMUJ
bVUoQCuCvloqUuGMBhrpJ9/quliCT6VKu4/Hn2MyU0ZJIllhMTwwmas6zkbBValaekhwHJC3kQeL
i0hhf/9bJc7fRw4cV8oPfDRajRfgZ/f+AxCyfC3bFTYRLiy78sPOHWUCIyvBSPpj4tZwr4/1EyCX
R1padErtzEz2xIZ0652QHtoAhi9yISQvPzq3MA6c3AoDlYLvFUY1/mrcHhEFvdDuLg9ntPhAimOY
4CLZEnQajCQFHq+F5s9kJ+HgVhsb2pXnxXbeYYbbRSOP6gYdj8S1ZE2OQunct83OxqXs5HRekDfO
mWfsmQoqS6Mrpef3NAgNMcIrNzSxl4e7oibtuMsp8P+CJlWa7T1XaCiOGfTK/lJOxDyrofXlL6be
78NAox3sY/V0dkd0UFXH7Yfj/3TYa/BR1IARMe2R11meiwpC6v++ZjtRZfKrSSl7eojnmixbeUG5
+CoQFFznCKJ49gHcl4i1MT9SlFQ1vhsGQWTc/fCV1Og6iokHkPMcT9w/4Y1w1habGp8z5gH5KtLm
WsTPN8Dd9LzQz9NPLn1aucrsywtDJkUOaHi5tmw7lGE6XC3//G0jU0ggyIFbcpYQgHL/+TuChsSY
eyFJW++jW72M9BVwIp6BqxHC84Ei85c4mNq/GKV0rhS1YcxHT2u556nu1ug+8axbEJta9derhWZH
QX2e/ELZsnmtY7wdIqrPP+zLU+5wvIeHPLpaEPgTK165FX1+IHH948WUts1h5LvdVL8oFW+eBUR6
oVuqXuR4MQ7idOjwsivz/CZI9EttuW4B6G8u/Kg4fRWayijCQK5HOktV6AzWQX6WeZqrZzg/a/EY
UtLKTagA3UmbmQ5+T8MVanz4LqH1iBn/ckwvG5uexLeUM/dEjWEjOd9NJWmvVwI4oKWiXwlD/3yC
Nx0PwYNXCyNuVb8W8fdOJGyay+ZrPgnc7mXfp0iw85thLuTcZReBxaNMkmydC4Ajiqw1oXsxYIib
tN5RBwHAu+whBtKAwFfLGZ8Wsx8VR8juJ6mQvoB69NQINKvYyPUOPkF/jIlyfCCF6+baRZr5aYfp
2cTNJHCXahl3V12+PyeBw1fK+FDZV64PJ/vi7Rop06gAXdT6h8veqwY3e93wiZbZ59LjyKBkY0BX
kIL0yqUzo/CeI4Q5Tux4EFsvrHkAxuFqzC0qI2Wlk29buQKg9aQNPxR8rEYlm2T/LLVMZIh18uQd
Ro5WSsZS+h8/okcz8oPL5WKLJLSPmW6KHUsGmYxOpXCuOXIY9w+wb/00SgUCxHXDZldcm2GlMiXJ
Kh53SuJ29ga3XnItNem0tmkGzoZBpSqVgdoGNxfUkrUQOkdo/kB+nIR6U9Km9mG+0SMjfGE+2U12
bTFzkKnKKYyhKzOHjxZGmIhDjZhBUWi7qLzBN1xdTB/YM/eQOlx4VrlhBt2h1XzaSifgJLm08bDG
WAyINdt771Yhz0zC2myEruT3Skpv+szsdWXa6Rz/Ri/rxWt0zGG3stDkPetweO5h0cMkMo/Z5kx+
hCAZhJ1+VuUf240KFT45EmymvY07Yf+3HYv/1BK2ujGuNqVyLduZdOy3O99MS3WFbIRk4+TsKtrX
veYuUxj/e0M0BbSM1P3BerxhNJ8UdLZ9nJ373hL+ShGw16o0EHiIb8YhuS5qycrO5vyqjh8FWwWP
nwmMkqRdv4Uuv6MsFX/DcGzbmWN1KrsG/Qv+Q2YyFouDH/RVfwq9Zg37BEXxBzF1fPAb5KBtWMfx
aesPs7lZZI9WArNQ9leXIed8jfejS7aZahQ/IRnmSRD9JBJoiabcNRM6J9jZ6cehGnWQ0SUKZaqS
g/YjXmZq06oWHEaWRmLjCU7Lfb21xUVVKgRZVo47tAnDaMYmVYtYvsFmqzu9YWxQmbk9iUsQK5yh
IZkIKLNroYFmjVMXQfPJyeX6+O49+KFi2Gadg1sf2f4nnFDvT9HvpLAxxAKIDDT5sk7E8EnmodFJ
Ja4teB/krQBDgepCpj/+17atiHB1cjeiOU5uBFZV9qd4OyauWNXIFVS4RTQNpxIWOLJL6ouSBAWJ
wYewBXRAAwKF+xZj5qeOvmtGM4+MfMjYa+7pm9RNL7JQU+SZOM2g+/mJkbg6pydMpKAINTsWwpmr
hlJWcmVvAa/ZNYjn9h/VsPvgResYJbSE8xsHIqkrKAHpr6hqCfgW9tdUg3NeChG/DsewbpAuQ/qL
OXcc0ajhXsGm2No97E4ccHLT47SPvI3dIK3Y/MmUhbfX3qGKSkPccW3xkw9a0BlEj2LXcOEf/NcN
j+HUZHy1EfS8n/q4kSFkg01Snf0eVOyvKJuJDF+jweVFlWGe4Rlo0Fatab0tL707ucHMd5zJW84C
0xzn/2GeOneNfL5Am7F5HSRM9cABZU+lMD1WI5oComzLsWFYH9RjOJ7bximkaWSryRBpk+LbGrW8
3Mc6Nf0ufkq/cZbclQG9pZxerKUHiFKnm4SwvE6EvZqMYqOuaGj4rs1GVSH++bs4ouR3WniyNisf
uZkNV7Zy5o+U/TFFCfWVXbio7XsWkx2D3CZtwZb0ABRc0b7dnfN5O6XfGLTYX1M6rqgmUbh2XXLv
PR6+b1/6fYtNb7DfwD/mH3GewSiHbsusDcyK/2wGMqpGMnB5wl3tlq3Rinr+SBli5yVKthgVFDwZ
sICvyNk/2Wt1zPzlOVV7d92iDpKodfyRS5iy7Sd/ZzgWhY817F4PMrJPJ3l9NBJzjI1a1NX5se6r
geNtC9G1qXy0UCD9Eoc018eeO0/H8X650sPuRbTaHPi4NBHqIcsXYjLAKsb5awvi0kMwYENtNoxd
j3L8SazZ+edMTOpeuWXHP6cghtwlej4qs2F4uZTGM68Uyy2m/lJM7p8DUHd/ZxTSJL8iaHpLxjId
k5nqKiyiejojgcoVAg3u6G1Fy32lcJHRBpByZ51k4dDLbHVCpqZ+n9vkV9uyEtc54ME1e8SiBF9L
dlAxHFF5GYRR9bFVK722S1D2CTngv8Idsa259+kCc/jXehPokss33XetMlzUdNjsyHcP/9ZQSdhH
bmF9D/lI52sehtyW56zqQg84o+il/Qp6wAdqnSzvqx0r6lM1RflEgvUPUBYLYb3dNgs178D1kxd/
09q5A9sUsYwDshk44YTuU6zHjfchHNUX/2wEDPg4CJS8PU7SLL4tG/JhEk8/p+G11cI8fRNunXyF
YuXkzwCaTEnpuiRgIFSLZ2F7TEHFtRek8l7V0gGInIWLoGm1t3788zKQ+gIp4b4qsRhiPnU7cjE3
OOzgWuK9M6ThFT5niF1UvYvlph1XxKMsxB2TfL0OsZ3LVg34I2AaGO/Rde6+Urjb8jO+zvWSrS5q
v+gg5tUWRAMDcvxQbv8kfpwekdkpbg8E1ksFsDIfZmVea8RJ7u+Raz2XyozsG3hBqZJ1jDSiMeO+
VC/XnezZy1fXzK2r4/+Rzz0sqi91/IVSxPu6N1/6eg8OFpVuYGxpwNeJjhqAL6CzkDFeqBzEYZeK
V1iL49XvBYnx0qoWrGOaUrwo9zI7n860IDQ6ZUwFwRvTq3pdk0Gq1zIhFQ7Oj0qBqg4ulKByddhU
VWqL59nZOyH1DOKMhexhhxgkkalZJhmvfl7to2kB5LNWWKiIM9y+R4VmnCvazmST4WS87Ph48MoR
p9CzvzKcy+Pr2ObbK5NmqGtkqSMnDd6oxDsj18k83b1ckvMa2PtVnaHtcX5HfSUFzz4aT2UK/+PH
9EgAShyqZpQZAB1kpvUC7u4UzA/v65z7ysmTbYLlQgb50/4Gnkm7W5a/0p74Ut6BzI3b/GnEut+X
FaUNH9W6VNcvuNxvAUI3yXNSRsJr2ub+LBWwqZvzGp/FshXa/DXqatcECv1WCc3mSfM1tkZiuU/H
hIGsIgdIHWDmi8dESKg/I0kjEUhWbsejxKyiKvyn1xv+9aN4VmKU+7Njqz22nNofYqdi62nKGis0
dRYTYP2HImdVwB0AfkWDZ6/sMwv5mzCWVGQYt/v7XWaKWKOuGzUhb+b2PafXryq6KIlKkPLoKioi
rvpE+oXKk1VWL5sesLM/35sKZjcKVfS6H7UYylBb8pfbVf/QHfWoJSV5OeouGIzCIcBEvUVxb3iJ
vHA9yc2b6A3B+rXy3lA7VNG28SMDMJAP0DOp1lnGkCNpjtIK04GKWFt0O4jLObzwXlzaZLVGvzVt
GPeR2A/fXdEewc9okLiEAb57ypv5/CRwjMNiHJJU3CfDAe+/NG9XZws1TB922b15r0bKDCo+sU9K
GDW+ocG30G9SbuCvbZoYw0qbKWN1l54DvxwdPR0AL3PautbUMh0fiwoDC1iJ0E2eggNPeU6qAptx
KIDixYzs1QxHc1huOq0e/C5L+asOrUWL+5j0Rb38Wn/uxkuvs1Tw2fNNwelEOUzn5ciIOd2XeYlU
Q2Oq7vDlNfyTDtPs3TC2rD5DpDSTTuJ+GHPUkS/Nm5dEYcUg4m5W/AkF2tXTmrYz18MIbUGgkPgv
lOYcdKnm4ZqX69N1OW7FOuIOLAW5o0wT4Z9tVS0fcDTUK+HVGW6vlyVDBV3IgGoxmkzfrJN4Ts0G
1VKOO2KxTaohP6vR/CBDOJ3hnP62Q8x10gcmX1m55Dy3vIi+1qwviFacyF0D+QZIWs6ad9C6RULz
+4AmMW9JSjlW/+5Yi7usOv/gqj2uitXFSMfRwk2LQAyziKRb6avgaVNMEM8dqQFVXvKRwQdweVwf
tx/7o5XAOGylnPYWo2qV/gnExa0slmSIjJk6Tfftf+OSmBwkDLS0BgYon23Ngz/aQaB6BEdaBwC6
sSksz13hty/LZUQfPl8VKopv/MTvl0HuxDaqVWLxwVy8jmySsLHzECioRpvG7c3poYsVD0x0E6Te
EQ/RuUBxzpUSXVzmyFNAOnPG2Va56s5jwfXSKwYF6WnIM34pAp835Pd4r8QbK6iTZwBjpyAejQUx
h2j23KhIlOkI+M8/exYh22ygiFt+kRnpz+93Ue2PDcMivDwdXJVZWQeTaW9R46HEgPm48e3CTQdF
NtPw1JkVFBrrEfXNjuDR24gluMFwFWDqcdJ9bbO0c2dSrvtsO8v3G8chJtENcGfEJRWqH0V//IvM
awQyHeiWNTV+ovjQOornu5zJkQ5RyCCTjVa4utf747n1sDMoZBW0mgCw6tNQqx+th3r7EnbRQeS2
F/jzIzfBKtvZcmCYoG3e9RbnZ3LNPfZTioJJ7liMcPPan9qzZjOM5FpoWt+PctNi9L2vs2eb/j9K
u1ABDwo7vrvg1OhhdyJBLgLYSMOUhngzZDq/qOfr4xJiuw2gqPPzS2yrA8DkGlyN7FUx/zzdsdZE
akVgpoJAo2WWI4Olj79ST/roVfXf6CO3HDoIkBgQCTfU4GFu31sWHHdvUWhONui8WjLVtHD/x/Rb
1gzYH56FfMWtkO4FkWzQTGR7kDktcAMV0MixVKKpRBOkv/iJJfwsUQJwo9D84zuAkFCdHxGH8OlL
2ZZNMbDZZ5K5aBN0eY854P8gNDTfwVOdakVhPprJKG2AawkMcETAQbrWEWiM/5T68FCsBgOEQuYt
e4qG9136w/gfIG88Lgr6ogEIhEej7Ln7Uj+FXiCxL3AmVZdc068i/P9ddx8Q2HmbNHNL2TMeVK+X
iWf6V+8xsfEVHqZxIeG9qj0ehIbGfHfLSfi481aUhYEPSom7xG2rRl52NN2zLed1y2WRxKUP10ZI
AXvLXmNyrdtuln1+UDkhL0ltmRXSoX6XYWEtIe83XwLo6zis3ISW1wzzFV3j/vuzJwbXmDO0sGi6
L/xYBE12w9pcWKVu7pt9a5Ajgfr2wQE/OMXMo3dlKQOhcKWO5wHPf/4LF5+kgDPxpW15JuBojsLk
ie1AQvOMVrbEKNKWqnmq5v+G5yKOqMH3ebzH6ARarlWnNNEVReeaCKrU1LmVe25xR2ptzwsXHXpH
NhQu/RkZdL6JFA1m9qeqbs35vMxbCynrP6i2qEbK8yECJVVObvku1Dcft9sSWj5WUArv3RPeaMqg
x57EQahCEBu0Q2OvHryxr47gBlXQvZ6o1z9VNfR1WCwjE6E+gS1ZJgyAI0izzG61DM6yUiFgVzrS
HFsw60TbfVJIYBxomgGHQbzV9dwgnYN1Xqmx3OL1sGUL4AJzc0zh7Jeqg7OljdpAVTffT/J5ljME
PD+m9YGOHqE4/btjWXSDWanDEadBlJnw0iyGNzSSinBp0bcILf23+uvMzKBPXhUt7LDpag/WxbhX
6AWYgTCBwJV0cZngi+Rdl5JNZ0He6zkPUqNntkMJ9nf3/z1+O/epdPK2X0Qaiym66zO0V8otFySD
PJBkJs5doxT4p2zIxQngqOdHmKq4hWcVZq1zeVZQ8SNeO2XfgoEDWcUBdgHkvQlB2SRQKfZo5wuv
1cu1f/D2x+Kom5i+O2D3o0s5B9pDz0IbKfzDgkYiIY8Tv6MQTiqAAjOy3jM7PxF+hGrbGc6ntlgP
DmFqNZqf+xfcc+QWPlhod4BM8+Mkj9OMiQu+bHR4OifsILnvXzdQT6ambMvO8n0kURkPEMqzgpE1
FltsAVgc+V4Tuw/MS+ck31ha5Pm7js47N7YllsJGre/BFLxz3bko00a4JfY63+SRySss55OV+WuZ
AiYApQaObXy8IfKmoGlQ3KKDVL2A4pDey5uZtpL1F/dqGOBZgXR3t4p9m5JcTj1f3l+6kzxDFWKP
Bg32kVykNLWvdkLEn/UDfGmJYLMQXSWDZy76tzXsR4pA4/JhEdUpBJPEjwn6B7NezDwVZfmVzTys
jxHK8ZgXLhKttXrtTCX0Rf3WBSxikTL/Vsz9OfLzjW9CFQuj5oNx7/7Lw4uBd7fi8nPrCF0PBDgX
ydauRwK2EAMHuwANyccy3M4oteJ20vmx5oK2lpyat18C8u9GhnhrmUMk22+82f9gsKHsCh14DxY1
I7X6V/9gJAv3oQ2PY/2RJbryWkBGEghwmx9h+Ia/fqIrYJdUsiYlMJXr1hAQKpQJR6aEVAdyc9Gf
ae5mWNwz3Nq8iaajuX+hM2x9syLxabbxX1usTZSUVGIyhuS92Ap6NPyQOqH0BGQG0QqIIoavOyZP
x2B1XDhGHTaBcJBqBtPCY1ghNvnJ7KaaIeFO1YahjzJyQCnjS2lXeNgQEmCTVHlkh/kJPHDYP2rb
SRr5sbOguapFW9uTck+UIWkQJ9Ykc9prktu9YfsOtbtoazqN4lTR7FjZ+fw1G+ZjNPYIXQoOhciq
qlEqjzTfuzl/Vd7O57WTb6nh76lGsj+p8miX8L20vZB40/Hir12KquNtoMoe4Isk6v60Yf9bP+8T
2CDQhFbvPtJGRCbx0oQuJtix8ZBwFtMZ4KiQ9MNU8gO8NS9xVge6lCCdBenUE08PIC5d2CF1wmiP
DFAve8cY4h92OvoFXzX1yTmdiIU7UR+WM0KYsqhW4+VRAPnAwrnOLoWnPmHyGP8hlhJbu3Ox3f4W
WDkVlp9tsSPWVtUkGGdz4o2oJh3d16eOu8KuTVJK8kdb1+qWRq3yDvkaK2kvt+jCtiL5s3NvLGNt
EUrDlwaZtGDqm4CJbHCCvGsux4SmgBsN2R/P2mLIB+O2blLwqugs1aKrfUe6UCwhDal1mEuVZ0dx
sojJZBIGjEVxMq/PZx+CNh/t2gVnnkmZQq78F620og/DbAOXPI1Mu/qKA7K9NxCPC6klL3xuWCq5
tZsICbBsiCqmrrhVz6EgC6+/H3r9JaEEPZVCpIrDAVvYkUnMlQKm7YoekQe5McfnYYCrV6KhpMgv
ikxAE4666gxvkKPG3wEUHANU/Iln+oa2B8bDHG3I9AiAPRSenl0OQr+rGdHacLSb1Ycva5/YHXZh
nBaZlgQZ46hcqsu5DsLDSQrr64UoPp+5cHz2HNT40jR7PWn+HVCTSzMZvxKN2PKnroft/eSN90wS
eg/WhZukjOpE8smtn0UcyU4FaUctpEcG6HT4AlVpZVlpSOktQH6BSGTGgIc1wTFF7uw6zdQ3Ah9h
lGYvQv53xjz7WBDk54be98McDFUMfhu/Zsf+X2EhbQvxU/U+u0ZA7SZmJCEQjTcP/qpJeBaqNKIp
bCTrc4QrgjWMY1Nx4HUKPn7XubPxnXnDN84MB64yqF7wA9xqdShlLsVA8JqcblP5VBSUeR5wwzsT
UTNhS3LwCJokrjRocp3nEDoyVMi8tLs/5nMrEGl6quVufDDqN+Gez4YMOurBXK8Iirapw4yFSM+H
35Yx6MZVJd3i6ri790P+hYPtV1tOkBI4wt53EB5VpneG3k3CoXDPA8T4XGMC7mhY0XUuatGHSXwY
nIs9AIr5DN9E2L+VsjQ9WyWYK6h76OigtxbuwomUyp1DrTknRnfShMM5sgtyvcPfMhiEnXU6UUzm
EFVelPZEPO43YPtEXbMMz+vO/sveyGzL4JWR5ep0MSuedFWvATjmyyvEeQshcOQW75p4gWJyqi5O
HblD/xPGl1t6sbs5NCtJRr2MPeSLzeUmExzvb2z0+ZK2CqDAky1rumWBvcSao1KDU+oiJ39uNrYf
oC5OPMeOO/s+TRsnRL22C21PPbWDBT++MXgIyQFwUEYLXbpKf1uIbjItjB3x8bw+n/CKqgJqUVCE
xWdOGV9vdBloYMClwIo4s8jFDyF61bs8qwqjD+aSp44QprSWtyoHDfyXWQAkDe8Y7VzzCQZ9zkZQ
1wz2Lan4hoYWvtl8S6mJh8I19oqqgLALkXIEVLXXNHg2Ub3Dt9HcHzgBMOrXVjbZ3fBFoAKXT5gk
LmCSFNF0OqNzwzJEL7wqKHMsbqI3t46ivTzEaDWBd5zcvRf03+RJJnfvFLkPmWE0fAMz1x8HGZUS
vUgu+P1el+nLbG6Z0OhknClXvzlmLr70MUdPD5Ke12QIGaTHyTw4T7t2w7iiJ+z52vr+Tl8DWSgz
tim38he9imuK+hmY/BKHg+6Wo6i1OQt6R2T94PLqqIgUqxWSFC5afk079h9rIPbBYijnekJKgXIa
pAEWyz9l3o7luqKy1TtvPJTHLEUXQv25TqYr7+Op7fdYLf1rTo+Q4WydGbcWbD9hmg263Pl/NaxC
Q1eh7uZ5JHntK41P2fzf2McHkEz3KQzfH75sQ3Gr01IunsYPWqNhL9fooS4prin0oe5ThN9o4fQA
vV8Nx2MWznH8c3F2OqfnRAMCQ8lUMkBSIxEjVcbORx8NmrKQ5em0ARTzBB+EzMFIbJFPA3kS1x0l
undK86Iba2Z7Rv4fdRgdvPaHpq9A6TeIEz5zWs2ucOAAqMG8qBadTzTdnelBSFYpgomCAM+qDnSt
VVctky7WHRyGoBHebCIQSe/VfwSwV5NkoObg325V84P5KzQXP9DzqSmDKbbkQUswC2T9+ZAVs3+4
WJJb3kwY/S5CSSu6a3lYB5s6AtABrOmDUhGCPGasoDtNy8sTOUsa+8bYRwPqRJRkgJJH9ml0v1ge
GXTFG5NlI9NwRXpG8l78lOa0iWuoFl7NatZ8xUv3OwDN3a/Hi3fwS5svr3A4OGI9yzehCCs8LwUT
Rft0bZg+haUcXraxdMZ2Si22MHD4OtIi4ikiv1SiE93I5durLvk2D1rKO0Vq5E6mS8xs+8fMPO0Y
p4YWJqjAFYwCuQofZR661tcyL50O9ZCuovlUu7mDgWmPRU5u51/zcIfnIk1KSfSp4j82cm3fRdBs
ROIblyKVQ6kM+gRE0iDixdS492FmMz64JtlLVbWEf2fO/1MwgOWss/fm9jNnAhdM5WWNRLAQYnxc
9EjZiAB/GMw7FpjatbIUPs9mvSibySOXqBld4AicOL4dVJrGIZXbnQq6QIf46Ao13EzAdrUT0Q6D
oKP1JPqVBNLfBA4clV8XZfqjGTc9f0P6WEVkQFOFSQpqGDUgzkGzbPS5z7cc40KRDP1o/TvtvPjn
98fiOSsqYiFiiJXnHV32V+oPoC0AoZoXqih99G4/Us28l5f0Qc4LRuQxeXbLIAg0RwEYlmjWpAtB
C2G2+39I2+2wuOxBQQcreRi1W+FYRFKP7poLAOhdQJ0WfHMRFddMeAezAFtacE8L0t65TqYxmb+L
vr4nl0W0kpUkAIO3S48Dg+AedfPN9Kjnv8pF0apfD9t+N4ZEPhPdxOVnXDi1/otvP6sWFYfmJkgd
i3Z9S0y6x1pY23Zx8temgI3x8+02qS+nbSOQyfzpqqbhLwmDGr2JQ3E8az/gt3jCpaT4ubHQEzlk
r1H7JGNsp967XVti4Ui1EbE8RYbsGo4PuLG2nt4/OEO4cCHJ4cHkHknF09Uolz39Dfytj8547y01
6IOh5TflyCJNPIndiyI8ZRfhmkC/Z1uPpf4DZD4q0ciTWwydzkWIdxbJBLd2B5Qtumf+iU+fEzhD
+i+5Z/Y9TNZaO6oENOmGq0dRPIVFo/eM0Bynl0lHsqS+xaBcEMnKtD8Y80qj7oUnmc4TshAYkXW+
gq4cQ4AxDHfTAG7VAASmd1Izo1nWYjo68KeyuarQ9658wWbAKoT3UvxzQ0/HIcCr5HZUG6Vi4kIc
LhNmim/ZRUkc/2h/iNcJDsGBbQrQIb3owgzcjiAWRDi5uDgX702VocRpW+tGgyudj3WVPn7beV79
j8VJ3kdf/BWfCoYTgTTEvzB+lmzdg5pYw2dZ8N4YgzrhumA4nrYXQWHmwxG5JBF9UtOD3TyESXPz
0yNvgNjsn+oiAtbrqrU1k8VQ5bz7rOXAZZzRw1ayULPWtho9eNDnAs+qhZ5Kuxaq3feXzUu7zDXE
QgsTg9UtrKUSO8/7cwR5hbFlfQ40Wi+XU0VAwr74iArJr5y4tjx/+LkopsnxzapOPwYbqkyZdT3c
KdzDeZg8ErNC9Ri4MeNUlMCsTvJIvJq/Zs62ywqxeE2UHBrffuA//S43Od93rXJUNV1HhuuaYSkq
A3UqEPyMrodzmyFhZd8SXjm11YjwB5mFVLcBbvEWCfgvCKUdXnMkKUeOI+DP28xS7qGEqoHHHs8t
UrO3V6FIstup82+LEIwNjJVGXG0ZTY36PnB80Ag6KeJTcnlltLKH+oooBtnZAOXcWiKYwDBL9X/S
LIb8TtQaMh6C0poyGXQR8WubtACb/inKAfoIQWDagnaisHQWXacW7Mh7y1qDGILtzrBk9god0pPp
knTGCa8BVqWJjpWrMhds4bWR2432/NsNf8Jq0KxJvERPrJoCBQ1vLbaNs/pqW2b3JHxvPAZiGKY9
iZlUpiRtLnNOPCQZEkMu4CUjBG79VQw+PWjw59Cgq4fLq8rTbmmR1n+5DYnSRbqF89I1eiAVnERC
DJsEijNAawAwkVwNqqFU8HiSn87h3nHQQETJSwJuSypUYTRh3lwPbUAC/MhikMKK/3dt7rhXYN3B
XSz3CL8nEj7ytvCBzTY5MWo0EukZRSX4Ds9vMPEivFp7TK6Mq19VZH4dxX47ROYe9IsUbewKkzEZ
aghhs51szsINvDMgE56Yuv1c2H8TnTwt596+Y4JvJ3KSZkANr3SIytJb3S6na/FBlNuY4FdIHjep
4cTmylZ02QgAldTE5GuY2Gn4ZQkNN/yzIraEE0JDcnFO9l1Iu0aToQGBUK+5T1AFFFR4lJ3m61yJ
kXPzJt50kJql5v3WFBBjNpOm+tE2koScw4wWU0ftnVpe6EeCQh/TYgdWs0KSA7jQCuttlhXLHiT5
ScAprbzgoITlYD9CpKhChF5f0vF+DxQlRSfD+B6QDT22yFVQWIZ+xYaAKPZeyk323kq0tWWyN7cu
vLpEB96ntw55DWbZBcdsd0PXcKcKoEql0HOO2mQLfKEY7AiKjm8Kr0xpREmP1mqQYYtNpau0mDc0
G47Bh+uP4O7JdD720BAqABmETBnLw/1SFG/NoYfn9/wLRMhHweZWFhToJUdhnZ3gTILMXWA1u5+R
z8/YuTjbqX7n18qx0jNCDw0S3Gy32oOAwoJvwD6ZiBURsWkHi5n0SpSyjWgOd6ayROwztEUAtCMg
KNEuC9GmPWMJDA8hfBE8RiCGwrY34wFmC3/ODSfROkdWptv5vyHMpooYvKQM0xBgFWzmBWqN6v27
kz2dbTD94rDabMZGSFFYtHob3PidyHIxTgb1TmLCY0r7F4ztKvIblXPqqRHW5896ceJ6cNiAg5so
U8uDE5ImHfKSNvglE1jB877QTD+V5/1PAvo6LsKOgiDdOwPYidxSB3bsEPwBnFlRcRH2Gt0fp3s7
5DiWTI660WtwuvoGVJD1O/aQd8PaxI1FAV3kvO6/mqz7VnKY4Cxm3Lo/7V5D3SrzUG8K2KtrBDLU
1rOkVlpxbHPSX67WMPWuOt4vDOXA/79g2Of6G+46tk/IiC0uq0qMmGDiQ0l649mJQxTB8/80RX0R
3D43uf3ISrZI/im/vuOxM5okXuY81EiLMlby9AYG6nciX0SppEjcBWJ6wJwuvpLdkIWy3pgHk/KP
AcS+G6hFiVoGd9LFMOiiNMUjKWsJYz1q7fR6yAYkW4LVSqPVI3mBqyIeapHVsaO6+1Atr79gXIE4
ACltVvutjiIunZeNYWXglwVsGjAzhZuARoLfa3CE9Nug3ioHonsLr5Dfvm4o7EqTnggZT75lWP8N
j4KpXBRaTa8dUdT/H9wijwxwubU4er4ewwrhywX0HvjTotC2fEkQ9sAQBMRwabgn/OrjmDDDxvC8
TlOgPETTPkeHTnl8CYHGwk0IMjUETMXRtcgur+85dZgNMG9gpHlXzdQDGQZtgvtZjH6nediH8fuN
AaIA526Z77ULXkLo0KsQsIbwS79KnOduoFID2Pk8p81jhpkS4A6l1V0iOjWYtJdas++BrkGmeigt
CxZ4mdfoRo+guhoacfIUeHQ3NRXijoynlh+lgAq/wULfKtXfBmIelSECBzXUxN61ZimLWvVWtZFt
6hLJn5cZuW4956vR3U/zBMvY7vjUBRfhW3rc3arMHOuSM14Y2sCZLpB4TORZ6rPm31b/ykaITxTo
59HQ4MulN0VAMl+VRa1aQyEpC4esk7XpmOtI21koN6xmi/c8dblwhCiHleSrKtuRr+MoC2Pv31Fb
s5mC/RBAYN898tcOfeJ6rq/wTGuDoUv1VtciQjxAsSLSwOhzQ3KrZNUpNHh96pEZRS9UTb247lGK
tIATD3Milpv88i1zQerJsoO7PlE/79OduL2s4unY51F7qvep4LGoAMixjyJcRwPznVYAaaP2nz/n
4U8POw9xRBu+ST6mc8DMbOPd6Wz+O6Z/ZM36KVrw2u1wGmYI9BK+iD/qqtz4Av/tL1iNO/4ew58h
hUt+ixxG5zasHGjYRCZOeJziFkBVHhImXepl/sJtkW9Zg57K75ZHIjveyJyHmb8xg4O+zVQavfOC
wcG4PQJiM6k+ozm8lMHX94AzyL9IEdmz4H8/mgJSdJMHaxDlERDcMdI8SH3NN58q/fO09v/MocOm
FZtpm76OKy+Gyjrstx3y0v0nfWSn9+S3g8c8l/g+Djev8j1qKYcpQ4g2mWjOuOI/HS1jXGvdm2eb
sSkMgo/UtzVgOM2DHnOcsj2NeSMfggGNDu3x1y5VZMOo4G/iyaf/s0XJYEpWdolKQmDwvrmMgurg
Q4iYB8cbiUNyQWk7eDihUvONpaIYVzay5JjbGLdWcGBVtG54XbA84lZbeeHe2NpV81OWd54FSrLP
bdzUQoAhJv+DMBFuSVy1vnKTKa4Jez0gKZFIXrc8S5/bEDI/+qvK4FEKb6UAlQBZ67udk8pgi1r4
sSDqzt5pWa8QqTyh4LunyhykyRzIBgn4Uf5IxZ/JLcCsfmAWu2r0TwsAS5dezbeqK3XE42vqhZzA
6E8avoQD5dojplhAIUYlYvNxsBmBFD/xPen2/nWmGRhi3G6PyabPp6ArlJuw3k+3LxAxrkBUCLMA
DwL8y/QUlkHxu7MlYWEnE+6z1G71RSo9AAOoqpPD+Oa0sbnJdndZnw1kbjAIUfBGdEr6nBD7PXkK
eunFs8nItCAgjWJrH8vb+rRtgX3rgbtmk/bGxon0+m1EHzUMFD8FwxAiuxRDPiIwimDcVOnUCorK
Pgy14w565ddkYcM5d8WglMuPrdIaEhI1nOk0oewCBtsQPh42DH/qYeO961ByhMS0U7J0ptbaN6T0
WWEJhIyW7FypXS479VXwNYIQXNTLPrEPt7FUrMtoMDEJxPSJx9tJhteE+SDVtzbXanbmjtAJEu99
2Ei1CgQGtrz201mSPCzdm8QNOUNJMo2X+W02yzGV5b1cq1fF3e+OvUTPCkqwWefev1O4T9iUYZkL
R9VxFnfW3GCPTmdI3IhzZwkInkn+mXwl/geemp36FHlUAFLUZeSuu+HlTHCMB3ZPULxdw4ZxfxZd
tWxf97cE5g5jz+e0XNMgUtYCuu5YotK3knbdd96udytCA8iG9xe6XztBpuPZzqVb7pv3qkz5uxO6
iGMuUbhC2gdjmH2ArR9P5XlPpXWaLVueH3BkS3tGRSAGXHR6ve8GSCdFgcKK501eKNhIC59lGwsB
1yWC8PXw+c4cB/3IF0SSlN189biT6o/7WFQewVWY+vVxdML33T1EpJCt6Njxq9Rm/LH7v4KzaD+L
jXQEFu1y2P/u00ips10WCod2pnnXfR1WSqfw52+88u/LhNFHTAcIKsTIt6nnUQyqvyJ9X+ASf6SV
uF1aozMk+on7XCuO6W6zLmqEvG9yZsBSN7Wt0175APA3ZrilvcVmSMh7DUJErPLnd5aTVyXWNObp
KJ3QtZhmJtu/dl/V1Ci7RPxGc8voFqI90/Y6SQSmsAJKroeAs3drkw7vqfGNS/+9S9ZIaLPfx5LA
/E4MHLM4zef5yeS5x73uOmSYI6caWigpcpCZsyvxykprVg/2iuDPbIlJU0CE4DhdLL2U5+K3BmyS
uwQsQXGzY+HvHPetN6PxmNQ+WadcCHFwYF4EVUhHYTz1zFM5dtKBjXI2z43hgfSJwjHEudTMH5a7
IHPDfE5Kt125n4DCqaLrCotfHr5T+CrLx3YK8dneY/x9re2KIVKMR7AwOY6wpkUhFBubeysihH1d
30ESph1IGSlTWRNW7a5+yDmHVt0njgOCjrFiCopdmWFUw7D2Fm+teN2Lg5Iq4hpfZdOxsez264aV
uLogW2KVYYCYR4J25uCJ7ARIThamh5to2gjlPaGhaxN4h5FaSW3QQsJZaDL2SaPLBGTnNzBTdzsa
Dbjfn74jkfM5T6GezyiQbZ+sZPBRthn8vIW6fP1cB+I5w2gn0wOdnRkSBy9OLfCFde3Vs8wUzwx8
ao7xP2uBV+5KkfQszrOA6VA3wvrwH37I7Iy7UNFOaMuwaVthCFMC2TyCYmpkDm3b2k+s6HzfiKCq
WyMWdtY1E2EKRkUcUaaDY5PB24ihaMFYQe3MqHZWpuAf+7PuhoPW8dWWHX4xPsM0WobdYUfEYvR+
MK9wOmwk87vp0Jn0eFfC+qtfZN8oPHphyNTxSfL44wHJIZRQ9OBTjzG2ncqgSjzeIrnChJ3nKk9u
XaGBwhylUcAr9vq4Mrf7rRbqR4Mo8VoF0+qGiCF5MiByU0RGx4V8zNS3DKMu/n9Gd64uHxWfVPDP
3rl0xJUqLwcU+qlFvdVghPvDxZtCZpidfzxbFstZdCyaUjJBNmB6/Az6eFmgIwEHeGZrgKXVoAF2
HV9k8puD6qY39KPRQY/W9ZXc1r7CTruDgJ4owKVVZhoWexsRT7eZVSK/BkJoSnceypLELfa1rQe0
A31EjABR5JDfXLaDZ8gedgJgh9a/5soZJaa5Qyn5zX04QNWCXifarlOpi+RBJHp1lL7PUjTnpa8O
4KzjsaCu+YdgBhjsrGLvY0go63LKDky5HKOn8Cd1U43DR0tFrp30pUJUWjhlPlVNla86HhsXNTMi
pwEeV6MStulhAcrlWk5wNGc2mQaIqnZowWIp3tnJ/ptLCjI73/MtWMI/ygwhn+Eyac3hgpPUXAKT
dW/svxoh6O+8t254GfaM5H2Ws4O4Igz9OeM5RsGLa4lthJwBcNHoejpaWJWXhOYseqtPOfH9X9ZA
eDVlpO3swiFFBLQsD73dz2H5flEU2Anf9CwncYd/1TjehmYTof6Nrlx0IzA0I/Oml7UYEsndwCB9
gQarXuE6fv8lBgfC3stUhBMway03Js3MNN9VW8q5zAgsF7bkXGVbaAq9JElXZnGyTgtqGuTDNHLl
3f7428nsiGprcA0nh6nUIoo3R0UYvD669r12uu/Flvz6dIgUMbznM1q4OV8zvyy1vI0ftTaMVuoP
+k1iNmn8elSZ5TVRA4oJgm4NUwdb0fQmf7XmvuAtB2jHp+7oOybj1/i7iFi8iJjqDSvqOPA9SVyn
FB4oyAX1v3v/FaC12pQi6sx1NXv6/zyzQPg+VtiWhOmC9gZBBlSdbxk6TyB45jAn4eIftYxXahLU
aufRL4mOPGu3yWVWbau65Z8i7P9swDZTrBdOSAvNodaNWVyHW/K45+0KR7neDgOcJqfrJ/1LAbQq
8pnn3Cm1Xz1HCYWTM7J9lqd7P8VBKbRGwNn/HgeEJwg5QUVxyCxx+9Pvg8wmrsPV8IaJwcy9kWpQ
7ig6UiuUxopynLElCIuvo0kXj2Ek7F08LSfoOfaKVpeybUeSrm0Ms12GGJGQBKNcVZ+m3dtGFScf
mfx3Oyiy1KuF8fowTXdlJCgDvnZ8IqTtWiQyac5+XTspjEAw+EoXMNWEHt3neMhS58duemZxUz8c
gWE+c6ZxFyt/xeG1uQ/s3KgDP1z0hAut8Lsd9DDUakFedK2XTxoH7qKKugP88HsPJvgh3a/TbvvZ
5zqTMIgJMewngcF3n5SKR7m2/22dBa2MITdLd9E6Nd11x1TywX/IjJAd3HG5lDMOSLcOXHfzOMZ1
ejbc7udQl7cOiBDj7BpuXpuMKvHhQr4v9oEp0NbWDMesNveCuKTSxYCXCHpIgdjunoh6SYFADOO4
Alj2pskP0qnzrpmS6N9dkqx4QE8E631C7vyHtR1lSEaXT0MRTRqfOFC6zwL17rQgaX5dPH4vEnVa
pTDo7WT6mvG7qirzvuMkwh1aawY5fsnf6ygQk1AoqRZwadi7SyXPbGNeAmBjCTCWDXg72fO7PVgG
Af0289PX4Iuwmpa7LmIN9ICrXBUXwaHg+srBYDYllEXQQ49KQqZgEEwfysxHtMaPF3ijSkMWOcpc
Y6vvAUOBs2kGOgnGXP9O5dT1M230IK84157eHw6QB4Bz1fIPqAkKyzP6A+rbxorAKz4Qbs2koBOG
aHbdwL3HJAmLMiAXYdV94IgLL90qEZXlNLqvqzV2PElKm0oFNSY9Cci9hqpoBTGsmgpyWja8N6tn
DFo+CqwAeZFzXMx5weh/RnnVM+4Gy86Rbbxr1i9URCm8BSXMCpRIUWExR/kcUZC4kS9e9TQyzsgG
R+cpDxII94MYbkXJ4UiVXgNVUAv92yUMc2Xa4vMgezwVciWJj2TP/bG1EfGdMqI4wZgJGO683IJV
0mT/F79ZPKcrumIkWCrdn8mHBThr00qPCwLGrnatr5XMFCNxpijcKCMkQ8awtQryP1fbu/W/ICM5
eCregUGesYgIEO8atKVMTavgkVDMdK/UngMakvxhBX6B4qZDIaEE/4rMMYdMLbVSlidmdLMcWrT1
VeBYGUP+RtVdl4lRTlbC5ZZww4euqv6jUgzz82VxfG9FlwtEC9oh5YCt75IKaeOGf0R5an3PZNS0
iye/c78wtRjK9d/J/YCI6WSqnOIPQXhVRpdu/F1gv80l8o/jTJTAImRCAPuzPkxpOqmNGTj4IMOr
jdtnAJynveBhKC9MVQfF45OuTtkq19U4rDj+PFII+nl958z5WqpgD6/fCQLuZ1lJMhWd9nn5CFZJ
uNwPk/iZKbNQHgd1YieJkfQa9K2x1TY2fyWatKchkRkePm3vP9B+4rOv1+b5GdQlGv6wniP3Fx/K
iqRjWvxjsBEeDXQnn96tme/VndBTYoz5NSWCxubLPmbeRi7P7OzbtdP89fb7jsvFjyn4+EfBRl7W
s4Xh3QNPukJ1gvN8whQ8cfxmu8Boztj+IPERFOt6wjNwyiku1nmbLf+BVIG/hXctarn8QeFiZMTF
UzXqGT/hAGsLUQpNIKmpm8MXm2jzYdGGJW1ESA6JNblIhmG4SfehgI2hru9B4VCG+70SjyK9ZOds
QmtMcMdl13mY5WZW0iW//z6gl2iMpqG7Y1rzfbSSGXovtG9XlpNjqWErHLu44x3oakhYPR3R513D
P4NJBkzM21HnFKbOUvBTgJoUk+mheIBFmxyL0Un2gqx+O+o/9af0vBeY1mRiiJssagta7zlYk0v0
gUWFeWwixR3jkHjnWNcoY+RsFlHg8vRAYrHTHwA1T+dvzscWJ5yDG8UTOZxZgtWJnwY2X2mgNAhO
poH7SWRPOCW5+OPxjp0+KDsRKD5Ly36AaJv/wGAWmotljbgyqs2fsvenwKYq3SCp1igpSX+cyLyN
8gwYTa08kIzHNMd89Y1SNewqz0lArAK/mtzwDh6dQ/0FlIgjVu1QVUjkXtB2ZRtzZ5W8XWucFMEJ
eOBYIyXuyq5sADcbuUmC/68VRh8PAlEgHEjsL58Tdk9tnB11mqEUTdSA7n0ZQjz2Wtt3JoVTAgu+
NQVeNNo9dmD4opULcwnD9aYLm2jMcQ2p7fMr3jFu/h8oxRRt5unTjn8COb/7ew1Id0ah5/mEJe1s
RCEXx6k/rhotz4gGKrv/iBO07tWheejAeRQwRpb4ysf4gVDMuvZIymiEGOX4KshQSgaE7AjhLV/j
HQzi+DriG67/GLdmn1zTHZiJ5qCBvupzrXUTMf1mdKLMJr33i5Kr3Od/NDGmmEb5d0Su6NOPybWO
ZZXql206FoEsfvXz+A8wQOETfI9LIw08xJSRAdWz2FhtF9GV5YAwkbyYZHX1KFzXbaQQ0ePWm3LM
2s5O0wq3o55kLssOma/WUhSMN0H6RMFn29FOvcsQX6sLE7XE84ej2d1AMVmczAtmuILRuYBrjU9o
dYJL6pCo4nXPsxOOLMR1Nc/AU4FzriHTAKHnVkoE3phmjF2qKJ+oioF/jRdDpReH2VLAa3Fm65sv
X2ueSDRhWFN0qzUBk60K0i0SqZVvSfY89bEr2DWC4W01EMHXuufWbbfQvW9aFy3zPgf5NBMUlam7
6sIiiEWRQTFhaMChIST5GC9z222cRXDSu61qnoY2MG4Xbyt/WrjOI43MAiZk/1jYUBSntEjLuMGm
6++TijAAv8ONuoU53BUyZQa32ahj+kXUB/RJ+UkpDNxmL7f1JGFllNxiht6c3/Q+wvFX8x0gqBwJ
j8X1ThHJTxFY0aPgPr6v1CEwfSbgqonQX6xpNxP3153FP/TvowPg/LpcfR3GYmcEDWZmSKyoAgfR
0VsRwv03RtP8jE05gnI3nHJ3+3T8yfd4GHlgGf5eAt691GpNK9byG96mVTR/cIyaLD4lgC8tKlti
9reS9hxupJboX5kw6R25OVaMi9gF8z3SqmRk3vmwLC2YUcV+NLhKHM8QjUFx4uzDZidKXPn/PaeJ
V+FiMPA890sYw5gCh80k4FBoIS6qs9bFxyZE5jt6TI6TjlIHKKBpIa/YRBcIA31ftVCq5BeVrtxM
HoGHKqLFmFsSUU1u3fZCTA0ip5iWO0pLC3cs/7Rnce+3P61ssMxDYuRRH7zY1FPW/6UShITPHST1
KpplxBdNZjD5DbCuw+riJ8vO+gWjHVkFOp4nAyh3Ly0Lv6lW1cgGk8as++xos+427Uh5QEZB7fuh
2+hDzhru8oClO90zGBIOvMwsd5fLpvQsh+yXZuhPxZAG+YMvPwtY/8JAPtv3ZgRwNonY+3g5OF9L
yrKGzTjN7HFOc9ZrVTvFiMQHuq/Kcjg/moy8PeUhP3yoyJEPu2aW9JZpp0/bnZ1/po89uQkN1fsI
u8OePJtxn4kv/vLkvB1k9ufdvhFYusbvEgwRxVB1Cy1pgUP00V9A2wKCD2sSQze7g7932bkmA7vX
O61c3F3VVGsvb+fv1hDUzM2GNH0Km0EDecblglOt9PPOybVYRcueF9S/Ih5rY404dPL5Rkt8L4kV
BT02T/Ek5XuUm9qPy3Q7M+3sBc8YiY1cbi8DLCo6D6ymyeLlST7Dcv6+Xr2R1s0CXpUNvnkrAYlZ
6XTs09txks6GajAsg4rkUX6k/xdtSBCdALxadlf4npukdy+JR5X0MvZF5yonEMFqhBH5HsjRUGEG
lUno+zfNCE8tlQrYlZ8hwbWqjEXnvQFZnKx9WiigQT1sQ0DO22kSXWD9gDDTg8GuvCmvNcuao8GT
IBcOGoyAEnBza3KzEobIGePaY5r3wN/P8cJ6ZVn2CAhusxIYhbLUPdXdhgMkJVybc05QU2ZhCTGG
/JQSWzCrYSvB2KbHFDlp5OPhNUj+O4IvadSnvQw+1yUxpgfw2xwx6kbW28jGheYNSsnE3rCxidfC
xFp633ndbTuNUEdvuepw9f4iQNanjr5T4VECfuWQatMul2ecHkZNbNwukQCGbiWlsBQLxvhJzq1X
CSKJqvTttuWDb2gvszttm+PDyaalFAeBfDPZMvcrVwujqY7LT9+V7YUtOliq/1BirBLWLoRq6bhN
k2YQpdjFiyDzpz6IjHc+rkbbN7sgDGINULghIX6qdMafvcIFUjf7JGPmyf6p5jBRkrTASCkVERpI
fUvU1PijPeMDtnMthc95g9NQX43nHTZUwTmc7PWRHSDnsiV/twyJh9M27NUiBYdpcGlfmFGIQk0x
vo6b0rFGeimXIF4ysD1cdf/24Xif9CecMLt8l7bF/5a15NNec2gbtF3oOSbr+gyI/RwxpzNmkLs+
RsV9qMSRMfkdsYNoAvgRJxYY2T8PKkbkXr3ZO7skyiPo2495lEU1JQD6kbI6+0PtAfbYLx6Ug7wJ
UAhaTwkuZKrl4xOoWLKbrBGkR/3e+cS5YQsuuUcIbuFNmq/SI3JrxQI+eycC4nUCy1QnES72+OpX
YL3wFDlbpt+Hf+2uoR7KAF5GG74QK3x714V51a7uGbgGE7uprRrmIiSRrEWIbDW5JSSN6Bvs8LMI
S/Pqr0XdueXvHxaYEuvwHp/Ghk1IhvJU8rIGgrhhdNeIj9zuSkQWdNvyx9EpbbxOdjyUFRRpBO13
DVGcgXOVxCK33nIcT7XIcvuOLtadyTdpcK+RhSFKwKEswfxUHvUaB5ANe9bYCw6SWzmKA3AXKY6A
IcCB3YQS9rX/17H9Nil+LTd5Sei0oT9J5NFnt3YRpGnoasSRtw15d4HRvhAU/uHHReggole9kgU1
1v9PVZVM8zZYzKtdyfk4xCbgwRPlfRm4oaMnzQRtuCdPFB8FApWOn/il/XMRaug2bnuOlJtf7/0e
4yExOlEBBUZCehB+H8V5UJhrqDoEfKVIPKp/SoqIzKAcKPHAOwXYsToWHL0ilcmL0AGCZn7hdIaL
xtzdprMVgDyen6xiTCHuyL6Yjz5VtZu0ZVWbWlP84IzihXKrsiMu1GtoKwtD/7D2KXwjrF+o5tWA
D+VNusAqPAQWduHtwSFqDvJpzjs3tF24ZZBnd7JTTvMxTpnGs3CWvdoTza2vg7URSKDkDwpILct0
76zukT7GgCsQt6mZs0etH6zmioVkgP1Iu0Dcz2fxQBeQYMW9kB7eYWJYUXvfo3+Lpu8+oSMig0FO
akzT2bSv+gxR4Qqedm/du2kElq5M+YAagG1LEtOZGFqvFGUKaOV88XAFgRDA2H4XObLSDLxh7OkT
sjEKhfoC2Oa4Zs+enIbZr9TgU0RIFJG9yvzz/7xkcLoUsJHbfYE9OZkoJ5A97ayG3h1yd7Zz7RRL
s5qS3OAOY8mhNVNJBoXzF1Sn9aiNBfCtZWF0WyqudVdb8FUDIQCGqsMA7uhFfTCPwXpqbUNlb8v+
OrD2x5/Col3SKKlRjkJ7HsnngUNEIUlHdApCSlu9weytpscHOLV9QOwXsDRlxEZn2dxuE8rAi9m9
4b4IA5mq/xUXDa+VPkrovCsu6Ees7t9SBU/7Zk8A9rHzn4p770ZyfKLiblh9dSBxdakg0n80O1QN
CWSSTEVfGKTnC8OCPA2JyV+BvDyCf8Z8fOHKJ7R/Jd2z3A6NiSXWiOqN7HACwVDmKArW/9bPW/7r
PXStnzU7ffdLNvaCMWS8RbY3mFDfNYgh76KX0QbpI+2BVSFQtXZEl4Obipzh3XJ231lXOXPi9deH
YfexXeH3hGKH5X84t4YffGysh7EsBTKxMDKifrv/TaCa5d7nvOZxVEZvNwPxWWFYgZNWuHeWR1T2
gvz1+uzgnbpPIRnG0fwvnkrcoWa8gjgo2Av2CbOcWXGtAjTqmVoPHLJd1PIGDns5N0dLZQJT9IT+
4Kq1w8Ge4HvOK5koBseEGsdfExaeNJyMC+B1KfQ4LcRS0xhlpw8+CStZuiKXPGM0zVm/bb34/VUB
qz2YLHjCC319M+BOffAQm2sgMf+Lp+m0Rv1/ZcoALahPXENK8PPnbDDM1DkFR851K7Noh416kgTx
unkxWBPE2GhuMPLJv1HFkNYUEKQkuKcfPjqw09EgcBlZNPqSLXRCxNMHobFMoVx/VDNkpCOW3/zj
+Pl76JM7DdHS1lp4Ss82tYfkyI84mPrWpmx3HYJoEAlXcSw180/lCJJhArP5Hv+sB1AlO0Q/8HSL
bFBnD3iyirLADL/K3bbjVY568WieuJnUSGNnONsBPFPuh22nfxl5JdVjcr1m6EDouj/x8mAvEDy9
1YtOaPg8Cwiwg057sYt1eDUrYn8stZ5GN8lXP4t7EwJWGWg9MKJpwI7rOmKhF0bpuz4v8e28lpad
8wxhGt4q2CnDwvN+5sKo666ii9zT0ii5PvnY5wUSaKrOhcU0zmjBWAkIPTp/ySDgd3CKnizeIaBD
b34E+KXK3QSG4KQnc8ljWpoJOyzdoVMS7GK0bnwM9xa8lS7NnxPd4TqRqfxgCWCn8YyosyD9sIkY
X0nqNjA47QiLs94TQEUF1u6u/xhZL4AY20JcV2xReAUDPhWJKDA1IZ6VwdeI3kxrUiWUU8a+IMBR
7ilNWbeid1HWSnIEV701geyuxYnyf0AhpllgBKbdOkTA/068MbEAvlQHUk7Nkrrl3LZUwTVQjFpl
6o6ypJsflxaoRyDcEWOsgErpreYnmepRf3Duy3G7rKQobGiSPpW+uX8r18FqpJCH6wN92LWHpxNe
Xvf4PGpdut2xb6P6OjDPF/HPPU92+8LA8WR9gtBWnxOSROG7Siz/c0uUQB+PQcG0Y8PpgC+vfVjx
d/mg3SSaLMj13ma1M0/srap5meLbAxEpGXFx8kfVbcWZo81NhTs4YacrQdmJJE7PcsaPznruuX7g
U7vOWtYWSPkdzzO15jmpy/xUEuP7fDF0H8WvpPkBBusZCTfuMPmwidZmTl68PHjs1v0QxvlAcBmw
bRV15L7b249Fnk4jBrEH7ltTHD+aPZAA6jgbt43Dk87CPJMwPLgYdm9eqpCtuknLjmt7lRi5Axls
+3XWYE5vlImvRzgNQosIGdqB/prlTNq0Ga/Ovu1QJX2exuZoDiUMAWxqoj9MOXG7Rzl4Ie0CrqBX
KsPTqimMFMA8U8seAjMTEQkUynFhqXNfTpWiOjMVpwC2YQYnKlSZhElRtYFwm6A9AwNu24HKw34C
4llW4me4BzvUJuOj4bP7xmjvv2UmMSiQhVR75aMxGMyZFSTbfAG3cTFkY6/SkMdeO4cp73rPLBUd
J4C8YZewHc56T8VgmbKS2BmnK8REI8FXdNNp8NUKuGnQ8lWldvX3CNJBrrfs7BaHuwVhs9MzGgag
2+w5j7sdblN69blH3mEDTjClb0xUK9ASemqNIrEiDS4/v3lYQl51ooo0GYaf3hVn7TqtOqlV4tQ8
5GGLAgXpHuvwToN9haq332l/YDObt9DJoD/c6pu/Urg97aft5gfAGCSkxoX/Rn45S2zZ1u7KDVB6
Um52Qv8W7eY/6MS8Y1z7FYrR4VbexNi1MLicrO9h9MKJHoSqyERSbrShQhx+C63DtJGHnOI3cInl
nRoMXdAiL6NbhQ6xTtYp1VBYzi88GgPNXIQNYVqwaGOYzUZfTiZ2IVFPGAq560oLJR5fPuY2IhDg
Jsi1cjrGw8LUf9OPMdh+FU5QdUw+udFVj6QCT8ca59oe0YB1KmNL3tqYfjQrUYTmIycWJVEGDA6C
Lv856ehUSvVjfRlZV01ES1rDpVr0vN1UIa028nBXbrKyapm66of7UkLj4JKtLEohpmv8fR7rBgUE
DxDOOkGR+SW0oV6LgUnwdeVlM/QlNpM8LPKB+PMCty7DLWw8A8xk3mSUU3DwOSUlhZLb3vDY03HL
4a4HrIyXQZ5zjh2RqGV8WnnG1RyM0yVFPg9v9W4q+RqmGfzcaKGkQIei8Xiw/zN7gZS+uilLa87R
xAlZvhvFjoWrqNLS4ECVtvJlKj4o4+XmlSGsXtkzzCyqh6oC/CdvEuPLxHfWhuYcOyHtqkHfqCfR
mAfTDUyh6bSt+fGYbGrucOw8BFR65+KSwYBNaokcT4XlrxxHLs+WZ++r1F3jlVqDTb24xuzIzd+D
i4y7zwaa8VWR0Hp2Ux2JPLMpwdXZAvZMdTFetMyJM5MXaiysyS6CaIXdELMru8ajGlEFJSvFi3aF
vcW4Bui5X/5p2PYcxX0Vhs1PpUvvLPuzyDnxpGb3yOEKXxnAJokThizrF4PqktL93aiC8JvN7xYJ
qm7NXqcD6XIF/r54xg6YvG0IdeHVGGUU1QyWhDw+RaXKOj8ISefvpitteJpTASuDVCn+ePvvxkyW
x6nimdxSgQn/hl/78DKd3fxiSiS+BzK9ycqXnVKu333QucPkwge0157GTWFfMsMU7m8vnaZGOdiV
czrp3az+lXeOQAy2uiXk8bd4UTjR3RN0poPhc6rx9JPSZduagvyyNZC3/BZy0kKizpXaEnb5BLqM
FRlLqRtHReHJ5hsTguclJ4VDU4itF9muN7DGlC8lNrO8fAv0xCyYZo3af8w53PM48/BEVCOXoEp/
X8o+YMqxfP2plt9KLbEIJbawuYNMimbPtqEE1khqk7PAZOMyVkS9k/S4krjgfLpq4qtHo8lSPRuR
n0GfbIumRH+mjIhJHURrGWqDkIfvF74+/nbDiKlNGJ97RdloJhrvM7kw3Qe8PEERqKU+Ea+G4DHS
tOoXZPMvQEis9ytpbAB6vnKFBBWxnVjMu2wgIPcmmugR146MIk1udIuJ9QWeq7QSrlI5gypsGcNQ
ZujG3WzhUABvaFczc52pplwYiVooQX/mOGPAtf6damlZ0/BorPSvEZ/AD9kSe4l1s112v+btWR8L
HJAzQlkh6SyA3sA0CYHs8qptwnN9DaH2dmn7ef1BFns5/wUPs0C5HqgMmEk3Hg0svTLmf0QTG0Tt
NfMPYA0BoS2pmAmpujOirBqwY0uWVHgyAeEDN9SsPbml7iCaVHGEq4bkx9gc+G95FDYM0jWEc3az
OIeES7VH6wOqqh2AnEd1L8tTP4tZAJL5qLUNxrb7ZkfOPBUaF2vNXsaOXGV0TxUSmwZd2NMy9Zj4
ql3sLSaLk5UgRBDZsdP+AywQpfFsnmZv50RLNeU3n8J+yU5+6WP/MsQwKa93yGXYOMnh6B9Ql/qI
KUoDBORgdQTLUB+diwn9wD5LwQuDh+rbRX0aDGroUYxqerK1uzK2gaUgvFouO8ecunk8TQ1O6KVs
MIjh6wTOjHNsqz6RE+YqRLH/gD9wqoOwbqkTQccJGx/B4GLrnzQ0IjoFYLRNvgpL6XzLH2GdZxik
xFyaSMXzYSBRY+5mXfpkRae/L+4J+OLfn1DJa9WbN8KJYu+mMCC4W7eQXV/OArOELnn+Si1ILYUF
FNu4QknLAC2BAKrPXV/pp6E8z/cGjJO4iRax1sA0FxfSzYm23huGYGMJl9LIBPqc/44Hh5PGWtGN
LGBzbugxkMzN3rn/v/7Vj7LIVniwd6VMa2YkkC1pqYU+h80iJ1CeCY6NMkxz6FsU+1Mhdzukddhu
GwnQzsVs2Ls1xiLFgTV0lx4e/+tzb0Wdh8Zok12DmMGfXMKn7pPLLB3Z6/UmMFA/UoPp6H2Hr/Hx
jigyqhdyzhYaKhlwJb79NlI1LlCwehwBDvgYemKjRxvop3yYKcPOPKiZgb24SsaainJfvVmCcXgf
jUaM2Fpb1vMBB0UzZd8JcOABj6AKUUYBHCyhBolvUB4kbrQQ7OFA1JshLBgGWxyI16n5LYUcrd5h
q6+Jx0ujn0fkT5lLbM9dGz0NmPGw3YoZ8z2bEmoBMJuyMrMJ4mp7Gna7d7tFTXOqk9Ezb3iUlRlT
EcrmekPEjP2StxTkDO7UHZja4/69W42yLhSv2UhC3eR7o9dkJXrKr9I6DmGmA1RHq69nZb4FsjXP
QFSsPHMLnvdRZ6tpT6EwOmcvb+eaydYmOJRhAyCKb8POpmQT8JLIG9AxgcML60Ppe0leJSxy6WeF
5BAm0SFKBAbPPhM4dJjYAEISNCwgCVNEw9ry11mqVybPFncjw0e/+yaU0yeWhtRC5lFyY4wiqQVi
CIXK1I3zh7vHogu6D8+ycxZlLQLUIvYacdKMVegyLpNLxj+xF+KSX9RIDi8J3aFH8PS+xmss3BLn
V0mJjI0xZwfBMDjn9PgxsMVJuTulWmgq9kcUY2jh7D9A7ckJhQpmUAqiBFhBlKOo0YWbOVUAEVIg
x8K8URwDjIEeNfJaMMCsYcCvS1wQum+4sYte7U7pWojORNXhtF9O+IhSj+8hpZtgiyjuhy+CE3hX
5sXCJx+PiKGWNM/zOt0Qtergyw5lzas/KkphjnlATxepwz/GZ23fHquqjUWdLfEg24b67bklEErL
jJXVxsLBzp604UbIGX4K3JeUYzz7UtY1al0p0z1/7DPGmZIe9roRjjWji0cImbEJbTQhGvXR+HSu
Eo6nTuHsF1D7PllNFUjaFUat3NKYUm2A3rAbX2or93SJwyg7g6I7R52jEL+rFv9U3ENspl6YcRm7
6iR/bc3CVkkMyB4/RzlOwod2UESwPPPrI21zcV/RvThskxuQBUfcEpu6mr84z5QLkpN4XugILTsb
If8HUV+jffevcPh/ixa7nPce5l56bZa3ekfEOptTRptXdMrgQb4cK6mKaFv+rdbu3DEHz1o7KSPa
MptCCnnfYQwUWEOiO17v8fhAE2FuaoWadYnCtZonC54I8+tcJmR0l1R3VXer8Eww6EB47RQRgbjy
4e8g8bkZES92ElDduUUfZcBFMMW8Uq9atIdfyTxMwdNNDTdjTQxk6b1gZt4BEXKJikCtzPemKZoj
KzcTuaq7dOViHQUzMwKqxQj6u2m+WumdfPK3oDvZGbdXa+S6vwFLa0ThP4j+BxDT16Za2JQXF83Y
kCDUf62OT9iXp3fEsMTx8JY7tbQeT3HckV+XOzKp6kabetPGiLsFVgfWmJro8p5fiiSq0mWOVtC3
DcwsSt+Yi1ZrVVfwVnyJuuhK/Usqk4UWH1zcnUQTIfVBqpAiWf31yuTiXSHUxMr++saVZ3hRNL+A
7Q0Qph6nqtUPxXpn9vIxwss4rWJsijByuwW7zcA8cEcYBrTsBUwduv6umne8LupEcpbY0OIua0mm
DeNE+X/bWvxfvsb2IfqrDgRn1wMmxWya+5CJB6i9phZZt+VG++vrzY/W5HaR3j9wdHxdAqZ66VWa
IZvSKDtQID/LveNcOx02daEcbIauWEUFjyI+uW2Ez2V7zUlgdGxpbspCgAy1fq4AvuvCTmSyRaa9
l8A8k/uiIIK9IqdaxIDjkMpCHu/ywgLHYvW/0OY/mgHQ5jI2ZsdSKUFDLK0nlgZKRuF+26AN3OGU
52UEuJhX4IvhjB4Uy2+gQeoQaUR827vhFDIAy/W5cWM/u62hMF8N0T0dmrEnGF5rYjXRrpdD4b8q
EqNLtYYcLwINutr/gNyPM8mFbDp8yuv5UHwyVJD9kFC/m3tgKU+brGQhmYUJo6WyAchOhZ5hdsuc
xh8I6AsxGzKLyJsM+dhVIBRKFTQsJKqBh0+LsJGr27hLeiGD84jog09m8doI6NbI/n1XYRuPxosz
N8cVojw2O+5vhY2MqzmqI7vxUPaZWXY1GDPWsUqpmOjKPh61vJvBKRNSvfjkycPGDh1k2lpNJjy7
wNsq7aHTVFQReccMMtPvpG8Ns2saBs2Svtxvc8jSjZZIjIVMpoUT0rqCw1u/xM6xuatDI9U3aBWW
3YaLUd+rjMIL32VBbfmexXBjCmF4izv6eqWdiWAEsBV7wQrDIxOYWu0eXNE5qMlAWKX1q+wF1E1H
0wD1BiSGQm/FFKRWYiuqhbQOF0iuQC5cVOYmuVnebvVrlyFpZe3Exxvu3V0I4dg22TydzS6XTUZh
XZESz9GP08GxPiUM/nMFpmPA1crfZbijTkl30DwPALKSp2pxx5wX1LJjXm7yEtIzf/0cb4msfZeB
4kNLzRBrAV+9zaAQn5pURrda8jHd74McUSi2RxaayWZivNk69PJY93dc+dp9P3yi11cXGt8DHCFx
I38TWk5aoYgZtdIaXSD5xJZSFMuR2GOrdsyCWOkruWsiKSNqoFFuiqPndBo11bA+6BUS/1m6mnAG
5KfcCOSFNJjYgI6vce8Dc3bw21wqqZVyEKjOZ9M+eOlilNE2tTjjwVmqkmIC89piKLLLcqISCAQt
vG+P6chs5MOGd7CHr96MyRlzUqBKEEjDBHjOyISB9k8Z0ChzCFwBesgZP+MFAQSPLekzsMvfKTCS
D2GWlRPqnllD4hzosFDzBs1hkKLPRYxyHcvyU5MD1aqukDPCAoVNjGdjayp2mbz7j61BLDgghbKE
hIpXx/KO2s17I6vFzRihF0cXDD5ohYz2ybEIH2uSMGjverEvbqwVXklczZAkCllHqSTqGw0GisTA
wKhZIXHqdBMqc9DechsdX0O3mlweEMaOWtlTpDSdqTSd/wiegapQuU7I816xvCSaaAqco4fi0ZkL
g5AqW5uhkihxhbZJZ5JHv2EsO/aj1dcvM9rp2J2W6WmYg2xAyfPbMQh8KD2/UkTsVTb+Xx/PMPmn
Sy2OizsB9I0UX5+YvfZtd2kw9e+u23kao71Vt+fGDusUhZmZwDNPNWavXZN2bRq6+J3/H4PjH15w
dUf4+xN5Vtj0pRg6p3dsnO1xYXYFbSs2qUXcDF2hQij3Wdfl1dwl+lwcWBnIVYdls6iKd/OTFyxI
7ljkVcemL1zREuEGvmdYPTbVjbo2FvxC5QlAY7kBbpQbRrVBNQxRM11HdDFPP3sW7NQv2Ca2879q
Yq09GTiSJdaYjxAz+evIvoeEfqQXc7slp0/ljdeJ90DjDCV/7Yw2nsLVNOEGyBqRGGuUlJ68tj02
h0ylf8FIgVH3/TFTctXDaiWVupxEkBW/GlE5Hg3wdgSqLHMStX9y9otBTJCrcSVYCJ6kaqQByV2C
+ro4OWbsal6VnKGuDHYje9zgvTwMlzbwF+9dtYHOz2znKsMjjON0VMZQbT8lYu8VVxTWKhzJDaWN
+9ICs92ynjpsuzuHslHyJ1dEh3LqtvngBGoqCOt+MXBPIEqwqRDM2EhAZ6oPxF2l1mSq5sob/e8G
1UqJ2mPuIzOOX8JfrVVK7BF+LLqwIS/2hkLjyXkHIV9flcSrYahLHXipVd9zWnjF2Rp4oBzM1lwJ
2jvpiAvs7oWA7Y1N3HeCQzoIhkdYIhdUPn9uq9JAquAp1vt0O6K90nr1Jf29PgPJRYMZ6oHf3AH2
hI0i9RJixE2a/jaTx2+yaS0DbeTQ0KrjvZ91EoJERhtdNZckMRZK24j/n8DlQZbBOhuriafbNQcQ
iJcUesPD00aKIzteRWA6FNTYFHFqpgOJlxPSgcbOW9oA3hPRsBFHiIO19tgXUnoMfY4QpFOGSbIU
L7tRxtlYvu4XE+CtgJyzHnzHxH9jlcA63fxftGSwCbGmy0RikpcgDvayIewRDPtNvn89mqCitJRr
WfvmG5RHS6pA9CI0q0riGbhG9yp4kQATIilWasYyMmuv/YVGn4m0ZzdPecfVoAf7sS3djzNIPeI/
lJrJuozWr1tAlYROO83eDw7M2UWczVdKErtqytTpEsXtIvpL+xPb2nF/QEBWjltcbjewe+XET+41
l8b16AVn3PqlM03hYkjS1RX8yKh8FZhR03/9GTknovZjvaieBcL6rCFetNdAcMn49S8vSsluXJYI
JFgaD6xupjYDw1etcG7/bDjOtgHCmhKxtqkn9cNCQfqDDIKfAdG0fAXXFf2gKHbdPoGpZRoJ1cFj
va92tUUgrN0h4QYdn4dWTgB8xLfnxS1Y0lqO3edzuwK9IHWG1sHhvBV1GktnAL1n5GEdpDOJMtOX
jpQN7ljGjbFrRQFrTDjBQZWtr0Ssp77vBWMzntLR2O6od+dUPAdJ38oFmlJ6CWMIL7Fd7WPjVRX7
hmSBJkK82orxs+BxtW5ruRAFj+jrzUiEXFLjmmkCMUaKHDnkLVpxJqaTlaDo2A7KNqhPQXB3+S+5
5rHnb28Ks9tsvEbj3kV9mH+8aKETKXDN+OxrweX7iues53Jp06cL4KZiZN3Ph0BXR/Eg3iz//P2M
cgM9W+/zSkIjAModksUcsHCyuH2v1aDvFYAsJ4vtl9/1vj2EdTTV5BOCLp3/H01+X1OSkJeWm8yz
VW+36qulUkW1zDZUrqmxCgDrJtmlwqjKSG0oVHQ11E6CM8ai+wsskGldOa8JdfCRt2nFo8TKI+S8
EwAJWDgC5Eb6Cdu9j0OA5++AJ5YQ6qQs5s9M+fUvenXq5k6B/NAN8hRHjcO4mDQkZvCT79AYdmPd
MbJT3sbEu9uYx3rjfPjJ6l2CxnU0oO/5EHYR4qJs/funjgag9zeDg8WfQReNqvkKgn+azSpVfVux
nG7BHR+GvNt/yoxqR4TbMLY62iVG/0RoApkbH70uEMtHeH5NeIMXS92I+u+LFwWemmVHyYnQN50C
xE2dHbhNOT85yQtrb+Sqa7ziGEuzrXyztgZOiE3cI5n85jrtfZyv9f8t3oQNX2UDcu2atO7+zmDP
75RxPuOj2L1vueKl7AqH9w6abYyWs8wVABFZNUw5KwrkClTP+UFzrDRzX68Oqd9W8IQBG6FxqXIv
1fDsNYqvxTtGpC4feVSGY9AHuGqAXbV516Ep8AoQ/xkjFzpGO8NUv5KXG4vkogFsby53rqLlcywj
Q+z4K7/QoHFga8GWkqoTWJCbDNCR/xWPyYsj7FBEl80uYuXjK3M3pnfPfMgaBgx+ZWJDw+KKOl8g
nEuffNPcIYxIilmcZtt7bPMwhYushuyeRwY1V8PVLE80NXfcB10nkSaBSdJIPlmrwbhqYbsNq9ri
uA4T7mvM6pgqbGhqnT0cq7/CvSiCE6JkAcr8wJUmsYG2hKn/xPAesCcgHXd4yiQG9cguybev9cyW
2DdeWSvvQJdTe+Bq/BZbhzldrvoG4mW2nxCCvVQPU/P8t8tE7XWw9C4VfzLwLkHJ6myE4INxOnNf
nY9SQNCo8twWU5OEtQZUSqxQ4dAeEvso2dijcGuynFQSiUQ6fHo2s/N7730kdlbJuvxepodhB+Wj
tBznIsUuj0NjlJemYDIUt5FbujEmEaFtQZq3JjVB1eUecHd6ZIgHaW8sNSL+eTc+hjBo735WG6CO
mmQJ1JqTtHohAUm8izV2A8iCl/gv5FSqqKoTpMiq6sAc+4N0UkpFdRBP1ONRMCPi6WHOoWha68aj
Fgd7Enif7RKwMBCZ+wWnbTcu1/2hTd73O2US8TotiM5b7GkRYXKzXudVMRAEhxLAYKeRnXMviMKp
EkFPBXxk3NhrfZavigd5JN2MPA3td+QvpL2ATtscEukBzD93eVvqf3tHM6QKKxceF0Pf+uBol4BU
hAIOpoc5F/PQu8hur0J2FCd2xTDS01oZreK4lSE+CfiOxv12WxhvhBjsJ9SDr3cXCdOwfcgkv8fX
YVvM8R4k2NuMb+xXh55j0gmy2Kn2PUfcZlAzuBapE8+db5B44CctRZrBJYS0VIU99RA9f66tOw/h
/PbUTsjjMFk4ZlveRgsE10NyH80M5eE1u+JsEsbCRk06ywT0wgDLH7kdIkpL8V5tsuFtX30JibaP
9WOk8ys+oJyWEa+BQOUB0pJppsS3s8NreJLxYZKVxdXdnkjyUI5+mTbEJ9TdqMKLj15ET+khXLLC
igTGTrfPZDOsiXmSKeDvqoErjxUn1mCO7uHu0AjGRzesMTFrLwyJHRqrWQH1CG7CfGG8cvPRyZwm
V01m42GJaXr9iCap1M33DsUb1hhcTYTXonx43/Z9Vlgw6C/1w/B+7NpHtEq0EGLwp3RENBQBIvQv
XScSsq5Sb0CVWFR+G845K2zu4c411uSTglD+8qLKxyTxXDCXWAqwil4q4D/Av2UkW1lkyo+5xYNa
A3rk9xfQa4IqIEv1PHlKyuD3MjK9nwLafH/uu56qr4lGvBNaku836zQsH0SNu45tZ2faEKSQxNEJ
GfPuP8Fe/jeEaBlgBYGoKISrjD8nf8jNQzHwMw2oTeuKPLvkkKFE06V5bGSzm8MbGYkdVHnEGoLx
1xfu+IRIjx6pcK8ohwCB5nieda9Dc5O5YglCDJWcc3xP236e50zj996Ktjc7Dv/k7w8jcYwKIvnF
2cu1ZjpdfTLikXQorik/YTPD8OKRbi315UtdhfhJK7i5qKhQLgmX9Z3Rj+MRhB3tdL67TdWCECk9
GL5QPkwDNjGjw6FceucZyev8C3Ugs+VNRY3qpQ3U39Fj91NchSO5tCayzyBjH0tVOrTUz6gSXF4k
d45bZcSfD9bvcZtVSTmLESi0PAALpzko9JuBkcYJdQH6d+qrMO4trjpVAsVRtWjPMh92Dsbfb6y0
zIb5D5ywDJ2TWWcZhj/4ZTlhw1AAv0HYHwx7a8/JjdFquxIdEiIRNKb3WS6xIfSw/1RyAn41zGRh
a9HY8B6rIbtDHxhZb1o3WlGlWYNuA90ZGGkHC3x2AztBnNfm4fiHa4jpdnecASz2EYwQx33QWy0N
9vdEBmqSbGs5QYZD/SHpK+Or5ELGfjSfzkyAXaBeM+B8beW7FX6HxQJezpVbgGCHuTE87UheKVfW
VR4psX6wXWLaYavVsIsbP4GphJYABN+flgclr6YJ7No+aGpUDbuLPCHI1Zvs0THacjQRnfD8oLeq
I/FPH57ffywDVVHWlCzZpmhgrH4mFdm4IWEc15EYH6grkOdaFeASQMod0M41gAK7meTbEcwIYbKc
XS5cymaSGxKozTwT6z2hOMBE39PB89+bh3R+qpsgZsGzqOO7NdWJQYighnMyhMR3xeelQdf2AKz0
rKL3lsaoTDTLHkIMJeSjogePmlRpFRpOfkWFU09xVFOm7fX1wnSHXvFeiFt34q0DO7wEsrs0/+r7
XZBS31gmFWPTYSrpCVsAQUix16R7T2jFYfERQUeSVtzd7hS53GQ1+oYtWSSfZl90RX1byoRo91x/
/88c4ZCYkBBNLyy6Wi2aDtV7lQl0nm9wbh+lITOwzYa/ta61PMWRPx9AU/UE8ejoUOfLDjqidVke
S21UVKsCT2wFUFOmRXC1qnpfuk4jry7i7NdOX/utapU2dpVVQH+/diXvbWG5asDeQ218OyBsTHoF
qPLrIXyRRbfUGllW/ewB2CEUwC8sBBiOfHKL9yrxGUV2dYjEYcRaCg/pF5DWh/wVazUri3/XMTJN
IMnHLzlmm8JHAk1cfcrwCSMLHrGYyAYRYhFdONNTiTI9iUcEYTffPHSGlDMaM9jlTCmCL3YJDmnn
Xi5tYYoBbsVKGcJXs5zo3kEBStSJpeUc1KGovkafTJd7ECMJYknn44JMv60H99W4D5SUP0nZli/g
sMqHpiLFajT/VHZbpG9lqondAHL4/xfnGVRAuWc1rCS1x0CfPQhGHZU46anIf2ntcaBDT6jEAAqT
Lj0Q8+k7ajvKEfC1kCQaikhbOvhiX7oaSEGpWmtc/B5ymTW8If/4SlWgvJdqiU2MaknR1kNEFKSS
DJ4aQHBkSAw/QzbOmjItL42rEJNAszcJxYUZr4GSqob0FoKl8bI7J6jToKQ9KA2UjNT1klja8vxy
zPj1tcO6pe4msPiwk41cnqX0v+14P/mrq3ikk+AvOdmBfNaZWJOvEaTlhtHQKwnocm9TXqNq2kL2
dN/OEF7KLvp10EoyPQCxcobI06lfSpYQGRNbyLKqWDcCwSTQEQVYJEQ5Ett7MhEhVMYVIdMs38fl
WeIj4312MtqGMn5rr60NNXrvrY8javuk6imYrGbxzmACl+YdK4+HJNXpLBhd6Dapzua7Rgtfondc
g4mSMgwDVbr3oNj+YtnMv1aDnTJdHxFZiia/9u7fscnRq9Nu9LCVVsKVo4VbI58mkhKqpHLIkQaA
Gd5oaCVIGc7j94nPr3OUPLVb1qwLSb9kofcVVsEY1VbGJ7Sb/lhGuihf/3AUOasmviiEOuAa7UrY
Gg3saPZN2bPy0i71t9pqWjZobIadWVUb9ChgzX5xFz3e6NQ+bTXxTSgvU2+bARUzR6yyg5igwAbp
zWkCS9sUnhWwRz2e0Wxl6py29bAJj0Q6jgVYbEMbZ8m+oXXRmLdgmEXlYxLBRJwsEEY7c1/8O3gz
vmCGtWNfdbnD0c85NPU+fMFoRSV+oV3eEj9xFPbU1kriVyExBioDdmIaU2dlUNBd2NLvnPec8+44
eePOlQBO+E9Fpwn7uU8SqAMsKxe3wyFdqA2GddWtkEoZ2YlYEHApqMiWN5uVQeUB0VXXcro7WPIl
RyqIoGVRyIwqy3Qv6pN063XNRb58CP4G+h13nSe+3UxmsBaH0fv4YFyxBT9b0XrD7Rm0dapatBU7
0w+9J+tTngobVBWDr6YtKcRcH/CUjmURuiJn1gyZSZOKC0lKi7HREHLq+YDGp/V9ig3gS4Vau/1F
qjl/4sUXW9GSr3v2n1PoHyUKWKEspV4bnrKjV7KkarRPCNsa6rori77706Volyo+BUetjfcQgyWn
ktzEgWdNrNpEx9lU8lLmIn1KiDdbX2QX1L6kBrl+4t+AatU7d6pQSi2j5xXfeNZtjbK/BQAFQJmq
JzBZe3gXe97dsMpr7me0vSWLv7G6Gwm0XXFabDlo4s99WIpES35guU/sBgZdlXMvZC2ZOhAdEtYM
6ZTX6hZicDwhs4tI8yqFerzeqUfGS7Z2nbkuQOSizDDEG0mVJtbghWPOOVqypHySeFQRve4qmA1L
U7x6r3zZhbIKUFo37Ajuw0UQRsv9nYzYIq6OCFfiTdZZa0uFSFX0ZsqGKkAECrcfUxhv+CcfLYet
rKoWprKYtBzBakSaczvUe4piJGo9bPqrCYtH6m908N/AO5e3O6heDAg+Y3o94M+Wg/zR5r3dey7f
ZbE+Pd3O6UULLl4efgk/B8JmkzcmUC5EqSulO4Xr0IKJMhORs4Ii5aqRuaZxXCPp0EvsRxFzQXZz
sLU/iAf6+6wElQBo+lchhxiouff1FD/TxjCJdY4FGk4ZrI5afg/Z+6R+yB+VpPCBhI7kazY0apT5
/61fgEy1+gjVJnieQup6XM9BJ37eX4RAOD0aafR9gf4r30QUVB06M++tncf7mXROjyjzbgvGbQ0X
j7TKXpXT2GHQo5moDSn7XKAgjLG9lB5ywioT2dlqh7arzl7A3aL70lMEBvJ2FM0yN5lO5B2wyXBu
y7W7ZoupF7eg5lBnr6MaypxKtoDCIoOgyB1wUTq8iE0LM850WqC4BlO5b2piR+Kxszyxx9WaDN6r
sQ5eFppROb1BAInFD1tqDoNILjs0gxf3sEfg2fGbTATKEQGE3/ru80wsaquVc+NYdn0/3cgrD+pn
jwscQKTpR/lRQeDJ1RLTq4IIvPLIV1qp0cdIJQM6pDkA8VU9WUAsr6LwbwgIJ1kj7UlaLKsQ/VdH
RT1R/hbx0lVbihvbUnCi+bWTpRK49j4aCJIYQbHIIDUv3C8KJSizTyp5ny8Nfa8erDZ8LS/Grtkd
WjcKavXM8c8Eabhe5dtXXSg+wr1PS+oyRMguVEuzjkys2VhJAHJKxpZWCZ1TkW/UJtju6MiCvE8Y
Y/bYHk5wxeCkp1gbV4RFCTnXS/sADhJj5uTnynjbSagBii5mAKhs5OpMFOMfYkH8Yb+iap28CimN
u+44OEGlDC37kH14pemjoCmPyUVz4T+lLqv+/9VOz8rvk0S5rdS+7Fcf4hwGFNNAGQpDN5J4DBlw
zpRRs7YxR8QNA4VF93opM+uQm/OSVXoGaXlJrapFTYzBAufgIrJsDS/l2T+rb10UvrTEoVibxsBZ
tngmBh0AgHUqPOqFkSOhriDOHhb7MHzSLHIiEU+ka0rjMDF1/Pq9BpTGiVzURz38x3AH5Ot18ycY
KlG2oS2ZowCw0OxiFlSAhA4BdPcxEaTfG+gkFemS9t6f2p7wxWgocSZBOvuME7iozcS1klXDHi8m
vh+5e25/TTbY/8mc1iue5kQIoormH7ycm2pJtmM2FSKYJlgdgDw4rBd08YDBygyc63xd1v6WnWRk
IHG2a2aq4dt0nEc/JgMCIZ1YZNgXySX+VUbeqIik2Upoq2g4OYmdihRMHFqleYFL8DXFPYonUkS3
nXvS6AycEXShA8O1vQ75BhyKtHO4GoPwguFKXFMwn9DBT1rzZSIWzUb52ZWJeDTpMwUGuT6rcPEM
1wTiHnZoB+Ry5XkE+pyAidTEIclQw49SI5fiCrQvaPKkxuXUAK34l9eZmBRDFJ0M0um2Ynd5JwLp
pRXX+6UEatcf+pdKypv1Rzqd0v+PLDmlkRPra8knlGc7tvq9cTkEzs4nf3rSKpjinT6yNZJyEmNl
SuvVxAHRpjkno4trklTjZ+zTmfxUNz7lJzO03rWpk5eAa98Rk76GsviHskY+4L0FMOagWvIsJlQn
SItJya16nuj5lGfAKSiMgawOmclkCzsVhRT1pTA7Db/+7JmzptwpGVm49qh9OhNboWz1gTUaMUf/
gkEuypVMZIAiLZVmRvjdkDrdDevJmR9/XMZ9741IXDfcGF004IKcWkT3dtP3xnetQGhZA+idefPA
li3XTf5epIReSbDNO4YVVgbhVUx0yLmx7OUkpaC+PB7ZRogWrWxbQ2og+5Mfbbtoa52iUv4m/3XK
nkH7Y1/6Z+XO4be8hKe1THtke1s3gcbOQ4k51RCVL/WFSc5vwfIJLpsMHBHm5h3Zgm4GlDXIjylB
5V+iArcmwUD1xv7rFf3wSHJPg7YxPDbVT5VMvGnN9Rop7DQ5RitUtO16IfLjhqf6HwvpcffL+8EM
WBTL6ZGmLk+Wtj0uAOh0DFfjZlWP0YgtBrgyvgvu+BTZVGwunohWVjP9FO2mr0PlUMQjYxmuaM7m
r35LLcticn7h1gw9p7Q7gx3rAj7a8oSMJILfUE03WNPX9UuW6p/1pJwkx4dtm3yUmfhmfW3kaxIh
a8I21Z6c2UnMpPt+UzG8JxX9wnv3dy08UeIM7v7ILoETEc+soRAxCMqUp0H4e7EpZGqGmidjFp7q
nSd3AQPe0os2tFzpLKEdU7fg1zl8eqKRCFL2xup4OFc5zikgwC9Vd4jQGiALMIERNrwKoPcSPL4F
41yndr8VBHaJ7iEF37YC0iauqyCIGWbkjs0rFQnrVpzX3y1HxDIZTFCF+x9HJNwMKO13Ll/Z+23v
98gzuj/8W1Vrv0RXZJftcWjmzwzHFNz9Lq2XdKL/pAMds+OrS4FC7uY5z6SPD/p1xlQ3lW0jGNIo
iAHvxiWEK1vNlzXTPoYkLaPLbLmFRPXqgUjJCUJdBq/+hGR7jgEq+onnR9oMCcssZNxAm6cnUQ/s
Mh8iFeAk3r18uJ/buFSz0F3dYW8JmOlY1KY26uqjseURv5OBniAEmonqhY1l+XCgU4BDj0fs9nHv
uGnkUgFinyp6TH8mZenm3KKn3rpZ4yWcGwkbl6+NOJoNgxxeU4UjDHQFrxpPwxg3BoW/VI6wScnC
kQA+ZUO1YfXO7mZX+Yae7bVcg7eYTlQqpYlitEyl1KkfmRGK4HwwXa6xPUGLwYeyQs1IsnYHNbrn
n4jDrzYvbo86LJnRasZxwdA/VG5PZ3rlLpjXww4Fn03gmUk5XpFksOWuB94Oj1nMtTGkVDB+WP85
5JyXqGdTC+Hlb0DTJgm1n61T/Nvpk0IVvoWZ/aErqoQYhaxHtgwHf0AJTqUX0NvQCuA1YBPrUbLJ
W39NugQ4FErDMa09YO4ReZ6lodhXdXBSk1MiBURDxczcO36GfRoPwaYMB4GtKIM4ciOU6xrrQzaT
dx+MmWI6Sf5fDJ3cyE6aBW1XNTdpYJ/EtPpWuLB1iQethvnAsl33msQOcr3yut/+JG79BsRiN4sd
SA1AC3IT6I/pJcCk03IbnKKEvEq5Hub/nRsbAm9DRcenLB6RIfr1DHSs5oOjBJ08JXmU/pwElCOE
MP7msbXB8jDLHlPckQTzjNn2O4aQRf5I/itt5L/6lJV/y22f0Rl0/kD8oILMAUbZ8fPYJgrykUtf
qCbxek9xwd1nV5kMfYqao1mmZEzLR6+eBdJVeHCgQpeKkD9+Irdwu7uJkaL53S+1sAjedz2JVCvi
Ypiyw9UHUY9hve+xXFN2wA6QV6uNaw/cMFXuCpLtkD7hnpZICm6PIt4kBTvDDmT0wIE+MOYIvziP
iLZlHnaPPRH5+ZhERexSqBBQYjyXfnnQniT6EBYbyx2odMFUWf6cfZz4xU02jSpofeLscrxxC+IQ
MdEWZbIbIe8M4JJYxSHe3kXfcAUyfhuuv9YD6p/nBPxk1sn2SqyEiIZ8762t+tYreuEM+U5IZUQA
ejYqyegOh+Ey5KNhsPeHLWBhEvMFGrQQwPCvdJiA6DOlAaSdFOqVCys/In07J4heGPR3PCV9R/KL
B4mFa4pbv7zn4+IwKslTns+GD1LHf5otRRuPgU9K/v6zWlJu5sVXgkrq1Kg7iwjtJDeIEbXeP36T
2FMJ7sL8rS01d2khEbBLEALdd/CaP9lV52XtK1c5bEtcht+pWWs/YbKBXtd2EHPWgsLentR1tV2e
+OCaoSz4S3zzY8WKRn1lpRqAkOW/0UtZKz08f6T06vu8cS22YiEqXWDbsZM1hMnMRa1+oYm7nrWQ
Bs4E7pynZsyddoo9zOhyT0Wkvgj7Io/cvb+B8lRFn3VrVuzZ+c3IIjPL16KGdFQse5kfBu0d27dH
Zbap4gUY8C/47MgRhoTa5oBtQfk4PHQAcJLDZTxzLr9xJKk8+yEMF/DH+GLkUIR+Ru3oN5wM5m+4
ZhDibuq6l4aiRCuGKrlCjc8h4hBbjK5gu88mxQdx0elYzsTf+lfHe+YwpHc70lWUdXul3rY606cm
oY2wytRKXh+p0T45mkpu+Fdfc5Zb0v4/jfMoTpyxELf7MIxdXWfyoQXfamPwHl62bcnP0O/JVkkN
JwgLbgNUDUITKJBrY31T8gNuKkgWfcopLkARX4sFYhVAr3WU/ruW0ObDXbrmTpDENteWRoBDpKfs
x+HB8NYnC5L4iAio64uIWeyozAUn4Em0Wh7+A823fZQIjc9tB48kxwNJzrX0rcyqf5LTvHkkixAA
U5HxzIjZlk/Gbt+bt9JFJSWU3iXG+hQw9RvfYJLktSiixe+kiTkB53FcUE4xFQqhcFiqvcfx4xt1
9GOT1S5/g1qSGwcg9wA7otLBEKn9pX4ChC53L0ntwNsawuXrXO3X4jTR2tYIupdU0vOMNCroubjR
NMwV9j7wU1+rpzV4sHnBhmdpjIkESHuOAe7Orq8Eye90y0vKBgv/3XVhb9x35kIT6UvpOxFS3u+A
xEtS3rJhccBPQDYBDkWsJnAGdmajJ5uyR5ktrUcjy+I04rRN2uzm7/3sLv+DAHpuJhkTaTGQIESQ
GAW53qYNuylbibpeuN7PF6iND8r4S6Bth8UG8AAFkxEtMONO9SIjAQDPPLX1nriuDQ0bxPfY6DTO
lAJoRMHzjLRvX7Gt0DgmR9JdznLOFiVbPxIShLDa7UkEU930l4MS3NzkQfvyy/0jtaCvrj7cIEHU
9AIu1Jk+Rce6yRDHYaOOgTx3Qaezskppoz3KYOOJ6QrzxcH7tOHEHXa87DxrQppYjtdGBk5Oz7AP
avHnPBwn56IItQ68Y9RggYQpJwV8d74MAc6mwDtSzgJ02doZBTp4T+51tujTSFuW2TN+likZ3Ovt
qc7neQDfS9TRc1GFRMnbB3yzajPfvtvSYZ55TI4olBSjGNHQFYWegQga/QLKq9ysEtJrlNlQvtca
NwwLxQKaPg8kOOJCfV3cnf3lyirz4i30gBmKTcb/DlRtecv+SXaoYYGLBRagnWZ13al1hOyQxzFp
4CkzdcICbrm3Inr1az2g2XcrxipcvOTml0wFuxdy2XRK9rZpYSl4jrQfPdcY/mpTRyjn35UKrEew
PnO1f9EnPE0XpN9YJjYZUpXZPq9qdT3E+/WLAIwsl83XmfZqUJfk8FjnVc8/uBBcva9RMNVzOHjv
AYPmqrWG3xFhNf+HgAbnqgGTJXPd6KTK+uoGSt54RX1GYOZUEmlLpQXo35rZ435ays/SmCwueYmm
EC0P3rG0j+MOr75NETeSZDa1ewXirdsbFTsZVx+u55rT9QofFfgUqOOhS4l+HWfOmOCViqHLdr3A
SdxQP/N0mV6wsd6zDCi3XZ+b0/71Ybj1STPOm/OcYijZHDbsa34IKQNzwkKn6ZrE5VJRdcqmAQpp
hs1CPmvgiUpvn/mLyeD75sEHr2PKB5SPRJsFA3dGpKXqBCPeCKZ9ao53/VadhfBc8toNj5P2fPu4
hnRQL8x/jnSGOOFXsj7amQZuC3hcBkpBlai+31qerZGvX1Mswez/6iysphLCzxjFbgwSieXEKxm/
ZLKuYqgLkLFEq792wdBa9s1S0+/ayMe3pFyJ1R42ZXkZGNyJZFt/wYCPVoRHzqkt+hi3m0+3QdvE
OB85ihZ60nafliBbCapNgKhBTePh8We02F2VIwSb2yP8caI/l+nZl2e5jBp2JAfViAPIIavrokGm
33/nxunmsl3WOlngsoHCS0xOm31GkgX3hjC/jIJiExVnZWRA1WgvuwqALEQAgs+S/I+LhLDOAc8l
k6cpXbhPaILpOISAg2RFqK5EOuKQbK6N5Q6Aup53pWuUNVb6PTASFkA2yDG0LDNqBkuu7nBiAZ3D
2DogDP3wyK/cnc7l7lRfnkag18zO2T3C3ytB2F2Jxxw9VV5IN1Kwgo1JxfxZYSHnM/ZZ5y2Xy2BW
W+zNvNVsATWSgqUyftBuye4z9ADFK67vshWzbwjLZ3eompg++QXokVqkDTjyUe4KACKSs4HG06Bx
8znAqLsDA24nAnktb4PbX9ED3mdg8UHRqHWthHZYaW/1lThkvw12yG5Z9xRJvutDr5ycLvoaEJvC
d77yTtgizS7SW2mYUZ8/6Xh9ILetGRhaetBjB2ZXV+nZWkR8ZuRwYc5s8/xqHRPb93wiS8qT2+m/
n1u5CDBM5mmzyt2pk8jqXI9XQZeM7LRhb4rYs5hyg5sjXNJGiYGi2dPi5lRDv691EM5Q3JaWiH98
B+uDXRINFhdk1H2zSxic/nh8xKWnwxJkBzYXzxYahn1m0A/mVXQJSs4zQMu9Xf0GSOv93Xte61Ou
GX5wMwia2QgKk5HzBUyDTUYsRS9kdLPld2Jnd4gGrWkmG695hh+TSAG5Xm7zDhrKzplkJcH3Z1wG
8//g9kn3U3StcpjQtjvm8jURNZyBRE1cXr7XkdtUP8BCLVI5ROVPyq6B7H5XyzqUYo+RLnYfUyPu
Coe1URxDj8JIGdshKaq7NZKTBTL4im1iCmQ5UPJwvxuxmVqNbVqjkMpUIN/KeizrLyhXiVBQzljl
6RxB3dctxL8skwN/vm43/k0RXTwlDk4j3HLowXJ3Yz/9cmqhnsDHoKYKBw38JoYZb6xMinQW7WoH
Xl8CrCo57PMhZkUXiuzfVXfZjc4cAffr+XZ0dySaBfI2rYqqUs3mQsoguFSb5gSEEpL704ZlXVao
SYfoxIjSqd7W+QXNsbIaFBspOne4G+NkehFJkESfoZWTbHG5v0fde7QuspmE3SL8tms14QFhkrNh
70mTkJs/VpC+ZTUCR6+P1Sz50X98WyIa/2FMWxe3AosmbmDcsCKExrRdwb1bzbnMSR0npo8DP7ln
Jx5GxphiJmMQPf0ia5cKJqIrAHeZj++zzYfpaOK4Z7DXrWxYHGkNVY7oAw+jpk015DzLRMDn8QBa
3gd8XSWPWVosffjX/019hBYF16bwgTFsyVwyBjsYNs2HW5H+UvsrKGSOCiwJ7cVY0z3pasS0sQPa
H9CZEAnlDuEG4lNxR3ID+qhjW4cVeYzFJvXg4r6Kv4ANb2OWWA9Nu7fqfWZTxFG+6Vy2jwdWCMjy
ZJ3ay6cf2TGGov4NUI2YzmV/ZOuOgrsPCdAAejpWQ6UuaI7y5UeagSwGA0ITkafIONKTlsmjGxNM
oppyTTrsfQ8qytAMv2l7iYS2EYeVK4uppRVnQhVrmU9Fr2+HLHR8ITIwgC3gA8WliO2ZT+rDdUJ0
NS8zbDIhPoSAaG/ZNK10H5huLgpB5oELaBSMeeFj9PLmahMTfiy3zNQ1kPlYM7pDKgkCoYmqix5g
Ron6BCh6rVOI2ybgTOU1irg+YFIhU1G5FYlDHG1VKQXGF+CfVuBQ0HyGqV1cAcOMbZpOUyNCeuRE
WSepGK3es7uXyYFDs0GU9U+jHkb41C+PmPPTnrF9SYWf8LppzE/5DXTmv+Zv0ItbjQglQzNkTsKl
aQIT4PcJqT4bX0857qYvwGFYfTwzgZme22lQCndqoWbLL8YmC3GzZXD5nvA66CBKmHz+SNiPu11A
T+MpoMS7vKwN+YFUoYreayINCZ1hdc7xDDZA+D/VfS8OTBaAAl8F36UX9Al4RkEgmFbddxJldA/s
PIfHObuX8VGVJT9qnNcG0bDNGhLtXtrnxIDW0zoXl62cPPBol0E+f29S9KVjgSh3QsZlfmYFMFTk
8r2msd7VKDxoFHc38/HJs/0FElc/lCXhm9Y6wmhAM8YXG2n2+UjKA9AtmWY2itFetsR3vAbiilce
FoWSHhDCJ1G6ngobKuDkUoaXpQS8syrslok0Qk9PyqIho8gZRa3NaJ+dpQBhOEiF0ugti1ma4wnY
4AoKVRNycX8Bp/kGU7q8cRY/Ee/XDBWl1GC8ZwDdIC/biNSSrENplRbH5yPmwJdO2o2Uaz4dCaiL
FY4Lheh1o4jUnx5nPoIHCJTWLn5fOr3OIV7G4mF5MfqZ5JLsu1cNZ44iIfz8h402HQOx3MF5TMB/
iTP6wwd1xwlTgcq1q4yct1LcAGcfFuouhEuOU5CTds8nzfrOFG6UmRNXLCP9JWzyL+WwIGbxUCHV
cwYaOT8Qk3pMB7rdHx4CGl3+qf0eW4vCmTW5M/wW+dILUF+5mMPvZMdPEbo7Jh8X0QXDeMIJNFE8
WQHGNqI6MjMH827XCXZdckLG7YoOuFm+B0JSnBe3MC4QofUtCo5AArJOk2FiV7d7Xseq4TVCo44x
S0RNdlzmpAZpvmhghTkiUNeVTEdQCC5DeHPwZ+fKipb51etHhVPnB0kKOE08vGaXztfg9lYknq44
0zMAnXVFyLk6lhEYFy1inNM7jfDPNl70ZSpwYEWoI1XOloDACG/b2TcOpJ4hAUZwRLSlkO9cPfor
sGzrcOQ3BwVgsxcoOXqmkSbbZ5mBtCuK+3rYnJD9QEqhWuYyE5JY1i22iafgZGkI1go58m/TDxsy
F5v9mzF6LPC1mY/IpLsrS2taQFSi+rFedjIFNTu+tg4dUTeR09kCoWt5JEWHDqRtR0Wy02DOpSzN
TekKBt5gXtq2VQvTJYz1/pdTzcgxY4c92IsjvzeI3zEdlumif8ufl8KMrpQefN90FzHvU+M4YHNV
cI3sXoycwiZIsPfK7obI+vOUWUR+W54beTDg4TSkgfMBdrsBFaUxJDAqH3GP4VQ3sb85V/gZg3nt
j18FgIcY52NJN615wE2Ybnn6F5NiDWFAZznoXo2RLb6L64IHdDniv2oufyUlQo8L7Y+R8DZSW2q2
wTpFdsE4BHjbJSKjiuGwoh342YLMTb2RNwkMZsVKMzmQCHTpKoP8amPS5LZCmM2eV6zD0ntTgRS2
LB6lPZGvM4KIdKe0OqzbnM6Uf8aUq6n58Lg8/56Ss86JpkZ+PvHWjZbP8qwVQK27A8o3ht72kXwL
P9gL09lZuF8HjMhiLLsMfEJT+fA6k3zJfepsJQd05LfN1vRqhb1dyve2+1EsQeRo5yDvtAnRWu2q
/mdAcQCGYCi7Jqwt+vRcD8WyMDclZQUbgHlYvXqOdbGQ9WY2ssb5cRDUpEV0Re2W2pX8qjqF0Aok
sJF8YOW1bK/bz75PkCbmC/DuuQQGUeDE2KJ0PKwHmW7pVVPR7cWoL5Ph0dgasWFaB7nZgiYEBzUI
AwmwU/AviLyWFoesIUu6SPCD00A6yJfo36r9pOfFtlAvglwgPf2CQSCPzLFs4w8N8T7TiJtpa42T
y9DbhFsomsbFKWb0STdr5ndTxyY34QUHzTlCO5DsKRTaZp5vw5gjzn2TYwRM3PEhhfwuHLhxjRoc
hKx4j+ZfZaLK/FdawlCagwqUFMULS3/qU4qAEbIK9wNutG8v+WJQEz3DmYmCpTtTqahFayzp4SAI
uakqWtuMEdQl8UT8geYDZhNjP5a2qdvpCn16ufTAC9D+c+5j/Mt+gwdooRUizjXge7BLbosXEi0y
FtcEryUrPEOQa7pgORZ6weUqXSbPIBVAMiKFq5LoWSq+tErlL79Jq34xBSbZ4RoqCfBQ37Wg9Cf8
hPcLWMb7efNuPOF2ElfaI4fJ1FkEg0fxSQI6zJxZD+HlXUXTyp4ZOA6pvf1zHktDjfV8euFTUurY
TFt5pOp7TzqxMhgqb94BgL+aYMTzIx4gFhaufEXLOOh/165RkVbq+EQeJCROr6BRUT6APRes4Vfa
C2NUmTm4B2oxPflpMO7E9ozk3eQfWKHpLv8FHwjseEbUwottsm4etg6nYa55io6glHMVop7r2zMY
03T6PY3MDKJcK02PLKGOCr36nh1W38gsS/pnPp1jgTLX35337VmX5YTgHLHBJas1mhO1iSFYYZkK
HHzUDZ1oOahlW/t1KVqK0GhGxZ1wSmXRQmvTAX3MuoIIhD8s5k+Gr9ZdIGjVh1zFKYUcGlnEp4wV
Ncgxc6q+cUs2wb++f2qIQp57ENBEZQO/6l9C46+yD9T43wwG6WO2KnHJI6PNb94KFnteGwWMRMXG
kuFDBFMu9LBNFSSe2CybT2ejBu8HVcxKPBTIqnr6gvdvj+JHZpOLWcztdM/LbOw0DKXmdV2vioUz
IRkGHk8FDKwwaJhnzj+xc6G3mCebt2tEahRfjAMx+Spq/QjSr7wybwVeo0BDhlUYWwgvx6hNUUWP
ZDxFUgsQ9ZjxhzJQlcMKQSSrg1iXIRUncG1gllmBDoPbtvLpE8h+Ot4enRU1yIA0/x4hAMdlYtj7
pqEcQR52NA0hdzrsxuEYsw11f1sjdroJGwRguexoJVEjrLXxTZh/FPZWGjduBRN1gQ1hAs1q3VCa
vbe3Hy76xk/WQtX2RioeVTgV22l5u0E0dHo7B/UPG6d5m4KsjuTC+/iaOK1QUCjAhAIrP8JP53ZM
rW+cBYgDWK1mlhbGocIwSgS76BAPE9cxVaHnoyh4AQ5EoYvK2YnabkENbwDkgCxrNA3nP3o6iyLo
zxiF7FKTqgzEgtOTyHMcMb2K08E08ioN5nwpi1LzfnfevHvA5ME3UeEgdj3jmvMj2G9EOwchwvJ6
oT8gErzLcChlkKCFbxrFWKPScyBjJNzd8CWmb5LTFIn/b0ah+hBOdIKmNtoxvzVPmDtXT4pDtpGh
6ZFG4Q0/rsKr3y84AfGY+e8wGxFxQclCvLPwrjtFhtl20/WQOM7ClFBVV+xS3jCpuJGOgX82QzZC
djP9U1N+I6FW7HZFOo4+yd8ZCRqq/p2tVt5oAFA1hTHRIWWOUdk+T+EhJ+JrMeFIoaIrf06UQgE1
VMwmFPyYsIXk8jTqWBAoXjCzUWd+NePdFTNJtBujCnUJcadZ+n70LIyO2TwdeUx1Tjz2Z8L80BdZ
Mhm9IY6hBpEKL7CWgeA4t57PJTCcJBE/aib7wocl1nkR4KIIaGAKdqjqh1XWAyXmiohydYGDm85R
5yL0ORgn6YAV3e7aRIGY/zAmlRwfmawWtvrHiY1KUpxUZNh+Mq8V3Nz2bQLa+OAGJCkYZmOwZoh6
06+rPjMqlCdcvWu1czC3mNWXP52WGu4J3IdRw16XJMmzrYETTmmUSskl+1Z/1S8IAtNk6NZkR1oT
JpRs6gWQmm4KfhzZbE9eiRPKY3glowmlZLx0F5smzHUQKl3Jg8z2CYdUMWoYTG+6Ee0LnvUaoxjo
UTKnmv0NcyZs3CzEd2fPjJE9d1P/H8iKCLdoctcfr2CpX27PXqo2RQ/Rtr1Jye0R1Vwo3/qVDQfW
s6R3WtpZz4yh9xj0iedcFjnD0qTxTn/8Ppp3fedrjqdXk6NAVuykuA5S3t2YjuO9Ur7bKuuO+oPB
FVIU5Fw+wNXugxudkXpmM1aehVMIoshtHRxT0I7jclTr2PDdQf4wqjBXCEBoxf3ZVTD1G5owjQpH
932/mLAcTASGQEgzDj/ZITzfFtPhOYp6/IyrgnZwY35CBEd//MsNIn0FfF9OW3SH6NRBroMzbw0f
WimvVAOrUEusCwPkBFmiIP7imME4GBEtlh+spAqy4EdMz1ggmN0HuWtgToWz+ixPuSKQKDtiCqut
SKMyhVTkJwM7gW1XAFIxoFCsj0fglVD4z/0wof5Us+ylOIGWhY2a8J7zzcO7jY7NNe7iDWf2k37Q
cKwYAy/aAre9xTyOoICMf9wgS2O0lOjs5ZRYZ02zMc89W2luDdha5HleZq98ZB1uWSckeQGLo63e
reMyeMpIoyWh5p6BHdMASRTJnUzB3SuERJHyxJifrMCRwQs9VnUyvd5e8mWPnFC20nXK+nI1QWkb
j5nUATZwNeNIafa9hubC4SDcsDC2R3AzfuqM82YU7jHU5B4JlOUkuzbqf8Al9eyATCGpBQbSeeE1
sfYDbBgk707dPtjeURCpjZLXHy+di5MIL8uXyllMFB/Ay2E2F3XSNQr3ROXY02bpSoeRgjkaXmp6
WBraPi1fAa9qCsz9/dmXuopVuQVgDjaWp5UmgoB93xzt64MSDQycdejt/f4ggOnMTSwqlO7cHcBf
BBm/oICUBGviy4c5YbXUmO3m/k7CmAJ/KoSqYUxIj79P8i+B+jTeJJAuNyXPGoKiA/GUoCu3LKg3
ABhPsW/zq2VfbmYCGlLpwylXNU26PeALa0KyeGlaMfvBQ2HMN/cpOkRIwS+oWug4k4YllDLjxMCt
dtQqf1u/frRuXM+t79EuE9kLh/B8eb3IhabJa3Sp7wpnyEpucP+TggvgfRoMKEiMQ1lSHFV26ACh
BM7yn12FB2mjw5qFm21c/L3pLw5ibTM416P15QkQJuqxFH/27kLJK1yCCsKVUXLa5bYD9L4JtVYQ
LlSupHTuCxzfW2MoECSgJbJL6Z+PyEMeKByoT9dMsApIfAE4LzDZ7JXL44UipbJjTSJepRI/dZ7i
bs6Kt+TGepy+iZcWAcHFzciHdzRiqQu+ylwRpIy9XPN40vIw9g/dsp9eZXl/e5x7TFc7LI0uCVgw
ziLPcm3i8IllL1tFSeYB1ON2tREZIZWlLeTN354+e++bAhy+0DANdxtNPfQ4hhKMbDNyssh5ronf
NV8kbxoVm4Zjk6y/CoTKfC7md20JtScL5oqTckbSsNtL+BsB2ryyiuK/6+5YzjgkTvxKE4hoSa28
JQGgczRTYCjejVTgdCqmZRAU/ZAtXGSnKpgnWb6Y9bmvW7FzGLZEExn4xXP1FD2t4l6IuGt1vd93
m4WwCaOeOaK8RfYRb2q5kwgVB4F4latQL4heg9iiIlPGPpuZ+cOL+Exdr75AyL39u4DQkPYHTl6n
dltrNhPb+WAigkbvtBpqzOwYj/10E6E62lqv8sblOMwDKL59OAvis9m14O14yirmlrCMJ4mhudj4
+pAMW17+1iAnkvYpw8Wyo6wtXrrxshgOZDyUleZRupfdqp6yUIraj/C9NKZXOsyBtyhEzmw5zztE
ulj8W4NHv+5lLdz2FKFu2f7Jhe5Ea+ni2Lat2bZEJigEnwqa3DQAciYXHoq/ejz8w2Jlyqu4b3S2
+YT2pwp/Eirhq1RN78xk2u3jFkvhmeTI7F+Z6K5/NtY6E8Cz5gb6/PC00MAgBMIeh8s4bMA1+2d9
SNGfuPVasMGE6JYJFgEoEeKxnnTylC75EE0i9X4sR3Kc4gJ/YRWUPWY2FE1J67ZIEZa5Z89BhDXl
t58LLF7SQXYdoA2+TQvRzZleogk3s0/rpmGFqo+e5qelfP9YzNsy7xN9p1Hw6XDx3UIEEVgJlFjB
Cvpa3P3EM13wSnDtJcrSKc/K0H6Bl2loPtGFWDDxgZJtMOQCxewyPwEVwa6JPCd1YKp4Enh1i/0A
7GJUFTizc0DCZ4Iq2hNsgpnq58ZFn8Wyqj9oqC+6x1pLvSGcTW69GyoGs4BBoh1jc123jPCOPxvy
sYaxauVdfnW0NrHATJCyjzCDo6qE1q+osXrC8LmyuB++NDqwR+o/5nZzLogWQTNUocTiq7gLamxW
cQjXrBET/40bzn361tG/G5c5YQjESGvCdsfjyEyBiSC93YRW+X2Y/bCokHRda6Jlor3nGP95mtUq
gizqnEBksufjrlKg+tbd+GOZ02hgkBBRHWZJHPQ73/qwOGxBC7NIaxpA8iUF80ksK68flOObPJqz
qAriCZxPIUcE2wq5CtPnnW3xW/yIullIZtNJ17K2WrcE6bqpObUIx/HRnLex7+60L1WevDSyUQtB
s02QgCM32n0FkYD/VXILo+m2YpWjMLeytWSuMv8p/zkuwfI9Fsz5aQxAXujvgE5X1oAW+dOjP4HM
2MzJuyc6O6z0HrR+CZlD+MxM60MdSn9bixqZZdEaPoKs/48pWv7fxKxfsxfYYwMff/s3wQboyPEC
G9TE/ijsZ3zybWHCI2/9Gn6Nl2sIMObWk4rilZ6WnpPTYLs5rgXyrKKw672AjAgi8Mas1AZdVQff
dh+LBtIqb9/7gkcxOPSsiaQXv7E7IYxKE5Ej7b45b/TgV3WwmTLVfA/rz/m1KnfrdL2us6W0qxug
2Py5Civ6A2zq7FhsF2X5323Yf0VlYHs38UY9oYeGXpxeEZk0H2js1bw8rmTq7jKMRpXsmZ6ctTDn
v8coYa2cjCUq4SbZaywT4YeytDnjMdFLt6DsROKwxddoD13QaTqY1wu1fdnvFLX1PHfbQv1qVrZh
wVw/7aPyeLbDZUrzc2pspVEh8+zVjwGDBaKORGS28s9BkmBLbOH5dio/xr0Q+HPUtkgWKdejkZCK
NXAUC9CZp01mJVrp3cbiz/P6ADvgBwXj07EaRS57kl/etxKvN8H/02aqpiqG+FV9w8EXZYS42J8D
vhA4WorKc+Pyw+ql4GRxy/qI7oan9Im3x7nV9gy5XQXkHETHbmfC54s1emCFBFn5UlObDAfistIi
WuIR/qaUwGjrO3DfKlAldLzSnnwZqAhksTT3mxNGImk+xITJWh+kqczlFASY0dFa2YPmH30ut2ft
Rt+bsByPANjyQcBOCDoRxoEOCZq+x82BqhVn++Pz2y/x+9nYNaOZJfdmXxcQUdTCgCAH7EZ8hIn2
9xame/CRhJ4Hr/WtvEmeue0F22rmFunldmFcAQekuY3IAwRpqEzV0Woott0lnrwudXEYYmrQgTTU
yyHzcRGiuhsLDZ4xmcDZMZFez/pzhHjX1K9EMW00WFkmkHJK/pwrZD7iWaf8c1rw5YexbfCQ3HO8
hlmgEnbTutm5P7++pCWF3vi0wyBHFJRyZnTAnhdYe0mPUx1d4G2iySFjGIscexfPzXjr/BfCKBCk
So/xp7A8lYS1sGSCW6/v+kHy5BBD2v/dFHfep8TUYas1E46a/BBAytKm1rLkijbc1Aru3vY+feX9
WnO+BS2Mnb//6Qz1kBqtYYSI48QM5K6s9L2IUhDzTaWcpw8MyUBlGN6EU/4c1wNmLh5uoYgQEfQI
UfsieBbOX/QYQ0FQUH9eBgIn/gcyVEhgMzeageSzwvD05GJDywSEukXf7UYD9wdHttIGEEuiiaCr
ihSig6oCeokqF8eEhXKrpKIgFCJf3jAg6AcaAWV1jhJ0oBD6a8XrRkfu6QWscVykZRMVf3hK3TRN
hivzBjVdFVxcvzW5CV0nSmX/Z9dzYHMy+InokF//mUZZSDvbwzqimPUiPIATtXUzltV4LRXJWpOx
CFF3GR4OwJi8AudiMXXgiaVO346kcb73Ys8vvZS5gImRkF8fjWpQj7pV0jzOZEgLS4Z2bj9sVT5e
/DFqWGsvmW8tG1qXKsmGYyqFIVe6vJC4hOgxkdVzgO2Is3N/E4OE1OUm40x8gvi6yLLvxwqa2bBl
UTLHiuJnmkzGlmcFuOY9oDDUeAG6fAiGSGZsOODbNqsyvjc9vjspdf6U+8+j9Q/Xfc+Ow4uTzFQE
QUh6/Bc0kkZ4mkW2dAre0DnGK9uHrxd2LkK7xboKyZk6oYfrRY9UtuP41YMDkKPaHX4C4rFkMhUr
l6OaSwIMSJ40M3WdZ+buiPGGgyUNst6oQXqHZBX47aPY2j0gv32Bc4cf6HhHDU27m2KCgSV+pMO5
p95O2sp8sdiKRfZzUyEfjLc74hKxIAqvrkBh4GykTLai86aiPEdiXATWFMH5vr+vXQQsdIJq1eli
S/mD6F/2sdBkIIVf03oDM7Fg4XtvBVMxyEOsiaFmcDr7HvD5Y/GTPJqvNvP56e7Qu/60WWhBjKUZ
4zRpy6G0ucufgOftuLSZ0EjWje4RrAGNMa4N5hjT9DJSZkZc+DUws5ZhJ95i72rQOJq3UaSsCApR
HPC28q2O5ZW76R82EUMPsgEeikH3JxKmsAYbCaMDKYtTbdDFmVKWPUlpGFSoJVeQw7+eyJ3rP67D
moR8wDo3QbPNZWsN1KYJJCMGRjT7eFzIEvVkJLtZGYP7HW+mnEuCNHfWuy0GEAAZfFW/sRy286PI
Cc5YHLhDABrj9VL3CN6p8gBV7er7wZgCbtGWvbliiUiBV5ocHjNFbu1E4Kj/JhM19ph2jhBGUGkl
Ebg20T0Hl8wRBerSm2h9u/d5QwWB7lFQGiFQlI2Kfy/ROKzMPiH/qu5D86TmQrQzUoIaLCOm8cfP
fC164i/AZ8P28kPUOBcxKOQ0zTNm6I1CAl+B+kozGekCkZvDVh32vCQhmZROEZS/99P1cutWi4qR
kETaz9dshJQwscYw5EN8xL3m3dqDU1RpYVideqPp4ZFeg3cAntYW0KGa5gYRXKhlWjzLCUnXqLmR
p81jehuTJB/Jdkyua5cm7I1pGUgF00GvOe0DzvEQugBmayXZSjvXTAmV6fldd45aHWXWpf658at/
KZqY0g0bcRl4/X/2jXvPDvXG3o9fOZSm4P3RUrKkbg6coMf4cP2+fIuilaAE0tr4Y2nekKSIi6ye
zGHmmevGQdu8iQSYlkjVQxnVcegojaavHb2jIpc4jx0UYv+o4snM66mlWMvwoo0hsFXQY5v6OGoL
rieOzPPEFcMmBkXn2MX6S08qjvrkszubuYXXQZbVpUkvgC5ppY9LuRJ87c/eewZ1U9Pgt3W4Smtj
OZIwoc2ShMi/cvbCAdHqofrJLhJwQ8SC/B8+T7QOgAWxbHaKa1HPt6cM5INx/wyOFnzbAiAMdbmP
XXuvbJcleNtihdLSkhc7VF9ZNBZXOcuGiaoBYeMwR0oMsBiEPo6tHZupABfw4k8Q7TaWELtZIIVo
f0hNBy2oA68WB4wkUf0+FtiYp/7tOicMyRAjQfuWm3qG8hX8tO9jH6NIE2HLhyOsRXIVEybDkFu/
n6w+ReFWfzlRopj2Gymjw072m9fQsiq2U7RZQUXacrDOSrFt+7q96VPXaXvG0okLi5Y09OWywTX5
kcef3xu3dSIaxnq1h8mK3i/SauNk1iLz7jR+w2+GuzcKKMXsjFuGvxd1YOHGW7SH1fxQj1Vdsfp/
7cRaOiYtCySb1q042x958MvjmtSWP3vaSZNE5JfTdgF01nPTg4u9jR2yaPmMowUuRhtHN4oni+rh
qE7394DKYCkQN25/Ulngou08dmtPZFgyoubK3yRgyZLfkx//FXoCQ/sMuHqN41RmVzoDbpgVEd5o
lwVR46K/Ttb5Nyuj9CeFf3larDHJ4DlYx2zV4Pyaq2HIMqHNa0t+4K3BUtDQ3hiQ//K711W6tqja
iHMsc+cXNpNeZRMt4PGTsiUgFtHyGgF22Rpp8lMncCzrTM3ldQwFAyOtydjAYjzeguXPEeIS7kJr
BBjUSEWQcydw/MsA/kURXkLhiGMLOMI6GcoHcXGdM6Xkt8I4wKChzaMiaBkxvvtin9rcvlQOW2Ww
NHVh/eNEJfERGql6qp2hgq5vvD97jIYNZM4LQsIID6VaOLMdrg2FlBz+mDL/sArkQh+vXHiw01On
cCnzUbDscMhGuTJAU86pv44zG8qBbZ53yeuzXyWVO3VECXGxhho6fv8T7GAFmftxTbEi9Gs62rCw
OxqrFVFLEb+kQA0/2QdFmspJoUQrjrGzzC44l7pmy4xqqexau2Vs3jii705v/Z1R1brduNYu6uAG
qT4VFsf8GsQ0baqfVZd8znkdFi3qk4LqB6JCwtuozt3kvPIf2R+S5BjfezFMDg6SxX5mI+8JsPVS
pY9vVMcmqscAWe6TO62Zfx140cUSDtYW4u6rc6BbCoTbZ8hhs/O+RDcR4VqTiY5xoyo2po1BLFFT
/tJOlpWji8h6ooNsjPgWnXjrC2pCy9B9p4ZY5dKvQGmr+Q55SrcL9/Qsfr7DJbVWUJU99nMVVz4t
ZGGddVFAuKKZkcYNh6OXXlM8WydDUa0V3wodj3KtTRhLRzkGeNauoZ+XSmTzq0lI3sNhO2CNZVSi
ux2VT6eEM485zTk+HqXtvE7pZATHXeQygnuoOqetcN/mBmo60J2xIsezUU6R0VDxYU2BI7yx9Fvb
Bt5BfLgeIyf89LtcbhT8LHLq7lASVH1Nb0mjAbQH6MrV7xkxVHBCbU4ynSkkwPfvKDJeZe6eBKYn
MT2v36dml0HVfzt4MGrY5mB14Ow1yWAgv6bqx1eHh4Dt0REAOO92oesnz3BmB2/eft3hFps1b4vv
feu0UZfGlCroyR9UZmAlHUNBgkjDHAq1Ns8miGfXxNuP20cEPUGkW7OBCN9iJ8OGPYHFszUtQtge
awU3bQmPsB2/MUF0cdsO39fZDvB6PgQ+6j6UbgAHHyAqtXNVeNZS1ol4XdZ/sv8ycGwU5NDoK1Uw
M3ItLLnrqs/26k7IOqdjZg1MPFqKkrnOOdeOHjir+iAFpGH90saosnzVhd5/lYEmYOv1isvlknmw
+GYHldPapZHwxDDe7Nj4R7fg23ItL2w8bputQzWHrzEZ8/dMk/Te3Px1CoBnB6q3l3Gy+/jwz1+o
zck0b+PSnRkNMWTZBU1pwaT9cbzYm0SL0IdEux2URCqBy5LhF6q/Ki9cnCQWCgo36FJax2MeR6HG
A/gD1ffa52S3nUY/0v9GrQuNdRBToXDBO0rOGEMbwmLraOU7oz7nep5W6BOP1mbDMGVOqSoLbyKO
tleF7yMY+LJC0eCXM/zgOECEwbi0PjE/3wrbkdi4YwafwmHmb/4bQbQRRZlOkM+KY9TnFuRnW+t/
v0OMV7l+NrstuZGcNFN/CA94dVu444ee4XLtPA2Unq+EVpiq7qQ3Ncsfr1OW6fqZr6UM/ogYVCXP
SHQyI0H5lEmVDPJp4RAb5+lMxyY9aKW//phR5h4RIkBUxVm/KwKCLAm4H51E9O7CZmX0GezBomWu
m+rNV5HA9W3lqXDFG5V0iAVynCVz+X6lTxJI3MqGyHnKyJKWNne+Ea+g0XA2hTuKMXG9X9bUZ32D
UP0yTbS+e9IwuoFr6wNXAsdIv/0vV5UAZ9Bg1xfCsP5K1IecKGlXUaSvLXG5LKe/zdaEGzwi4Pwk
Ju0XAfwOrBBOC1fC338/VYasnQQaqdhZlupymL6uoLyr6fczKeNjrTVm0v6H6G/9KursCp70WYZf
ey8TtUhKHep7CrtEXmMciSdKV3v0CaoluFnXz2Tx71X6zISkG82qwmzCWlPhUzLQG9FjLOhRI4nM
peWAP7UmGD61P15jLcZUuVfQ/mvPkJ0L0RtY/e1Nb1gTlbaNpUhRWX9Ga4PrnZYlAJzfvLEbCPo6
yy0b4VolyyzLidJQIkrRH89q1f3cTY4P1rCIzLd+LuTMERP/1UF7LbeYiFGpbYZMpyU95fPv6K0S
654AK8OJP4HBai+vXLcVwn3xzQADHR14W0hO6+uPU2AWoQA6nAhtIy/AMVRyt7mNoiDKbIjETQYz
gyxeX2uVnyqRQJGLeEx+OLPBNZ1u1bOMbrvviaH5AURei69nKD3UN4yAuMLPfvzemwfODjOEMiXf
phelJam8rsqQTUWsDSnnuvAKZPRf4sQxFE2eEpLIjepKEDj/w68AyLPwJWIkXiIQ9Vwt9/RaXVRA
lUnlZkPwVzmuEB4nEC1A5T1XpB1lWaMg4S61/0vPwJbCyRNqp5DNwYokovC6YRLCj1pbrprYLwGh
ScXLKGouUDSe2Z9JigKGZM4GNeGS4SuiP4tIlXy09Yxon4PHr2BDaeDUvCJr66LPjda5CDYZYMUq
dEy/BKjHefGcQMSDwcobHDQeVNC8HBuWjydh8eitBulvFjdg+2MtsHye7sbRl6Sh+L6ZO0PiircT
vxruk55TA6Cga8aM786MjREw4C7SN5hAsBfwRGyEbpIcbenZ6rx1m3tdcgVqBUxbbwlg6glbtqlJ
whnpL32vPZISCuHJkZvd+pS78uPa60r7/rCRf+NSN2zwnldO8ZeR6b+0BXQsLnoK7THgkAGoXtS0
LGJ4RJwnVVLROGnke4N7znYLm2/NS5CoHBCwtGoKeTzsKje0aGHdRKjE+x1gllthoZnxS68EMB98
toBWN0QVVREmaSRqG08CPgesdYyBJVSJHUYxbNYZcxFXwGfNAwi+gjl1wyrfhu6+M9h7YJ/fXqwU
ZkW57lI4M0ctnhwavIe80zixQCqInFzpA7lCjX7Zk2s437C0JOfLVSs6GBBw0P0Y1/AEU7h/ITVd
4osJkxsM2TmFwbiAFkdiRsznJjthFa1Jeb5I62G1jYkOygCqYNMdpO5OVw0aG06+51EXwSBrRTrD
a4Og7NG4W8KFPyrvHpvzzV4A9/fRNcOG4q1KCVb8JvbG0MRCo30enm7lygSj+tbKQhV8+OJtjvOo
Z95XJn29IcIJBOqvXkRPbhx5OTVfG4h0iwEpAI0I6WwHuY0dpzCs1xjJgr6QR9R2BAUgvDwpc0aT
hSeN4oFXT0HLFrXi2FBEuSunyY7Ialm8UXLyvsesjlnhI1TXYZdIaQjQKegHz8uk+nr65JpG2S68
QMXGTf9I18CZFVgFoFBxzbUd6iShJ7+2FvrijUpR9KvuEq5nZuBHdF9K39N6FjrRy4qj1Z2at5ZY
UCCqlQNWg0/IlgLqKmC8ye6IzSOFFeHP7fYdGkRLpTrQQQXgKHJ53qrj+5hV7tmL8CP2Kzs1WzIF
AkY00mghekkHXxX7+ccw17TQYzfGU3FDyUopsvuS6JBWZ7MScS11gNMADkVvWv7HNUObcs/NaDe+
hsNr8TLuhclD9qMU9gSCtB/pUvQihqTptkuQz+RGODSB/2IMv4sDqFYtILdRCXd3T3sxdZ72GRU2
eeI9qVFKzWT8dFg2a8chYKfa9fF2/h6GY4PFpAEbPlV72JWRbNwd6SUOrzU/j1fhY9cI+xCKP9FF
pWjPqp1Oesc8JTca/pBxaiCxWg3nLKr2Mj2MPGThHq8ccloQ1mibNiqvuITT8xJuIdGElf0hDewq
umxgB1rMXgoL7IB2B7xRkIAbVp7faKWRDJQe8lGhYZzOQ0IdXODEvOPRgAC1SET5TrbxPakTfuxw
S09pSDGQ7E9ICp/leMkoSvsvHzQp/rgT7ZN32614WZ5KWlLqomvRTSI/7dszDc1IAjTmIN1llyEx
ymb4W/gmpjntCp1gui7Y2jMUAgNhSEklo/bI1oHiNqAv/kq1Ac422GJddnYJE4+ACZWMC/D/RDG1
hKF7mcvxvjA7x065z7i3YtBswOOVzmjV8BWC953KcLlPm48ogQqyI4W2kt4nxqq0YyYq6xKlZCe3
5gTgl7EMeXPnXJYB/U1rPvWrr9YrYtSHCknSJ9ojOUsp1Vxyad48TlqDte7CaLt56n3j7TWE8vSc
oTq85QMttj+XKED3z5b2nD6Og+eDWvMzNvq5utX+B8PX9kOeY/Zp9/P/GTsSZJ4inOUUDuOKDnIp
PaUFQEn5DPcb14omjeL4jP2sHnvuc17C9gOs2BQOBKeToj2PZuyzXT5BFCeF9lqyYdRn4DB7Slj2
Kp16pMRwFHbslxRj0i7t+gjnFlT3JwvMuT4v+wD5frUH8JOE3LOcOeDfG0WGh4rmUlljX20Jq8w2
dVx+QFBz7m2VsLKzu6ywxjnj1HhihOirlRrWpNHiB22MrwtHCxEAriFPpC+NvH7YDFRYX8Cfg5YI
mH9UyzU/o0IkP3XHv6mPeBe5FWrBBB3nFOBNtTEhzOwNK83UY69jzEKVAD6tEFksf1/chL9R96Al
pep33bk8kFpbOopeWKUeJnZqUU/SAe2ifa6ihM3Uywsjck8hhFw0A6fUAniLYBXL7j5+P00ZRli4
bS9YwlRkQYL46fxA06BzIRQz4GGdvArYoN3MMPuKc5yAcMd2LkOekHpqgfX4jZOGepER37/qAFuc
Be63c4jRim5cvLqCct63sRNWbjc1jqMculQdjQK2n/BbhEAX1ya9HUfVxIH027JlklQSD+wWOJqN
ltShtS16RppgDoCNXDq4ddd4zackzPNO3xFiP410zzCnCU8TKIYxsFDNE/7UV91rdvGNXB2dCecP
LSiKWd4KUh5oZRa1drfJIdtrqZhk+ggq/IIKT1ezkvegv9r8kKElck/lERJIDuCU+zjSSOiec/VP
Yy5LcCRsZDNW9nflwFeqTT+dCHKCdOR7WUGRUKyNgifiN2LApj8EqM/bWxHBYVcVIIKP6nFVA0WO
uey59f2hLudfQ1+DVcj1WBOFkkLYFRpCVRxyghqYH5nkWrTz6GIf+zZ+4sdgzQERWnYYe8YjThln
ssX/qBixvBo5CWaU8I1+Nuia50KflIb0uXDJlmqOm4+b9MDiB3Fkji0Tji9QVhovf7xYKqmgr9tG
RuF2fNv10JfEW08ZIh3FYp/GlytkRUHXKvCwC8jM0vB3ZzFtXlhMenDMif9t5+o6iT/ynm1DNsuk
hmRVUCrHoOY7Dax678T5ILraO4ByQZ4o0XHUeztVSSwWzqDw4bI+z/pSJbmgdUk983154kfoxDmw
aw6gPaCl4r1Ge6iXYJQ7DHHT2OZ0pJg/U1+XkPhnmqx3it1VJADAGcEABTDAAOg+Ja0JYWKnolPS
/YiwA/dt3VQIp44Dm0xOksKRRj5nxYmLzEiGOXiPwhJvlsvWhkrCrDpET3qRC4qKDU+WcYniIH7W
+ghq+K5R3pAxoE2QeNJI/o/sERXcufgiWnZS6CfeRwvDhuyItTJ/aRnavZo5MPx77QsPBXAS7a2a
FHYyWF+tSscjriN2+bldU4FT07xL6FEfzFbWWz2y9Wkf8RYzxJg74R/mhCcYpwiL8nkVRdiRLNX6
wn/NwA2w7eMUEMokV1ib82WsCBoBcz8HRLJQuV1/6Mr+JKh/EotdRFNA6w6S3E7LWV3wJIuAvnK9
+CXu22meUov0Zdu/F/IzKqHfOt2vbK0p2+5+Zsuse1zt8s4YalUGor1xdX7PMNdsUG0Ut5NytHAU
jrNHjH0rBO45Af8heXlLIc70PM0GC0OOrguqkCWiBfqTYKs52svF+2Izjc2t4f2OzlIUOrZltV4B
hiLxNBnsHNoY7OiatndvYJVzB1WSEKTq5/HfL40MmL3wwwMT4R4YztipnLCZcjarCkK4qGUvGPpa
94bn/ZkhqF07NgtxWATj5PCljBrvr7+mbpCp9GN+tO7Mwf71KmqTF2J5Y0k14tgdNqaB+sVzw3hi
8QgoWKxmn27I9h+8FksNYOfpMcj8HUGKBrAcwpq8Th8VIXHevNGwN4/cRQ77y752pzcuqi+bAEIh
AambBJ/BtK4rRPXW0KVD5lf+qPOcJlK7laI+VJOWfs35bgVKF//1o7erfqkNuX6/fQEz1ANNlM44
WTY4R/lkovnABwzJAE53C7iTqz+ktl+PVYxgsnzZgtkGcjsv0VnA61a5XN2tJNonX/J9IbtCuPoG
oUQEnqeL/ZxVnyLw/m4KdbeH3eeFZ5WKUSE3f2bX47TehZ8WXViRLYAmT2CEcwGNJNt3zuSJh4a/
Ue6EQORqogdXkRtbHcpQyivN3tFUZZPwNyzOQcs21Niq/nwd0rp7ZUFZ2OkuIz6Fm+EqULHcgoip
6NJ3596LhHJu8FVIF83YTT7JeNLx3j3lwnRZpipP43yzxOVOL2xaxun9/ha3bnTl+ojLDNKLLXqC
j99tTzU7gINN617eksKJelxtkx6weLhavUgoeis9jWi4Q3Q7gGQuFdxsFyviQ5vMUNtABzjzMw0+
PP1CIVQSnvawsxVywZWpBj3zdX4N2eiXQ+uThcbdPMn9X/6d73iCjxs3MQKoMfGWsve+V+9wSYKZ
USwOhpj6KRn7hPBoqWgwruQgugFAg4Bgei4Lypz+9yRdOxIGOkDbiEVeTzpO+jRBy0V9GqN/RY3b
u5WGy/8HqhwDw1/gAwDTz32rENKt+WLeC906ARhF+A3LD65qKFBEsVTsCEaW6jNqJo4ic/QeQGGi
Qvxf+NLoMiDpJpeaULfjt1TB3V+vU9+zwYHY8ut39Nd7NF3qDtxJrhpoXhuSQkMJWfD7319UDlPi
gDjFSSo+eaHRyhPC3XYOV9/BNRbg0rOISCNNPXV0jXV9bGj5oO542T5C/1OS9iDQptnaz9oK3Tk0
c89U39iscnI+5lFDaGmtA4GAIK0Ur3yR7k1SGpIQZzNuE0KIYng2IZPcfJLO/bkvXHDzAQtmXHvH
exidW1yM5NLbjW9s0mzWJgLanozADWBfQBQHT1B7iXQvTZE97n1AZ7bqr9OP6uYx71ndqN6okWNd
Umu6KnZ/tTOqG6ECHhS36ARkdVfF9+176wIw9ZF9512JGJafoJ2JOwECmnkRzVmrH/bvo91oN4hN
sv0atO0M7k20ZGXcnhorVrr7sYbhBk2gccwh+qTzYYjFFYHv1SP6vxYJI6TilAYO6NfshzJJFsJf
v6Sk3H+kN6Q/i8yC6/uY4OgM9TRenxrEDN9jl1P8yrSvA0pe+bO7AVBQrCfB9v8jIuTFlBZzxdgu
AgGupvMlLSJzciASZsg71TZHlsftoif+tscYY1PZ3O8oCwVnBhBcBwVLlCv/AO7PVRhgchCPXZ5b
GT1umAIHekET05OMBTzh1BP4lEKz7qMfSuwll8ekNMGY1lKlaftt7GzIhJ+pGN17Uvlf67I0FqvP
0mjaZCX11WS21pELHhgg6CVvzKhTGojsQws8CWzTzruWB/N85Ze0BwGNlMIdc3zLgxL7A6pZINMy
M5c3Y8BKipAnRVxBV3YWZfRvTuAGiFmH1HPXIcS+kTP1TBOGpGTHXWGnn8lgP5GB5lpG3QlGOoFI
jcCtBJqnCrKd2Zg1/JQE/jdnouZuAGu7uJn/uC/oMbQZI+K/JbMI5EjUWya88HGlcGdjBSJyO9gq
21+fhnQbiaVKP6M9m8E0bI2mo1KCa4C7YuwxWSfn9dXrvIGr39B5Ahb/El/TVNXSmGyeWTbD/4gI
VvoTaROyltlaSe7lDIDs4BT+P8362OtL8s9VJcUlv75GVpFyT8tSBxp+1/g25oXgORFZ1Hi2RUft
jCxglNBubamO5aHA7Pj1kazu9SxFviZJYzEBr8jsxie2DEv2Z2kat71drdBhNNlMnE/GBuFkxHYy
dwquWNgX9K9K+Ly3PJeePhQ6MBfILwzCuva32hGpB11fuLC+N6LMgwQR9xMPGssfpSDsJgQ5Ja37
+RB6nGyT1aQPhFBh+eOQVi3fsDJV8D8JeaxormLpUkMb4KQTRi0o0jBPFHO5IjCMj/Vep39lWFS9
9lfg6xMBFAJy1tpLA4ILyq6zSbRuyK+3A1EjFwb9aGF13SLPERZMmmnkWmZdzyn9qcBWopAxqP1s
id0RQaFrMRN+1c5qU3Xgf3w1QexBRGQJMCO+PEPLIgSPdXI3hQ5LU+rWFnJLES+tXrQTQsFKurB4
QhMrzTqrVwnXDvbx3OEheW2M3lOFi1sQcIULv8KNQOIVd4V0LJklLspbgGvJdk9kREK/eUdychny
FrV2paRjyKOOdfdmpdYtDk1wVqA+D01twgvv/eN7P+wrt4iKbvHHYqoPWUbx2pAjcF7ykIqFhkoX
mjczQ1QNMusu54J5/ZQDCTJey7XPb4KYiwjM8wYZQV90AnfExrfTPrBsAAoSf8KsspzAWLAJR6FB
ytavd55411VxT04UK7M0YcPWLotiWug3KLuvF9/EqvAjM9r6A+NZNwIA2dmgFyeDYcSsYe0Lo7zo
cr/x4kx/QByd4ViysePL/UY0CVqEUP2vZJp7l536z6opGvYjfNOVIstvcXchIQuv1zYH1MB++IJ8
fBkzty0xugQvPwTzhb8CeHjKlN9KHD/lZGcuVLCfvo52cEPhXi40twRIapI2fRIE0g5ZzzmAyeiY
nCKvBkOuZbVkjVjmK1BsPaQIvPP+7exrId2z8NBqkKNHvbxvP1EcG9ngKBmHkbS3LuaZvboZ7oFu
fc8jHSGTZv6jrKnn60HqlnZQZDCU04Ub55bZ5HOYW1Rcs8iE6IDEjG0Y0LUBcp8NaIt80Lvbktrd
9Wofq0TVMLP3nxnMKUz89oWwAZh/GYkbky1xflyEWPS/be1LrrRaAHyKcQ8LTPQjkxVB/Y+aIK/c
iafPXONBLzSmwveRR16hIeVH2X4/dxOAqfUCYbBEbL+qWge9Dxx65JAIUgUhtkzAGTjVKuMrv3CH
jTxcBid6fBF84aPSdDb4U6q9VMDpsMvV76/kOGRiLo5xi/B+oILujQ3x2tLdENYqhLmj7RNy2LCT
PvWaXZQLSM+ZVhxlqs70vQdtv3vtAeNMfG0vcN92ekZ354aL7DrliKIASPTa196gygZJKdAqEfVe
t1VCWANbLlODiP7MxGsYwcXXI6N/3cCdgHa0wHrIoHucfNGfyN8p9rmB6REiduYF6vlmcgrIcapd
WBiPA/NuyOfck5N8qZdI7aOixbbfEdHlbXlKORxckP6Q5V6j30L2EJjo4/LPlODLH/RirrvBLqBG
NANrqw+8lzc1/AaB6dymkQU2UyFlH8GMunK2Iietb1YqGbExDA9jfb5q3Fe/pCrQK8LsW+vxMKIh
ua8oZ8AZ2OqltwfQlKGtT5RSQJDRIWvfl57apJGneFftP8lqWOVKbmzS8IFcjV9hnPw+dGnjHWHb
h8DaUGHT1blH2oHIq5QxQPovVd4GWWC4XHaNLayONvBNPOQAAJRQYH7Xl5iIY6IenvScyKddBZz/
Gv3em3TSuviwK0mo/pwi1/9dlT7PZULIOfYWKF29wgE8jVVSafwWbG5JJXOz6AsqOfOuNqCs/XbG
OtjKlkMKGXsuL9CAx9X6CaZ4SdTdGEiUp1Ea4rRsVsfwrwoL8/WhjhPrwHxTqXZ9Ral9yexwAwm1
cQLY46ik+31giCMIeQhw+ySqMpQTyUgEzdxhnuLBHeqSBm4xpjcEuw33pTgrE3o5Z0sOXlQg4sSM
dimlSBpGgdUviG4HQ2X+qB/ZxD+kxo70o/dGBMgJj5ZhQNTcYBgcYk5lQsvPaHdnfoXoIYOUI4eZ
VnAwAeBNQv5w7xw69eCtGKgpf4sXmgRqfSjoafCdWjuFgyF1rBACMUGNuUyIVDjUvauh90RwyEdj
PX8Fi2GdeNNspScTDGSQrSaBIlJ5CAnm7wMIc/cqGkMG6LKAsiizuisFmiu1lzSe0KQqZo5upuCT
Y2XH11LAIdwrTcyAscN/VLK0vu+4s+s3MZlWcfJ4ISZBUXAeS6PX85+PrZe49LWW1OaWTv0zIw8v
qcu/BTKmYDTlgCj+pRyi2GPJz8blL/edYDE+3LAOnA7u2clCqU7f8wD+ZjsbQyfQn1qPBFLujv7G
hyIWdryDDrhiSK47G7TFwCjn+DeZ0vHftQXu0nokdNOw4f2m+v36A49rt92IK8cRZX5o4sfi5C+O
BF9a4F7PHCiXiAue/S1oKr+UVQjBACxLVsyC1YTMG15mKDNbvIrLs2rOJStBYnRMxqIrQd+2qKVX
Cploltp5b/wxbddsNaldFiXcrBnjm7IdIuLNlo9igRWGyyWYOUjqqCFxMQ3a4bH0vFR86XPyTbDa
Ii/YmyERbKVzfVMwU7/aMkp89qkFBAcifIoLG2s5RM64iIfkXCzqP7obpYZj64e3VcZwqyaDjJ81
0NsZkiCpFTGfrBTvtfEBhoaEjPYkv8HFtL7uevr1USwg+23NUPF3liWfpzKzlaPPHMhD67bkF+s6
8iNm7Gbz0fwWWB+VNFFkdiQ5YV19zfKm2j+DPaVEhXQF1SSIEZYL5dOcVCg2KShlFLyzjSXS+6Ty
vyTfzX7bxnBqLAl147kG59Zae37UmnsRDKFhCaaSlRm5w9oMPJNyzTMWUK0462DXLxHoaf88lXH3
SJSHG1SmZNpwFcVjpGYxl1iVRBQvxVEQNE7RMxotcr1qvfFHyj/saXZ/0Q+Eda0nCvK+NrwC5PAv
wTX3UyIihsO11FgF4qKz0AtdWKs9X7pwsU1x7BtJt9h5h8vBysQvWC4oaoVef617MlVXId4crNen
ZwC8C2IwJwQgxGyuROPLz/TMplHlHyIIogd/EnRbgt0saZq5xVbsw0RjCFsWJbfw82CZ/m76XkTB
/qBbTezAkrU+IsDujSXku+iGc2TLC+RT8LnU9SD9/YHRqt4J/mBB2Dby5S/Y0tx87ShlUB/2cm5c
BIGW0EkH+17fq7e+4ROYWl62A1tQhC+oGBPSkSIB21Yz06cy/LrdVTX6Lx/7z+52TjQrmfClBFiu
IJi6n0R6GPVjB9zG+PmrbrrYHfGDrXB/xGxO2zL4O0AO6boA2m07475Xq7pAY6Dh8QcAKHHMD8vO
86WML5TJCbnOO3Sr/ygNh5O9rZ0fxpaJbYaNp3DnSeA1DOZtNaznvyFoq01qc628wKSrCQRgRJla
N0lSgzaz1txJ10ZUPDzVRLLkwLsV1yoN75kS5MgyDSew7E/DVtgHkxM1PHEmEOptIhZxs8wcF9O+
pxYxUdjjC//OTfQFi+LjnARRVxBXgxunvXOVgicUDn9SViShawdsSUCB1gVJSvigFzgmACt6vgiS
SYbtsm+ovOYCflWVgAraNNIAE74xXavP6E9YUqoxjpJ5iAwC3P2sbCw+6Hkp/Ik8zrdePBs7ZDL/
26d7KIpugu4omRLBS5WHp3Q//9CqZUOC815Ae2i6/0/o4pHQ3yZuwa/7BiJyK5k9PbUs6gN2KrOi
bRtHpIhgu/NP01mm8PRo+zryGwNjGsN+JB+GGrTS0nOLWlXmgugCMtFzHq4aQcSnPwZVeJ3fRSWX
jyPqq+7YMi1gDq/gKHwkU/ZIKnbaLOhbnn6bSFEP96qaRQ/8G1QshK3ndXp/hNVXjws3KDTeTLlI
Gul1A6T+EyemiJ4pyuub1cN54u6tetFlErL8Us4LESV/S72M6jbPaZPaZWbC0M1fKsCkHAzMIxsU
DpDmr75lRFdxxGiFEwbZaW+Lzw1YzedDEkeGvq3zSDfQLi9Wjut7cX/Iq+BJlQG3HhxTK8SUO6qb
TXcKJLs2gJ8i9o+KKpXgCw3DQ58IWCL8F7dgwoAKXvkbmS9vwe+8/YrNDakOciNloyqkqBw49EAt
zA4R8wJ98EpfW+qrFGD2g1WJxEol/6rU3Xg8VuJ7ETcu5Z/pLj4EfN5ZIERf2/XAt7YkD7z5SRaG
Vjq+JK2GG/73p+vQ7aJ/Hx/I4ZRHm4Wf/HQ4wXtcxYLZJDI0G66ltwuT3y1VvxH3SJGi4KjRsKc+
sm45Cx3XACEuqshZMjQuEB2ajcGIzp/+FVP2Ia/fs78UbKtTztyWY3jmI2ZOrxSYINgByx1PxR9n
3wHhkZhabkSeDc8HXVngb/41oyE+h8MfJ+elv8GWu16BqJSoXe9BtAm2t74EQPRk8VjnmNmIYBRF
6WwUyzc0gs6/UOzcc5Qbcbo2SWsT3w1L80CEsF6IVwvFqTEhAC5xLDqhLml5bO9wVybskulbv+Rn
CxKxLbqZNTtG9CGkVrkXIwT5P9UZgdeV1zkBXSfbSuCWIsRo6GYpVhG9jMvL6dEfzNo8B84yCfB7
YRlHb8EMTiW1K8eT1xXFbpovTDAaTNnw64eHu+MLhIOXFMqpop3yR+WNh0dJsxcjTnuhpYHeU/3q
Sv3N7wKdbRT0TlS6gEUBJxoXCHmrhXuxMx90TT1eY0tMUTRSgW/fPqFwH4iSjOS2x9qDYp/Cz6Ai
qGF+eVYdXjs5JLYzsRSQyuR72ZH+EloNC1QnXtwBENoB5HFosdljpKxL4ReVzKvxIiXuAyrKBFu2
PbadXGa7/+Pw+4OaWSCzm4epYVhlD/IMiYOL/lJWq1+umZMM08mnttX6rJECMDs0pdAwl3xBXwF2
DuOqs5kGELT5RgmGc8bR2bk94bKKmROp6USptM1Mc417ig+9ttdT+Dk1Iov4622bHqLrCmARvJYT
T1dk1G2s95UyiYs7wurNyTPTq16NTIOuU0DziCqUCYj3IIxZhwsZ+QQ42zViS1YaSwoWW5udyJ7C
60sInF2r499C7hMKAFTpFbkoSNV8HlPEdzaigUHw04G3UDbyuslFKHkuAQRQU6+bn23DZTRg3GZ6
BgAIkwlGj9VTuvF16nnI9Otq/+a2UHhV0Pkq/fmwgc3wzl17D7BKUmw0w1UrqagaQsI614qF1Lsv
8DzAILjgkqHr4BW7XPAN4hg1ngqNG5uUhl+9IYZ9umRhLAmh1sIPngkKMJ6+/1uFMhjDHFs6Hk/2
eJ/xzINFxwAezYjdfmwtWa6Rj9woKZ3BHhV6qeF0YNwbMfNN8w+cTN6c4AHUgf6GhYPNELEnWR/x
i0z+R7nMWfqEOEeNw9KwuJzPCeP9SEnY+Qv0kqF1S2djCdksjDsgVGTcGwwgNh3gFtGEgNZPWEWz
PI+xxJob/Dt91RGbXalkcjD7hLvyqVjytfGFEr6zzmpPzGpQpUKHxI71gN+KePVCT641T5dqULXv
pibJR05EHpX/lzjH7NIQMmZBIfFySMbXYFLN3Wh9n0YuSgAfLVQzQdtc64HB1X3Gov2jsnosF6uw
VDuhntFVVAYdQE6N97HJiX6yXG0n3fmgMkcX4OenHX9MA/tUdG/sN2G26it9WSPfxlDDpAfDdSh3
nQ6RAmO7nb2JnbHvvm3xgs5HOLVx0cXS61VLD4a5cvR+ulBasgzWfy3HqUabRFjuvFjw3Jat8Owq
/NyCWItkymSSDHrpTd951MpBwF+E3jd4oKCswYZEQR9oYvt+Hs1e2vJSYcGBpuxhBgaw9SVdwIkr
tmZE6BiP5D4zfvfQYhhXLoAxaR7N/OXqpHX0FG5dqbhZmjJsVGAmBtjy9UvID1lAFhSYzbd8+TCa
a7/oXndJpp9LaOhwTIY1Cb+h1eq1JiEXpSbxjrjxk1pUGqcyjeLmLsGwiyaFlbyHhkBcC6I1iGEl
9k2fZ4BfnfA/PKdcrjEN+/NO5DYSXSgzPTRbx++EMfJthYDU+caWP6tBf9VgjsghQ36gQ27NMrXe
G6k0Ld1Nh7VFjK3TRvBioj/TOYh0GgeH3AOHX5BVoObAdmVoJV5MI+NDz9Yr5vqBrf4svhU0korO
4E8X+TFgxS+ifMpKeHqs63iVoxjSBG2XXlt0UfQskNhJcIGiQ9PIc8HcRGZjPHw8OtD6YwaxqXqJ
ryB0rW9r2+ux4NHjgGsFOF7VBTV3ySg2rEYgELIqhlRHEWGB89NvJyp/GIfTlWZhaGOm/SxsSZaO
WRbpPfKaPtpu4OukjkeTOHIozNCRmHQ8SsKf1sdd5U7z7CnF6XRgQduV4yqZjem1qCtmZ6hwkBpc
pqEpi8sDPTAZ1HXIeXiUo5BzGJpMakM4H+fiZxTnG7ucDs2Ew+dNv0yVHMw5GjuftlVCU5DL7W7K
64as4wIY6/BIaPnpYfy0g9F/9dwiQBXInAww2xrZLJNtvsa7XFvqyg07wZGzLoLvTA+C4za3Jh/c
Om4BhXTDoo0N0Tkf+7HIdHJkYeoDRQDBTv3ksr6BulXYZKl3VN40Ou6ref+ExGIOYRrjz5mZ1/KJ
Aw8rYAYehxhqAW84OsG7zMwllHZdBGkRTPlDDtuyXBHSAJmizsPlmz08072JVr56K94QeFTLoYX9
PVe8+k8k66h3hOXojI+BT9EujuvAfZ1k0d/Q8r0hrq9MbpX4V9Co5jx9LlHJzUqhDBKiAPSz41iQ
s7X3Y/Yvx0Wa90YMZyYU4iZWc0uk6sCk+kyFlFgyGTCNIua12MlVK2SXdevEA1ZgFbKHEkkHj8KH
O7Rb+C4myaQf2Q41VA8OkTLQIPa5IUVKa9B6/ZedISqnaAIV+WDSjCXvMoMxaUxjHYU6WL4WUlKv
Id6S7kes5ou8CrQOSGTLiefeB/ikLdHHT6LSBdKcl93F5rvU18Hwt57e720lDFsOGidAbTQy6WSt
JYEJ7JizGgTPVQLSvauSid82oXLfTAuWOnkpEajmScQhqWtvCbwJTY71pxZIIFwYz4vMnz8sVs3k
a35m+LxlWokDJLKR6yV73pTfuyOS8uRF0rBjYh1cUkv/aqoiyTaL05Q3bqaOCPwpNMzzoHSf7wVR
q7UGAK3yUnEeEl849QvEoDjEls9ljPDrw/FCnJ97RAJ2Fp+Amv0sXhDx+SFiLisW2Ks1VCe0KcgZ
4HIqAoJ8k4jUD1w6TbB3EQ78c/bGVvYM5tPEjKPeFCFJ/47imXqMCynDpN56bKhWtg1LDV5KFEHH
4PU7Fb6n+g4GRv20nS5fO3TApDhATRSkqV8kj/1tMir7GmTfbzC/KWvPspEQXE+WzuljujLtT88O
pLNw8zAi46e/ybikxwi7FEdP5zFl1qB2sghHJf55766KADhdv/r/0urIRFNmBwULrcFgi0boFwBl
oSv9kFsfgJW4cQK4tpSREY7zLaaZVGXu+OJJ55hOHhh71YmFlIT+881eNutIHUMXuUjQsHwBaSEU
QBgIxHOwQXI8GaZwIFDFmSYd97IAS9VzwTEk/CVXzhv8zDRKzuK2TJViWUaAxSZGed4/iWcNskGZ
GHaaAVXuTo1FH/hZLQLoNpRoGgza+vaJbpAJKtWn4ogdPbVcCNBSBGP9mCpx4+eYTrt+Y4F0cWJo
nNlHzNS3fiiYvadnPf8JPJU7n7UDi75mtV+gBdrsSDpPIA0Q713LIyFBw7yTfdEpVD5zxXBxoYjH
xpjTunY+Z01XQqhB0Z/czHXt7XQRonnMeojjUj9SQ7FsyPasb2k/sKgwSDd237NeZD0SMhsZ3xqS
xh5pdZ7lOxJpPyPHX0og5gjnKh9ZHUOthwKwG0z5zrUeqTgm9dCmJ6BDUilOOW/3YsNtmwS8ohAY
oJRNMadx3WjeGUJLVmU1mORSpMNgRNGzl2TF4bbrLJ3oTBHjvh/tm2dnoukeSp2CE8WyomDSoCSk
vX7KE7VC/ozNPh8z7gutMB4ZzfXkcMaOsaq59eG5xTQHexpnoKxaguy4V1MKjeZ4ARWDPbony4pF
AuIdRjf8ZyNRcVIxBAbVyJ32MsNChfZjLsgyQeRHYB/5Se7GmVZcWxRdx4WokVKA5YLQ+CPEJfzJ
Wq0fsxQbmSFjlDzHK7xhsKkYUvnC+tv9C4dz9MTlAeUD4J886Lf6Rq08WdIpJY6rME8SE1O6n2I4
4aciiZcfjSkKZg3R37TrsIm8ZE+/VyJy+PIZI8kem+bQBdgneKhTNrNYfrE16phnfczi2c2wNUnm
IvMPS3H1681Eg62kXzM1VjT4SMUaeMpemQSbW/WyUVO9U6+u0Rd/XcC2KNZNHjrQ43TtkbAGCTOm
EH8scSS/BfrBLWe1M37G5ibs+AJz8eYx1CMvTpnLk2qpKyqg7wMZpJ0br1GUJNidr0S3/KlW057F
rUGlItsGncMk7ur0f2khgBH9kgm8QSINaGOscmQTHM2CrWBmpvc9uj1u5iSi3mQ0rnFMSsxZdlYv
htnWk/2a8Gtc4+LnJS/EICk1npKCymMj5BPu4BNPin070fwQNGqAlNEUeUaqieC0g15dQAfwCXg5
MAT5ecM80ZRgqZskLQfIWhj4pyTTFDb9eY0CSxRRt7kx+aLp8WDC98IDAI087pxcxpX6d/WJ7gq9
tpZ+3dT0baQBjIHMtWwQFKRECVMKNmijdH0nZ8lWaboqPdwVOFVF+Y2G2k5bwYIfQLU6NBY97XNJ
2nbUXMsUtWxOy33rI891iXwqmRjifnYd5KJWOfofDYRUYBl2+HlI8Vbt7q8bipwgVwoSMCHexvcV
tPGl4hjk0d4jzUldpBa9IwC6LtnR6LZcjFMCdfr2kH+mnpFV+QOf8wnc4UWkt71ni4LhmJKuy/J4
Ib/Uwip9zlhf+8MGyicO9ynuJdSCsOMZ8T98fUAMYRZMzS5o+zggoty7pBeET1T5+oky2lAv9WNl
HqODK0qdOtSpZxf8uCkaXhMq/xlEZnY/TcN6QXfyfDLA+OzeqEdMNAlp4KD5iL1sKOLCKBWyC7tM
6mrx9ySUo8X02VLWXc6njpgb2k/xk8W2sykNDkaSeuALcZC2kAStn2ffkvxM79gEySTn46qQ2Nog
NeVS1ZKmow3lmg96oEzoQzcC6hW4vkvQu2iuCs3B42mkwkOIzSlHYSIQOEqClgYGXqNhqzcnoEyv
0XRaGe+psQdBxa+zV9KWADGZbqbe6f/pXUPVjmysekTAKNpUAegz1sC8cCbHE5xATganlsxHPnqK
lJqVAMnbXAnKRYfNS7Blu1yN9gcM0unn5fLjyZ6++AD49Hvd7f7Qk0UF18yl2jkZiwCSNhS+4BfQ
YnB0SfmIkw8VamL1+lNMW6JKkwHZ/0vHo4Qb99Q8kl5QKGJQ4m/ygcRpWd6niC+5GUFvnzyUejfL
39xIfBCmDuQbcda4H5DKBiLMJ6Zpr6/0azVQLJKCQ1TZ40R31isMy8p/LELw5z4iDWkSkJ7O/v0Z
R55po6Ncpt51xVnPW52v4VUEGdxPcP3hqRNfy0MruotLeE3YBDlfdcLyFx1bTYi2bhDzcEgJdPCl
+Fptn/+Sgh8C7Bv8MPpbHmEhyjudeXRo0QthC3HksnyQCoz38gJna+57HI2SCFZxkZR8B1ZJuvhj
rQOuBQGn1b71nbXpaB3817xISk0yR+PLNsfkvx2W6TvdPZZPkA1ZL9J9ltN1FpRgmvRSfso1vIt/
Y0mCASEijatqR55EmuqBlLAT+Rs0fmj1t7NLsM+QSLKb/kZqKXhMokwlnv3wS/4ERI9/FqbAQ3t/
1Ti2z8BCTtnvTEBPFhoF8/xqt/j+JGeOMQg+SBA7BL2X2TNOIan3LyVR8F6FxJVOBhb/nN2un3kU
TZEddnVz0gPa6fi6OZ9ucl/giNk5GXpRIN7PidzY7BFdaOUJ7EToMgX0uXeoYYK+OLuBddZZJq8N
ctW9/WqfqAKnCTjjfJAMcHorDX6lTp9lPvc4rFdHsxX/mRDjzDzwRogr5G7FSKqgp90G5UlPx3Sb
BoKupJKJFdBj/SZTUaFdQDpqA8SCWFJ7dHAmEkZi1A4T7k1VOYLRYIFsGwEzrDqEHglQihYipWm6
/DWZFioeR1FYdakPX1pd1hlFuDae6Jv9SWX3veeXXE9oZmvJ93EqDv05K+WgyjZa6dN+ASNxkHIT
kLSK4hGiyNoWJRNgt9iXezDor5H20gFmq3UrncwmRBp5O1ZD9wpjNiys7GPksiZ0VPCTXBmcOEl3
euRKEcWGJscQqTKoYGEbA14KCWoTYxBTiQ0use+iaeP3lWb0JhVsHjSb1AOjbr8Z8mCPOrEJrxtT
2SuMIlIGk1lJH9GdlNZwEiWXefdyuf97ZGT1fbvZNfX/EX87aamloaVo3uS4mIkHACMygTRLzTTi
HgxK81hjfiIXhlfh7PapRLLrSDWwRppDxil80aU914ptwU0KaErNGECkB/dFuDCcA832v/dVXpp/
cHEEJXJHGWA6sm+cSEaQrJ6gCCqXXgbPlMU/q6nYZABKzSjY1CJv07UHshyoJGfBrB9FINgrmQL2
zDW7RuDquOzUZK5ZYRvoEk1x4n0K1aR5MVe2rFA4LYsQc5GpkkdXoCNR6atCJ1lEm5DEFaO7TmSH
orSaMagAvKAJS/uyyjcM2n437shkcNSZdm5kI0d7GxLkXZWVpKuyeuzpPX+r613pKYkhtuhyoRr5
44yhQ9kD9T5U8GWn1D/+9UjA0qn313wSBfvx/FFEIyOtKk48wefS0j0kDKPvRubRV7E32f8VSyOJ
/S+sWhSbdgJYhmcbI9H4Oky3rna3ZHQx9TQONESbJPyVJLlFIoJM2/n9DC3TSAWK0aiJPlCpUjkW
lxTRA2BcamLeSLVTIbfkALjj9Vx7GinBjZ5s8LxYGdCZuZ4M1UPgBRtKivtLKWs3gEAHzNY3IHp1
thhOTeRdnhaKtsqNoqB+2TjYzo7PV9zvhDKel5YkHjan+EC1ZogTG1npr/qZmI3DiVwZeLmmf2Gf
FGBOEuDksJf0lGMewYfuguQDBbNClGqSTZpi5A9RDLxaOphKSEXFBdKFAatqqiBV6w+bAwHRvHgz
iK9HBnIDhXjOfLT0RkYkKvijdiqgyBhrCh9/50kbKzfc+iyjOGgKSRfIj3hQBi2MTBM3G2JKaiEt
u02WpkSrhg6y9GqXF2SwkNiJOjad7cYEIPKIn/g76W61rAFybF/GszoriA6HOH0QBhc3g5+UiM+J
rww7P/K5zN1B8kAhAvKmyDGZF4/SBUaLy5UX5Z23Ma5+NnxI8599oLGoiVANNUrMDU1DUsicTYpM
Ew0YV2bHyKa9hPFGoWKyr1pDhvWSitQbcTE4BgGoSZFfMEqlIChkrL1F0p+SZtiG9waWUMo/EGBL
4JFk+uXmnQUil5po4UNgMEiTEg5T41cT/9a0WQdAmSEDknMRiKYGy3lWcHU+2/saGYWWEFLbwFMQ
EKLeSM0TbeLoZ2jB/fMqwzTbhKg7d9AcI63yAYwDNGjI0yUiHLw5CrMYO5Iufrnhi0dEjvAtVb7d
yLdf6NtSIWuhCLyU4hDDEP90g3cF3wJQt1ZZvbfnJEcljdh96BNyFbYqm27mKkwxThU538C38fWt
Ik8s+XJ+WqAgb1omvGM9NlW2IXSMvlqqLvcB4A/hDIpQ/dffp8MBjBtT2yiOENqyJJq0D0P7Kp3g
5i4bwPApL/ITkq5M7DljeGtboe7ft1yyklRp67Fb/Q2zO7MCUzwqfYQeTJvrbJ/ucHDzWhWHgbDt
CmZm69Pl3D4TQtZGdPem9BdEkU3ak4mSg7zuz8Uope2tPDFKrC6Rq33ekqBg0cdfuPp4fL2fwY8x
4MWxAZx62SHwmPa9MRd8o3D21+gojMbbVFEMvh7AzXTaWPMDAcPQikXL224yZDXnm6dZMumj4xmn
S8TelsPsaq3SRKuiXjK3tw3oyX2So56fUaQVvzN3qXUt4T8p0RxSAggNbTIg5MdGRiDP5vWFsE3a
XNLUd01TSI7RYrIw8X7iU2HJSZH+voc+uUE+8zo3AjUzhbkNWWYpxVSNcSOy21uOKjMWDVp66U5B
UZTh9NDwZgUd3FrjviytvTCkJ03Ha/jnK2D3PUMV7MqDCP7mr/0rMqisJ+SoJfomjrkOgHZ1qeiU
YTM1NowwKq3GiCfK3bVlzIi14MdP2Aj+IS3V3lqKumPKZnuIevbG6ZNsG2+hi+r/t/N7iLj7onlh
MEJnyMSsP/3gIhcqhbPl/sPWz22milKCNCRNwnwD9xWNaDHX7vya+4wmAVqiusGcXr3bQ/4F/XRu
JiB1VMXTRFasRV83IkLeXyntlmPu7iQWSGxVWheAEEP3Uq2UWrG2L1Jg3N54Xc7zu0l4yv2aJjqp
LLnrCqvI1xFqoQBHJdCp74oj+cdkwcBJK5x1PwOMGccLbw57IIC9XMUzBD9T7tTEvFkb2SjpJWhN
JsAnjQZ9vBKz1DGaXNG8P11tmgfsRdCE2UNehC6lO8XCuZ6onVwuJndnh0m5rY0aP6QfuTxSOvf/
KY3CGJhSEmxaCYm3zqWWBr0awyqAkJ/ro7S9sOkt/O28WNdzDmFX4YpxIRgHvIoFZTPeUAthVEwy
783ZsZPGsVfIFEtvHcYTTwayMbNoJWON8HuXqzoPDfYlVV9TzuMV9Z6qiJMtA8b1iS68SUVri9qa
zcgKDdvzG98fvS0baJ5BKQ2+fGFo/dPPzSbBmAaONZF1ALhfXHk5j02MA6f/6Q6WIEdnNrmMppPK
qPH/2IN4uHP9S8H/tiOQBPlUWii5OZ5rsdUC9Aci6HMg/XvQmoY5b8R/+0WQsZSBS8vcKDIfI6h6
28olyD3JMF6SLdQQZ5XMdk3ds7NptWqF9tQwGbvnw1jsfAxQDZwQTJ28kdCRzCADbrnBn+xle/i8
L2lZ8G2OimKH1BrO4rlyN0smmeDMgNFdd9iZdCFJ9jh1W73H4Y2DwBcz/guQlSe3CrZoFAlXUTqp
RVvP0XKmbQgpsyH0U7nkrG18gLJLUlb2YQbCKwc/zw/vHegplNzAabx2IFdzTNMy+IfeMUEKlNX8
z4yfAOUmHEzmB/hFI3NC/yjKa/Vw23OyxUSjlrin9P4m2Jg/d4pV5D+d5mWcQHbXwSPUNfGBVsJI
EOSc2dy9lupYiaytoTPiNBBcU5yU7ICV7hIUZ2yRWT5Z6fcnHIzchP9bjySVDt0ex0Puto2/8TrB
48xEbkm/6rkWVsBiAXE2WCc2JkpCa/8GAtfc6BZYhEhYcS39x3OJc+ujQSeGU/bQTarFEJqQWFlg
DJ8OV6vmDMimUCn/Du7rWsiBXFiYPmI2brwWk+QlT5Nrx0jBZtrUisO7uRr6DHbs72JlzTB4Gahq
UNik8osGXNJPzQfr3PnPnNax0RixLDL85kIh8BWAZeGVVVwXcMhQoYd4aJCz67qLJjGh/DsBMKC6
Ef12YvD0udasgRyBzhzWXVr7551q5ijLISkIyoAKLs6yDD/bVfY7qQoCdde5BlL2d69c/aUC5kon
LbPiBlPbdlk5p2xClAMb+wU5oiMc3mAh0ekyWRgoEA8XOWsUE5oPMYfEAFiAK43atbteuPUTkGfY
9UhTeBuEaoYSYA7EZ2moaCokb7XZnXLeWY62rJ2A71aJWXuHrKjJ/Hz3xp6qyGg4nEneU5vLoZKs
a/gfeLK/yKpQfj7ID804aKods0v+eyGCAt83b6o+9n7b4zOlpaDsGpe0p8KEAEjOJ93pCLTb4iI7
bANFNGrF4Sl6m0IYzVkdSykQs3VLw9Q06tlYtnEANkNW2HT7MC+SLrt6J9s19c5RZQxYCCH8vtaR
/JNexbEXnUdHW6b0IPRm02gSd6iKLmF2UxQmHMfKZftVhe22gkcPuWy6xeaMacb2lRqEr5H5uOed
RcAf24UaBkSs4QQOoSRTNoKEeTPmQebfItMZIFESVTOSOdQeV+eAIpK2xh8SDSXjb1Ukb9Qbmx13
5sKmsGJAl5mlTmCShOYg8IdpDk5X5mDDo+q3S3CkQqCR6pDF2SmfHS0eSe3B4k6jIcqJwBkL8dk8
bd96t7tZu4eNuRoJcn7ft5TOt+Aij5RLLx27oewFkdY9ghBxub7WjInmd8+WwGdyOqxtqtE2Ud35
A16YAVo63jYUnF+5rlfKzkV5iXfvlTtmrot+1JnyCjb6qcR2zwKkrQRnnt2e91wxHkcGIrWDzxcH
xsBCPpASoUEC/96V4FvtKws55QA56ceSv3nGxdG9vln68kzSyeR57Cjq5My5VZXyrX+xmGTSdPKo
mxQ8dSmImTRZ8izkCrLJnOttGTVrzbjPAaL6OA/OmsuE/HZsXY7z6mZ/joJLIuKQ556v9gt8eaJV
Nh9BrnHly4+rRxWQ5c+lVrKReMaolk0tJdLWXl6pfMnmcCZr8HtAGfrt5hvbWOO6RhUlNJBGjYkA
Zgp0uDZbRlRUE93l8dwnO2dMmd7anlvrQ5OG0hYLT9qcLr3NUoPwIMbUvO60vtTmOD8lywegcEW7
rzeJsJ6mvyUp0ivP7DkUI5nZAjQC3VbbNiy2Pwj2xnwWRTWT87BFXvndb3KKER28wcPaePT4mX+i
LYdZcHZxKNrTzILRcvoJDNWULuAnDAaVFUPGA9EvCwWW2movf9ZerSm3ZlC2/hKh1S7s4VRkgWKz
Jo/2q15Uf0pPI0+I/9rBJQcsS0kkR5VVNhRSRghA8TTyMoV2ZMNjkUOROi4/lgUoi1akd+7WVqgs
OT0ZYy6APpgoD588eK0shutM8hs7abgfChpyxGCW2bVJjEUfy+9v+E3T208HAn0zCJcdFK2jTcDs
g4dDDU0nj5eGzCH06KHoUWx6XDEmdtWgSpviF6t4mKV0nCJ5HscIBlvnTq0zTpuDbnMatFHgAh20
BZsh70iX1ssenq2zuL9/T9F2Qqo0PnclL+ZXMOJPPP2HkIdgg4OMtgXCRbM5oX3n707YTPIX1SCG
GPgLz8x6QpSIig8Qy00NfNYt8gvwQysx0vQLQ4SnK38dhEVejvXLkv5B/suuxtwCneSau7nu7ATw
l/QwnKp25z5sDw/6qpRV089tdHv8+p3/N5Aa8hXnV8a1R5CiuWFePqb9WlHUStfjkYrWyrEl2m7q
1YU7eAmeKRA+A26szbwUEz1j39m1p+zOuNKKU55fpIwNsZOROwutMyIeovv+ATnuZU6FCjpCklXl
0Ype8oXPcezMAZH2iipy0vmmOrT5r4Xhs3/SMLemQtzdi2iAbrM5AyOmI7uPMmrI3TBkOYydl4p4
kt7xS9xFUL/k339nOFFG8ovJ1w4WMulFffkdXeZDC5hNC60l2a0PUnrXTN2kw8JX3YiJYJYE/lg1
fyU6zByHE5qp6sv0FDWF62NmpCSckaan1ISDxLBlYwAbYdDNorkuci9OJfTkxWf5zlm5qPmABMdN
KNuipe3z46yu1uxsc5QI22NG4ahmLAg3sIjvvyJpj0Od7XvklyHUXyWXd8h59ah7ihTkyG1tCyOZ
HkjjjzXrVmtYg/Dwq7zOf8h32PXpKFL/7UsjahnBwJUEq43heKzlcorgltR+QczC0+C3Ov3fzid2
A4PmMeBpAgLdTejGMMLyd4bFM9biHbfI+0ZZMqhVtPtlDpZ5Ha32bxa4G/p/SGBr+yhDIJZ4BYdG
srvY+9KgTChl82EUrcKO8s11bQIgzuQAwwuptC/R6+FttHFjWsQKMtDzJTzzTxxtjaZQW06mL9I6
rzso06BjftCwautV7obKty7vHn//JSgGa9f3I5EHxY8Zpo38jR/j2cBX1nF+Pw3A3Yo/cPCdeENx
XPihylFm4W/OC/ze3D4VOy86vhEl0lcOyq/KKBQjTz00lqRWRSIVwZkE4MKXvzLgD60/wQTzmMeR
UprteThBSHsqQXYuNw02QMUjGWNGPHHULjZbXU0bytYMtja82A0If/8TO1TQbI4c47qgUxysDuHB
qhSd89uSCnjz2Fc1HoZw9IyI9EGg3KUHbEgM+0SLd4apE7zU2lELHOj0d0l5v5AjolyFbA/HRPcY
RQhbZJuAtp8EDMi5BPJqrvOLzF4jNIkbyg42mTBLdWzLhc1DIFSq9cp8cdkWbr6r6q66fBvl/AS1
RZ9m3Me8EwiNS3vd4KRLNCshceUnMTpBaDqfJLFyrO/4ZZvQHhuSMIbrWTmylpzuPDLoZiBhLMWA
XzqMwHtlqbNKb5sOhMJONS3Wjth0yVx7sgAwC37Zm0bfXN0kDdIrfOcgvfFPxEQOK/Esryjwtthh
5A0JPkD/6ZYYH8v9Ur74riKM7AabaXy2WHQGPFh7yOcdHsWNmGNAmSvz6MKD/gdUT43xfPks6oCn
xpJeKKGEq2JvBGNvfDJbJO52NsDEjpxhk8QWsRs/9pi2netd4x6dDARaDuuBWBFibflbX0xZF/zw
kU1QBYh67pRBXlCQ2maf3w8A7ooYvZ12TCXIb+IiGDGCKKwgDO3LVMmQ1yFziDzZbUYwXO94MSss
IFqbuRKy6D3NUDRBDuAN5WaU6Ne6UtpMAteCh8pFjLCysjTpgsiuzNgUV6suID12iUA4kU/g2f+M
Y7A9YsHBzxA0/tw2CXskhTpceWu2ItJ47ehvxdqOId/seAUjqSxUbWypc5tkmkWQ00Aoew2+RBhA
QcVqt2Co4Bi1kqZP227WLmG7bGol4SlVuZIK3waiE6iGiSF/JtZlrE5qLnbFHumt9QpepR31G2z8
cZxax2Ii2iI0vppD+h8yg4ikZ1sY8D3geKIVhtTFtt5vMBBW4xzLaodHrhDW3Z895TzbfKAw/aZt
40xsyNxHQNFvAgRVgotdNHTB5N1y/bzJE7tQNtIE+Qc+I+tQQ4IHKH9IgM+W+VDedFH+IPrfMIws
RFWdDaADpyqL9IAiHqZBf8ixa28J8EQ4fEuUsRNejPpR421e34R4AKsfMKp2PResiLinwl7/PLMQ
WXRUYv2qrBUan+Uo9zFOi/ahFHgGAPc5ctHKtC59nzGEPD77ffsOdn3rJRmGujdAwX/D1BBK0uiU
/mXwZNiM5g87cpnHcX+q/R62PeOCqgzsRRW7tAa/Kn4G65rOCd3F5KCVisEZ223BdJZYQSQmysHf
KOUSRBquQzliBLEETYUl1IWEYTYU/hrzRGWtwc7S9Xp/MxCFNC2VVDfwPVVmf3uAFcgAbdK6drZB
5YmdFF1WzXLtPrudhHkIyiwGm874DO8EvSuzaBTI8KFXUrJUH0SbvsQclkZk69T+jeN5Ldi4ZsKL
44B+0yZ7yFnGcTukNXu/DaRmHdhxh56t+m4Js2ewTzigm34uzzNi3ODX9dddVQsN0ELdK+niFCct
xvef60suH6yfXLvAAV+/jdMlN6MH6b7UejsPg3Rb/6SzS3Tnlga37iiBOCSZZQ7feLaGW04X6K+1
gltkQShXiA4C4pZ/twhFeCUYPHPb5yKGLaQRuHspJkeXsaOl8CpsuYxNuOlldPSdgHMhaKLurXGA
iakotlxtjvPhIsnay5AnGxnXRQEz3/shDgWm26AdU40UetTUn75qkPcirgtek/TF+A5JfLEbvjZr
OGXTEvb8nlHHaY9PGEfHBHFkFP8mHEhkEqmRfV8lRGlTesWW+JHc/zfWniBmW7nBpVbBaXkRh8/b
6sy5j9kusEa1JULXicnSoT8y3NOjypOPfcctTmOt6v8u8r4zH1LeuJPG/4BPY4KQwguvdqRl25N8
aHGJ+H5uepkKYV7nVoKF0u4rRRIbQADOaptc6C+7G6GfA9faR8+5VDw5PHx2NPgIvYxY4zjN8X42
FWToliHguJ5J33cyOa2IrXkC/S6poPTh16H20xFyZBbp0OyCM5I5eD+wqE9HpEsWkSobY97JZHIx
7/GJ2jb7qOGNZFJGI+iM8jcBCHXfPuqUkalCH4vzHjn1xPFBJmUfHeoMuhV1PeWLB+IX3JltD630
JlF5oCXACMTX1ml/AebXAizgC1u9bsyu1OM0jWNvsrZhxt7+6ncdsyMs5Uzfz56iC37wojgz1bPh
8Yd2g1jVnR/2KWgjJocOQBkftGPKCqVj0VGZiIKGhaNiExmgZBfrIHq09Gu9WgEJrSU9w9ze+k0r
oPLor5k7LEzxoRhT+k4LmqG+xUO5yE8beAPOmpzHz32imAJoF0ln67SC4AKYYdLUFUGma6JQcunu
1RDKQho0vkNI7riNz4BJ3+ZWiVe811+RO8GzDs0odjw7M0aqP9C888qBERM8piE4IwpozylCPBBu
eJosrK5ldQs7FGjZWyuF8oIVKews7RmL/WknLCZ74TYTiyZczAYApL2QwBuG1ejivdedO2s7Rhut
cWNklLuWii4ckDXNyPILwhoezUtcOmRPBPboc8PlYrgFpYFVG1dayQsZ60o0mNpct+0OXWrkWCcz
NfUvcq3K91k5DHgqrTZyy1nWnNr1bMZvuYkyLVOi0LJVBmzBtNkltJLEiWi6l0tkTuxhWOqakbvi
nQk5KgP34KQShiR28LHOOjS16pyGZA+Jk6Knie2XSHxi7BqR0E9UeJ43+O3R+WtKh7RZhpSgZuO2
PrsMOBVM3TmShtdLkFQbvBMbxkoIg2LBZCewdaVGaPDlrhn1DiRmSANWRcVUBzCT03AEOdy53sjj
azP23gaAtSqdPWYz7gvGVmBzb0k/wkaDxyJ+WtEM8K6pqOtQTP0p4JbaRVop94JFZrUj1B+FlyhD
pVIescQmMZSHAufy4aWCX2Hdjx2McMSusxgEfgRxo9zyhF/IAssInEvykXi1B29gzrpzYVcf/rI5
k454zGLFP1cWnguPMNpOemirWiLFi4JaPt2NeCfxORl7rYaKxAGYCFlMftRQnKn6v+jcSBV9xl3/
Be5Z7HYDGgOgVDnrnSX4Uf2KYz815qSjlZGVnmJ3J7qv7O0XmVa9HbvrtY04adtYGF28nAIpjOt0
bdE5xH118cVk3PM5pfI4uQUDJJAKZye5IFKRa1ElD8Ali/7HnVN/0pQNfOPK10TfwBNeddV+mSMT
clPiC7IBIJ+Zi/vlrkCdeDNgQXhmfp15zMiQySomggnhmhdlJA/1T+QHkg8x/IzaReF0kRWxA1h1
LP1PBKsxTcVZ/ycDgDhHNStmV09i8tjmeAoq7riV+CC5VL0jiH7yzxVxw3WgQaFt2toPkuDsIO+M
T0ttcO/4uIonlxJiKUz7hanyJPEbKxnAwIo7PSIy47LJ+GlZSK8htx9Sug0YQpzeP62tMRstMYn6
/txEWIa1V/lwOlPaGowZY4jRR0ozCDPSETfIByoBKGFW0qJ5V4ySOpL6hlLdvfTUQWbGZ/VJz+IH
iL7183xIrJ9DY1wCoP921dQgt+WHriQsI66k9Hnkt8uUwXtrGdMPTEwLgPaegNmpmgY6ag+rAz6d
GEhMBtxb9rmGXY/zer2H4u7jmKT26PPdGJF0w1CYt2iMMUkc5xZYqfe+sRiQ+sukqHX+eY8flkIs
hC9QDAsab0puEWBGvtdBOKoixl88mfRv/LOZtv3Jh5VYHYFwjQ7kSarq2drw/ym5tVaW1o9VgxCk
pqVUz4qZygIyTKzq2BtkccDC1UyP2rpEBmCwkyu+fsdVAC8xYqFJNL0iyPGEwfP1wvvhGIKydhjw
N/pjKAZxtZfseZNFVmW0CueG15m8XTk7ZQRq22Xxwa5itJpjXzycNUWUJ8gBWGVxZCs6vyqJ6prq
u3K2ule3l73LnfUj61CCbXWiuZFiG7kXmii6U7/4QsyoyvmYkWWukl180sEHvsnhwWneXM5Q3RHC
lTMNgFOoUbRvNwiDvHjSjujkMjAqBRp/e3Csy+fOvxKixEtMYnZIMFKWBxT2PMfTzMOmKqE5T8/F
k7YKZMvrEJzuyWpUBGfrqfrtGBZPMAHHRM+0bg7P1DK1z3QnJPK2XbN2t3t791QH02wZW/zdnAIQ
QsJpqFcyrit2rwcLUUzQG+MZIXgo5hL1XeMed2FeHNqiRzyh1hkpNVc/X1PuErjRHgr7vkWp4Hwd
rSL2xkSTA/oX6+h3F3jKYQ2Z8BOsB+SpqTLX24T/Grpwrxzg+OJMLJMocCGWcAlvxnbzT/Fh6qLw
pXBizulQFvABSIbbt/zuNNd+BPTKm0V6KVKbT/Dq2acFRrPGnbKTWBW4KHIOGbBzK7X2YMeGI9J2
d/uY6q0kS/UQLDGu7mILpbMW8eu/zRkNQfeecooi4VBXxTFbCvSq6/Y5mG2AzSjmT4p3uhUzpHW9
z9DHa+j+McA4XLPommF3atJxaS+dUHlXhha9C7S5v2BkMCy87h+KEHLPkZN1FHtgUfQkZqHt6vIy
EymHbw9IdK3RpUHT+2ax+2capsvMk99A8qFfuyYrYjfhz1n2gTtQnr0JNI5w0EhR01FLLlFY8Tgd
ToBFjQm2XuL3BpmQVL7m5ktvGZTgSJCmzUvmnQpZs/NY0qaFRrVLc7/G+HWE0r1GeEsDwb1/c+6m
H1rJVKgi/Fae6zu/P+rKte/ZhZrX9x3ylgbaDBeMpzaEkLObhCxq6bnMUCkkCR783K3ICoZTVUeW
0MIucInku17JqdQTZFP2jMab/eVmXF3Yax5+TjM808IfZRRFfxYMptwVvPmRL+f5tjhVYnuw/yOE
ZfRpHfdMM4U7kdqpheFqQ7RcKgNdtilnkdtuiJ+MIxZvro7w6cWMgg1th3UfSpNfbPtj2YuJViHM
+xZRzdGMZVqLOzsCNwL5PH5dUiH66CtRf4MLw73NIsjB71H3IFgiemu7tOi27vyKtQ7LHsmvPn47
3CKsVA5gIoRVOfVwunqFbIDUEQhR+ahDjxn+Cq3Yvpdpj6SC06aEn4SxAl62QxTvIwU2s9JBYBXw
wC3ub7CKOSqJJacuUDeVs++A6OTbdGFGEzQ2SCHP2+86dXoXDOaOcJiNi33UG7DMFXmZlXvfRIcY
o9h4ZMPc08axe4GcIB+FkuFMgr//AN2UhtD1Xje/QsU7vmZZercxIF3ol8S6aPe2ALHqAuJwwtjd
+1kAJ8XQ3QkQCenJw5k0rpfHwo7LtvLIxylLdm0fu47grjalHpzCEqBJE07VPqv5LkRtVAcJqbUk
IOsLAlBasXuKIGCR6Vj/FX4jcmKS3qV/LR1s4GeZMyPtQeCP3kmCCctbaQxzSKyb/J5boNlsMZD5
t2LNQwtc3H9qz0S0ofr9T81x+PJteellyojq1pfrTe9CrQ246aEZ6zmJoqV19sjuUGgCrxW1DIeh
w8as9JK5+T6Dmoq59hRIbCcO68t5A32Fu3ziOiztUDNZcP67uYDQvPcVGCizLL4jfHujh9EqHJft
bbkRkovW+lUMb8vnAwqq20AKE4fqwScO8yvxA/cfFb/yZgkjH3XTQc2qvnKoN+JPw0UVqfS8Bhpk
i0Ef+XNDmsvCCy9msRFeLS0YPGjkXI5UzMcOdmAwp9LPBBf9TbrJjDpxMAUk+Rky22yp+vRsgMre
lnIA12uqAvHV3LpN5xoX/3pq9nwUFnJhw42tKJJ1Lu5E1EFh1OqTGq8fNLy/Pb/prU5XYIDSEdy2
eLvHZRxA/TNC16AFOM+fmF7L2kZt7wUlJ5D5ItLtd+l479BK2VyKlJDP1Zf2THXTSFeu/cnjoiSZ
1lD2KcsMGHX4WizfAVBrYadIfSBfm4eb0aqaW/uKLL4/Mh9sWaeMrIek2EQcMODyLpWGd4RPu93/
Lz4aYidRPXlGZ6kKCLs+ibqmqmG694kQ5cYTUhTB6sC9ddpUkzDsIGWz8wn3UQ+xwB1Bu3bLfJJY
NITAtFgM1UdpCZc97jZpb5nuWAgHruAFaC9HYbsct34HhGVDrOtlxsqf9ZU6ztz0BRPK+QUFqkEF
6cMIHp53PDPzRmut4DBN54sizvkLoIe6GHJz3NCQtDRLbEqNODu2kBTdRyiWiFDjrbU8LX6/xgZS
8qBDsrMaPWzSepXUX1nkqAamw4y8jLZZjngkA+hye63v5aPxIGYhfkLhh3GFLXSwNkrIjbygmq/o
F2djJyqX2txzplKdkcwSzDwvd1FMNtVdbHGH2U4CyyQsL32qpgzzXWY2pHN0ETXE2p5zFhWnPWR2
cvp9Row0QAb37f0m6bbM347IoVlSXjxNWzJkewcsG+L8rCvQN653+iIUuFkem1ilctEcQyYvoH6h
tQxwyuu2R4GEVey3tVNOExIfYWzvfMHDFVQI5Xw0/KepYyVmtNgvk6JTaYB2zML36cJDOf6iYZdX
S1ikOwSyVDw8J6R5vk03UrGHQU5fxHXM8QGyRs4KzIOp0le1ZOjBPUGVxfv3PL4u2BoFY0p5dmrc
JhZgp7f5ah5su6qS/Gktmkxy1mJrgaBs5nSAdodLrj64SbJY3CPP19PsAGGeHOmQHAtEdmJ4Czcb
pV0PZt8b/XPsGy8u+qsmnpd3jWC+MhOtR18lX+mAc//yeam2ODniYjZd6WCTpB1iUYMIv3GbZ0VJ
sVkmk21TC5LsEO1nuRGsQLM+o8r4M0vgvytx7OIXzLelh8FqpjdZiC4NXj7XCYmPalbidRcQB8hs
B7lYG2jDcjUu17Jj8UwdLOSQ2PMI1rYhOG2VYoeQziAn7t7Oo49O9wO/CBwGg7y2lCVIWdhbu/aa
a41orVNFbIePnsCdgMprT29Izgr4ivJOLL8jvuAtsv7ZfOBrEkfUg1jdLJgkoVEWzECeuxuBp4tk
2ucRqWKwRwABhh9pxuNO5/cpoa2H3fB5/3F89Poen8gXkEUu1xW8sSDtcQZRFPzAzEEGKzVEGAtj
B2QSGQK+5XWjV4ouvUK+a+tu8bYjt1OsuOXboLTH9bQ5ydJ5hUaYZdqUiOUuZs5jmoRL/yG7bCVY
CIPaF/4C9eNRrlwhTog/6PdKmX7n/PyINV9KrARE1gnvhNBi3V82NX395j3qEAJHxKJEC8DBoZLw
1FI5G0RhLZb0FqS4iWhv/pa6B370QYeq7r7WtR7PZBk7K66iKJF58n4PpchvuleAtUlbrXx0L9nw
Phd1f582H7Xtwv/7WNvgaoveO1VMAHi9cmAg5fJKbBYT6Iz9s4kTUBFBZClX0yaPqTK3BZf0K1Gz
TDjtCRgrPCEtaPij4Nxkqtg5tkEAeYR6GdsmXvYgPnKCAVtNR+TzUscvuN2vKjO6MeoUKf2uMrlh
3Amk//rnpmgZgnD+dHvaKuwN607Q1ne8NspVg44W5dN7OlypzTEHH4kDjkgrEjVLwIhYfXVRoHai
KWgaQc+Bua6rESVorHHiIAYKkPCze6mGMnzzvzrJvSlUGdUsgnuLwKV2y7ZfwnLKe8NAzVv+p2od
u3f2+vpKbn3jArPXc1HtwMcl+wDTYeAeJPuhgsz2LFWgPnxgU9wYRCO8wr5Fqhh1UX/awPsnR8rQ
8vowiC6jpc9ZHe14oRCurBfm7X+9cu+Z9yAAJgN4ysHiuqpbJO1CL/KnSGLe6mFl4wfb+ehMOzOu
u789+RKhyhSqAUdkC85bKx9uQgtqj0AWr4hKOkbyeC0+rPB8UKDBOFedcq3rmP/0suQr7mBVXFIz
BYTL4dyAAA3VvT2j1E0kBfJA2UkPy8rlWYPGriKD1WY+YONbozuzI/IZj72tGYWMueawradrnduC
K3vY9SedNhhQZL9cueNOAJo7A/o7tdjtojDRenCgbGhsp38Kzaof1e6kiJfzQiPfbWrqAx/D303N
wuCSPtqxjAXPUwYICcUUxCxk1ISO3wpkjmAs/SAdoQNoJVWUX3XdOtgLt9WeYptR0DIWbIviyFMe
I/ZFbujLgVXhgM6NH6tLD+0OZyJwEMb+SvHfnVN+jcPu+MBurLI0SZZqol/3EHWrKVuZucJqPoHg
3Tn+5rJteeRQwdm1CDVmUMoy66htL9KXm8J/QOF0ZRq0qITIpeDmuyNF4fCoYhuM7p5tXElNZKGH
KV+JRRXCoeAbGgaIIUFtm2FFvjD8/IDWQ3nIbzoVhMjudK+bjU9CKu2mG/UiPDUesfIr/3como51
W13OYZF3xpeiCXQpJI2Xb76JCN5JTUZ4O3O3uYW5WpW2dkSHukBanKYsC0WD9OGkVgHpXXyZGEWD
EZd0T7HOn6DeNibJAvvEVtWEk/oH4bzeIQGfHOKYCweubl8SHXNqMn8ODlt+IxiJQ7zNlfG9QYUv
oasDevx8Vgd7Q+iKRO73MKmOF1WPzCpq3l3YBwIgGYYDlb3xpUqZYhw+KxfPaEBMvgG2vmqTj18c
6d7HTsvWD9bYouQanN/x8VY3moztT8PwAn4coAQ3nkSLEy6zr3fMycHLkaJMCNGDFklb8iNY2g1a
Yl+SfKxNzWe0IgIw03Dc0eA9DiP/whqGzLKuBVjVvRMjsoKXcy3pE+cKiKObc39+OVxQM6NOX7Dx
/w/rnY7gw/rTFuP7R5XtNI89IxRaMUi0fJYpCn4CEG8glc99/5JBE0b/zgJKnopivVX/uw8vms1Q
mAmf3V3vicZIXksK5ZHO/iYsRmxdXqUDu0dGZMoaLYj5kh9fYQHi70rrg/HEpZR6GB0ypVvPjt7s
3Ewbvw817gBp8ojvnNUXt5x3vDpBr9Sp1HWdMNu5fcPAkjF5H0I9b7AhcN1y8ES9Fpyjpk/iYrY+
83SuyLMic618fwyyvGnhKCzIzmIIeWJIS0J1dE/vtxPFLcDhXbpOdJnkarT006rlbCnBdRRhIAQ5
8U39+24TSy314/tyRxgqkDtFJV6MgtxXWX3bacrgeJBTVPVR6PH1txccjEtG5gcAacx/p0F++uqn
zljMODhZBwGGBANr9opmd9hSstDppNq4wO6UDYEGkIQ/yzly48dBP0h1oIz8uAjbUwSurrhkiOWu
9Wd2ceNQ5nASntHdx/aRLNkEHqTm+3QpfLTE5twipsbeCgo2lRq/mpOFqNJueqcmjvXwAn2QxJ+O
1suY2y9Q+3Zr8TWMyUzEb/61dt3Uw2UCokJlxuCsnhkkMg8r6iijTz3bMV5w5DioUHnC35iHOmqO
izlyoVZbLut4QaUTfxeuApVss/6V/pLFiB35ucyLG3vrTiuu9bynM82soBd+diwA8N+ckTcxDdwC
hIfaFubJl0uXVaKkhts6ooM4V/uVvyquow1kjEdHFGGeYTDMLkjznfhQZDqMofV6ZS1m883GxWtN
FWOhyLOgTk50T6uNFQNvUpOk6zhAUyVxvlymiDQx+x5iKbbelBW796Y+wbeFTfkLAgkWAdCjKTQd
sbrbwGg7KTP+ua7FfeyLPedTrP1VhWEWDNX2HgTHaJviGRPic5dopdqlYIM/KPSNeaV+vj7jo9M8
XDvwpdk1cM8HnYmqKQTmGmGg6z+dMWG9jtjJ+p1h5MLw4MwMjH+CF6uxIMqZTerqd7BEMcbgilmq
8OvI3hpy3gZqHPzgHhmHx4ghDrfgo+D9OMpOrD1tUDTo5q39Vmz1kDFRy1vsr1jUmjkN1QrTkuUi
0c6ffxoV63Wv8anl8xuc4Cv1+2eVgOxkvYupkmYkYxXDyUiDESs/BE0BQyqXtIpyLjTfv5Q14c4H
Rjhbt2d/JXuX7QJAjLJA77CJIT5Xly3kZAh+USQavNMbNlmnzNnQxW18ZaeMLY81hv8aXwA8xB68
po5ThvXMMFCyafiwmjpDhnGEZNM30IEAwrpIaDhkUfLMlLkxNgQZUHhIE399JiaVX8B18ZtmUdjO
rcuSOhTLnIYyOlS3oeEGUpgcDbiMzut2FFsoB86v9tqKlfimSBtHrR4V1kL9R44f8gQEGSFoH1AF
rdu1nzBYOW+uLo9SM30cqYzGO+4vnYe/O9Z1XMO3Tom2okeWJ8iwb25lQHIpqevE0U9iZam51qny
qzMuErJh+h/ZdswnlEf76GImyB+i9x6zERru+BmYZNRubhedFINQLoICiys7ujmmb0Tz+Orh+ZNg
kaGNV8acCM6vTZ1uDcdCCM/gu5k1cJsq5MKLgLngVcAh+6DBYs3ILe43XNeKiU6SyawbwBNbBWGk
8k9VXDh2caHaoKX3hZN2FxN8pqJeup3+P2lHZI7qiSn3M4PQgLcV5/KnnqUQ4FutddDrPIo/Omjg
NittnZhrwfuqpwyUZXPlD1o2b8J0TS39awN2kXGKzk+7N6PWW6HYdnLGv1isFAafeBdbNFAIwLdc
Qoml/lpAvRHAnrkXSGTZvdEn+BZWjR1WSGQDY/mtTl/Zi5ZPO/A7QAcwgQ8KDziWgblwqPWwLOak
GLsAzNeIpEEFODpQrw9LnXK0kyuBqy3rvt6x2jv0U8fr4N8bJaSzOisVIdDW9QfDGFesvqmru1fr
9YGRm9xP7MpHlg2SMImwdoNwjKfc1QOx17RwkJsCsC3IIDSvKHCKVYWjVdAswLDqwk+1FduahQGo
0XMD05hiyBvRDdG1kuJqOHMx5wj5S02L/gXrj5YEMeLlOlaMj5AfdmnTM6JayybOrXKqYn+r6j5c
rJqlwpqBiSzFJJ8z0xV0xGfdnfa/4NqKecm5NMZsglKw8IrDkncV9Klf9DuZprQ+WAnJRXrv1zZ+
pEK3i+c/DJvPDeeGp2Kw9SscjrdvxarO9c0CmRmrhhFsbpcVWuP1HUtFeNMjcN6eXtg2ymZDbKVJ
GSsWafa1FPVz6D7Np+MK0ERU5k6Q6c8AJvgTqebomHFHxiC/+YbUQszof6wqgU/dZ16XLThrbbtR
CeB2W0eeMyW4eTF+9WnW8cB92gjNrdv0HYXliIitXSBxSvIxKcKqaB0FqnpMzHH2q5q0LWkwpIZ5
7H6NmBRLm23Cwh8+Cz/xJULM/ZOI+t5OPjst6/run+6NLSaYMW823dBLWj4E+wAvO83SfiQUtyht
OEAhUNqxMFxDLMsZeUP4ws8/DlvA8QFkczx5haM9i5h/JBfSzz+hTeh0DstrlAfwoG/jqLfSkTjT
eery0wkwYgz3OapkbrEMaaaWx2pJQU2XUV2YtgyE4YTTQrIS5Dl0fYs65IBQ1Gh7tlwKKjOQEzzq
K0MyRCgCbLm3IDpLrvCKjxOKKE2Hq8UoOQIN8rHPFyXeMJlrcnoDk3vFWM5xpRKxzVN8LBKEKxd6
EiLVCipeTMgNdD8MAPW65B4MxxqREG35Go0KYfONsw57V6SXzm0tPwPUo/71IWnnZHdehiKyTo8A
7dYwEmm9xdnxul5ms5xjr6mh2LKwmSUB6aSvv7t0NcbfvZS3UaoAubrtbYR6diZzCdWuVT55L9V2
7U8WfcTviAE7IGhV76zBUE0YV7g7W72qmtYBl5PkcbMAVcaNqFhjCGm04GtAgPIqPAfduvFjMyhw
8/VHUKc62Hmk+CgP0IBU79tird3h974VzjN0d6uffSc3yPviGrkkWiVVSsrzH7KDH5LwHRcg0Vsm
7CZoC8ACVbeQSNfGFMgcVVhfXwkpTbzs2s/CP8pcONqacCPQ5F2BsIgftl8kzx6RdZUIY13bxVgI
ypXtRl/cpRzAtmmkclAuWabaGM3bC7d/RvGQFMtRbQOv5IwinKGJMEGvaFGOowU7naNoybHqfIJz
5PACrvJxEvb0jc+IL91MmXP9MF20wwO/4N+jx8bT8DkiwN1p7rR3qps0mRVYADCnqAw28v+d/3/a
pqcwIViJdaAM52Zc/PKQYigkb7QWZEeSvhvcsUhxpfvyq08u/YNmWAW8+Pzip+wGoHezv+/QtJMu
zobgriQ0sT0iAzDQECnAhlJZImUZlLaot5iWh+xhGA8p9j7lZvDOS73apvgHVo92NGTOV1mtoj1e
OTV2CYDbCskFknmT95s/filzYCH1eIIAe2odTbASREE7uTcVbsRb/hXYhg0kshmWa6XO5MAGAVXI
ATtcb27bI8ZiW4FogZ4XFQI5xGppbEWzkCg8B7OLja6PdfQVI3Q/bT1aeofJ3LFcAfCXiW9SxnUn
p7o9FZn+Dx5WNi+UWHpUV7tnCfNiEQF6e6SI/Rg22ojdQ+b2Z+1HvFfcZGtfSh0djYRdUmTzIuue
iFPuBgUIFUIxHviiEU/gTyiBfVCOQk2n3QZrVwQ+IQPk3/JRbb0LR8wewprITrRuyYMYJ13ryusT
IdrlNhBaizH+TrCukAEa+7bJW2vraaGoHsPB3pJpU654joaQp8FFMjmimnQgiqBArqorz3D7Wr8H
3w1TG0RjldBqHMVfeAbckonr+DgYMkFGf2JOND1RUePTaDZG3mR2duEhmiRRWblzvLC6y+8i9CSn
KUzMWFo52WdDtR94vvrYUVVGsBb/zt+LmbYNXECttUUCEp0S8RFBHThKYkJX9+zeJnPQ2N15jyK6
VggaI58/vcVkgfrFHxOhAX/NBP5j00MQJdefCwxj/BnxjteJNJr3SpxEmTqzuTpQj8gFgTunEYw5
1nQRdcekYrIcnFBlygjlUhZvToasNd0DYr8oOlyXHwPXMTLe9gdTJNfAKx+kzt3opnHA1tBwUYyP
9ggMTl5dqKasNhkJimZ5qlE+lfMEt7Fuqb0d/NW3LX5T8Ij+DOkkxWAbD+X01v3F1qVvwEpZgt0p
6CAUddWRNq2KNc0eXBYZO2Bge+mTwV2dM1S2u7ZUnynbC2ZAqkdqsT8okaxGheBjifkwfW5JIMKP
KVkhwrqPqLWlrbCZIswXUPE6vvPJql7HrZmE6TzACxOqVbNqjlQSP12W3gbbVtES2825FRCYQNzh
XmG9K3/MRq5pO4gEZdpcoZqVaqJIiNekGXyC5eB2ui0C8TjDO26Ti3KLxmJFtd///8dQtAbDo/Y/
5sjbtT0W99gQU9sK7F9gr0ClKkud4HLaYjJlscTk2uperCmc68L25DWrU4rKUvmMIaHcPu6oKrY1
VWw7WH2434My8pfOB4et/0QT5GCj7QbszG1Xox8Ov8ViOVCV9ypjQ2uw1TE2kmceDW7sLg5vidjG
tOWvnTeQW41Nz1XCwnm6umruJiJFa3WMaaas5oWHjAcLpjd8KedKlgkzmBhllr8BSXWe1fIy8Whk
vy2rqR6TdawJfIuGNpYTwEvF05h6mwIiWoPdqeZWpI1OebK6syiAG03hYkLR9/NzVwnfgdEq5TN4
yjZf/U7R5II73dE/MVYRUF4m3ZTBwR+2LHJfc2DsFjwnOHBjXgR2MU+M7vfQoBBte7yo6TbFnEGc
hYGDrca6AedcK7KD6P2vS5W16lYp35LAFyr8Gvdc0OCXMXTCPoLok/1iLCYK4MTUi5uz0F0m5YST
g2adDy43lNsi+M/a2giMNLlMUH3RqvuShhs3FiH68bHQprgGJ0nsHuzw9rWRxv0jwvcS5po7gNcC
fgjupNzrXVjGKVhNfPaInVcbwfpTKVAXSTgbuj0MV1dQRzh5xaQfeqq0r/CCAF3cj4ithtw6uwy5
HMY/3MGGGUoNwsMAxUAUfwQCEBsPurkcM1YlNTl6t0SNvrPR+gKDhfsVegkbK4Pr4xE3sCdxkv7V
ZZ/Yhh0tC2zMWrm0usRDbNS2IrvfLr9dgzKUq9CTdqbfcyvOlnXB7dXPqR9hxAw+IifuXLKbXp1L
kJqELLveQHalTh9uBOB5lSutXlBIDgx6KQNId0vR2GCGXdAPewS0XZ0G+Hd6WV3QOnLx4Gqw+mmG
9dUfwM0N7z2p1UfE84yxbMYmCnDvHNINKYlK5RN6pAb5pdv+Dnqp/XJzI6C0uowxMha+d6DEa3iJ
6SFhp4bRCdlV1mAasaD9xFAhaBwGQq01qw1wH85Xj34iyA0nTQ0T0IXie9sD1CTJ3W3wqHIeTDbA
NeNSk+dWNaWz/4sD6rj4eTfQvWSQdjyN0tGNjpipofSiUqN9lxyZRZ5vQ09Np9LqIyest5Agu4pp
cWkpYKDZXe31Ntd9E7A7WCLodrgg9/BuwCjpPjuNbNJ5CfSBrbX1XTjd4icVizM92XYbzYyqupy1
MCJnHSghgD12SdUh8uGa4BmBoAsgx0OhWawQmlcmG2rtw4/JY+JHYyoFAutk/UeFZh83SK5ahvI9
75MQlXSmtXqKk7rHoSIKh1wJnmEYfAAhGD4qn9dHV9eI5DXJq+h6XYpaXSWaHmnvi3QLc3GXPqrV
LAkXM6b4qW8HUJx9rBNz2t+nmcPJ8ReWZFFL4hH7zx2e8dOoefPd+mzn5GZQxPtGsghyRNbQIH3b
gMx2lz7GaWo+z+WFRaQEp35HGZZ7OPE6t0DsVid6ji0awpZuStQvB8vcT0tlj+AvUC1bGBrVCW97
4EZAbluCmjKvt3hNsANU3RDKh/DM3QGZnuUxl6BsxCc1D3zvFJo8TrZAkG2Yv87ASpTqk3mNkQIZ
MWvRP/7eTxcfpgkhK40rt2R5OMM5EbKRkMohxj7yUmwQD4DjzRB+tifDeH70omih1IC7nnfVTHfb
9SsJHwp6tHEpTcCT7xcFdZysNQac3Jdo5vToAHIL6/23pANnd7q0Ut2HblnHblkfYkQtT8/jBKAK
WnZX90O0m3D+zt0IsZ53+v3deMDCBUzCoz+DDz6K0Ek0Ij4oLUjTf0EnjCCufjD0fmEH1BIKRJt2
K5GBntrpcItUkevZxXhNhTfNyiR7Z/f16Q10DMnE4LkJp4WleWf4ew7KxoWdfNvbhZR8ThAgKzCn
GE7fPDCxbDtUQaaXvIxW8nUvqWUb7GattXyjvYtkuQB/5Ag02Q2MwnA4sK0XUguDolXRIjpld2y4
VH6DGTWzeTTUUDYZTpS398LQrinwN2MgkgvTWNbKXhbm743seRSxMVfTLc9g0Pn9n38//7Ogot5D
8t8LL0IZmG0cb267wg+k0LAMaNj+w1rscBi6ZUmtHJLj03IpLqnF2ANxhchPaC5EZX9rdM6ottrC
4ytyQaubvce3nGxSY42CUpC7WrK9RI5OlaGfsss90uflk/aolt4Rw5WkTyUoIHob1/FaUM4rbc/7
r1rO10JQ/1lPJnF5bYgiQxgBuv1BIaX4RA4eP3doFKlswHGaCw1jNX5bX8HrSTHSP/ssGdEOJKtN
b/djO+M/qK1f4tVSLDm8Bd8VmDT2P2NjD9PlXb5YQiyLB2NdNzq/5BH+UuqLRyh95MNQJ30Kq/Fu
1iFappXDpYaXbMeYLg9souMTQVhWN4UJz2qULNV+jQj9EIHHQnglW+QmRqlmAtKiKPY3LCLA0UMm
RYv+bNtjqe8mLZFsjaL6jZ1N6UALJsYXtA6qW9bDWGln2dDulg6XNAQbzI+qeJGjuqftxlf0Ua38
OOHWLSpTVjKXuGrAnvJFjZSV3ajhm/CpFBkIPs4Iazu0BK4v6NK5b2Ksx8UJJCPVSHKo0aJMd1LT
XwKsZZ04suUab1up3cHiBuFRUewQ5q7Mgw3LaFaux2iBgn+FmbNWnQYuU0GBw4f6LPaV7seAyeN2
KHZ/kdaAUXoLqon30juc0Jy7Eh/tV7l6WmN5fCQ1TIa6Q2vsdTu7+Ya1B4Q61dacSp+gADJTY9PK
NhXY+9PSc0olLujrEATlzXQ39rfK+Oh+K6Uy7x704vHaeHtaIKEz7uq5OoBbKLOR1g32D+Rgx1J2
JexpsWcJmbjdD0lLlO5INGWD80IxAAE4BVmuPgvVPTl891pTA+KYz/8TI8lKCMmaNFUXpXr4xjI3
jUFoWu3YkQiFYa65tUuqcVFBUFea8szxLOp/Arl0fU+9a35JtkncefzVL6/tiCClrYTgpPo8iu/u
jk7gh4+fjmPJcUfNTHg8l0++43RkdibYdQyUO9WSRYbr4ZnMtvos/mwVIvms/gUfwrNWIjv9U7Wt
bKu/aoBR2wFQG9a5u71Mi7kzomLWSdkZWM6eeycMuIYhh495s3d88hCj5SgWCcsiV8KGykr4O3FF
R+3k6yy3s4h4dQa3PF0AgkZcWthL8IuSPWCgp1eKqPRih/k3wWAH3DTPyt45UsyEegfs6MirAzXO
FVhWvNj1DRxqx9+xZqpuHilbkeX5vIprGub4CNnaynlKJnlwq06eNL85FtX6x0fxhIx1LpILScIu
gULkttuJYfjBwlxXUpxsjtdeTlWKs2Yvt/Vjbc4YXSHjSE6ArQaWOgTXmnof21r8WVgPVkvtOanW
oB1slSSBupjVIsrMfv8mBVVn2cp8wQ5FIBeN9ygYCxVanJ286sA9pjaQDrPiAtryR1mil6PiMQlR
2Um6XRPxD3CIo/6lyouGuZ0iUyqiYlhkuGoFwxqMegGfvqRhD0oIaU5cwOFZ0njvkXzw+xLf+Eoo
8XFzxRNIn0htSt4b1rHuoJtKiEPv33NFiy/U+t4BbuQUPbnndSEUfqsFhODHcGUl9JB0ZcXWh6mb
CM60LUuuWWKE/x2HFkwPubAr4ENyibXaQMHk/DwvQzRSYVdOxzby7XFOL6KLvEkahhF8FvXU+bTV
UCS1nLVPWPQoYQW5+IbiMpQgWWFqJQPkwIsnKoOqrzbUPWIoXVHjdFqhhtNeqhKkLQ6Sq10Fc+NW
mQF4I6RAuZWQSZFlT2Xl8MnCJiZi6lKbwzLwZAvzWQohHQ2Eick2+FKDjdC7US5cx+1WBvwdlt7U
v27hwv0XyFOX3geaLX60yJNTzzpOfFydCt/hMuH5XL/J+Jd2pCrIjpmN/zmm19Ed4phjcNDbOgyW
lbo4aO0sLKH7w4Fgwuj0WRoTIyuUNMml7hp3GTtZ4bl0rNUKasbH/RvWp6qlMinLM8hqgIcNnZKH
fvZZWR+wUSnFZ5ZhnUAMisBCsFWQZbKHNuSmycvIryOA7CizbC7w2daT33MiWlnyp3lR1RC5MMbC
yaZNK0sHnWse2hvKsWCHvI4gVBR/qyCljbjzQWrExl/9vVOIHyaz3eNM96jvDtk1ODLRxQVc0dlZ
YfErF8ud1R2EUT9D5CrnNkadjtyLhsCW4HwQZG+KPwDGgEnLzhCLQaIF+w99qCPpdQU0HJZj5YSl
zJji4ujrioWdbb8aJHnoVuYvxeJjM6gDLJtVz1XRDjSlpnC9gFY6gU7bhLfIrOzW2y00QkV/i6Rk
M3XZqUom3NrCOn3I+e/u2DAt6T+UjfDsoDPZzY6QDsmfXUTjjyrvK3WI86sQUnjFiR5jqIn1sqHs
+tvs/YDNXxpCGeCnNDVmPYpfjCMlW/ruIkbsdjBCpPxRH7IXpS8OiMSQr5csaFbkjBg+YoeaCI11
koDeuphlrxOYQqvRQveDvAG5Lnl6gG0Nskhv+i7eRdzhvCdBXJV5ZSt/lNv+NEm9tndLzF3vUluO
qBz5a7DRIqnyB1lFfB7dpJUTwPE7l5PbfKj+2cyZnbW1HaKPk4LFvI4Wk3FVQWAw6eUpV2TKYW66
GzW1+RlEevcgFe3dMSQUKLDyeEvPMygbNzUno2H7bA0fPUnA7wfpLAaNtp/hK8ZERSbXVIkpgYbo
Gu9I+j3IifPdvWWWEu1FpytFpcaWH8AGMrIHIlE3bi61X2zSHrVjJ+WnV+pjMbGSN8Q3X7dq6Fp8
3X6XUbcxJNpmzVyArzhx6CFNntuFVhIT/BizL07hh7dy1Hi+HIPjyvBn1YGsMzYwePACW/6sheKS
X70zU7U+xCkeSGBeXPJSe+AFFI403OJw+zv1NfhQsugP95TV8K/aRB0l3UGLbLjK0PUyLKeYRDWr
XdP6tkURaRaox0z87kW0jySAsWNC7PFwbRQYanWPcDXCb8Nrp1dflLSlTuBbJEBxUtuy8Um1aUvl
6YnQ5NzY5CP8aR+0cAmXxCWjD+6ik4mcb9XMCTyKsMDvtBirQAVqkCjLFnbZxGBNLIbZGJtFJzH2
f8kGsrTQodeky/cyj7Yyi3bOc/fVYUxKBh02Vq5dBfJG5cL7ILqxh79xoJztUcLFaUv7STjAaJgO
3a2WOQiwGsxzkcP97JfSajFOdXlMwDaIe6yz3NdzPHCXwXxEvVO8hZ/bW1FPECvOlrx/ExyaBQAL
Wjt8NwOHo+DxrHqfuyznSBiVV5gKISmIt4ftNUjcbkcTPtxzqsK1hOvyj9X6vNP49dgqqSy+sJF0
9eAQ/cum9XmJ6LqfZH6ZEWi50AiYuOaZcGTD2PfwVpTNc9rPfcd3SAjFn6eAS62D/NtvwQiajMfV
vk9QClHWWsiKzoVqk3jHPhoJLc2DPxHqVoN0/yqCzlJprXW683BcANm9n9OYJ6WoFochbxtANyC7
D8URkmiAcpnhPpqK0Y0IfotkZkuIu6zUiGqCgQk3NJxVXg7jhozQPLrZb+0y+ixhJiaVsRST8Fhw
FFjvM/J13E6vIZKF2n8SwF8zKXwQP46QYgA9Qn3hzsiiXkfpBK///70/np3QjHzEAKG6oZ8XoSb2
PfLaJfuW3KS0EU0voTmyHgY2UTmheUOwN7/7Nn0I7i9Dwz2PyHgC2sfxDC930FjDZlJr/iu3AxYa
zF7GQrwa9VQioThLb16zLMrq95E2uwmiooRQproOFX2X3Mct167iQQ7bMdvkAu3m5LbQWXhSwW0g
wC613cvOzkBkWk0qA54UvBANPzslA6HxBHJfSu6h9S4TCV3GQP632ZaFcp3ggynT9qUpYEJUhJQW
C6A/YKaXPfOCZAa4NNCVAhajS4j56OvlOSdjpZRbiDN3ZW/ZE+il9G51F6rd2Y5WRAcNOsnWxBnJ
HYl5igf0F2W7F2e8QXDJHCJR5+FV2m1j8qjjULRji+byBPwGkTK772j2AKol6VeVPg/ZrJ/3LvMY
iEgqfVeqUFticPkhC9wSCgsJJvnTWwabrPk7b1GoceLf2EX735a+0Lz6rj6Pb1IWopDuuRpfr9iw
69ZAtM7eSLcmKOt0YgCc//Ps1LqgdWU5RIaZmTmXhkvGrx4jYOdogbNiJH6+l9bpQwQY84Qp1Bf+
bQAeT3W2JlnNowgwFkyliDMEl1WxxnZ3JWltClU+WIr5rM30puH5f8oBiUNa3NP9C9wxwKprJfmL
e1bm1D06umkCHy6EUIaXlfMFzaKXM5v/SkQ+/hQwRRqVgT9t0oGiycOurRADA+ihRyofAXZ4Ugnb
0nGUsI/NZUbH4adtz/7RaeH43tRLzOLqH/nIwxsEauHYRaHkUduEqHtbuWLSVt1o6nzVhS8FR/qk
FCgQgqtY3/eMWRM/47Jtu5asgc37ySw6GwBUqPjbGwgNAklE2GFgWeVi20ILrjJm8nhAGh/Ia8MQ
/4p/Irq8wXzy30s29VwU4d+Lfi5ki5y4CTX9yLY8clGtioKDM7ghmk6e9+gGgM6i1bXqym6XfD3s
bh1SBs2XvJjgQLzvqJyaJW7E9Oa2HMdNuQ5+r9repCihoGEDvYMJZPATdr5EJTkkJMLt2hEwWQsr
sdLzlNlC4Wk0PgHFEjgdT2UOzualEQSN2tTUZF+VqshvN5VRIorX1XfWAC1I9hpFW2/iVwMLhb+H
DFhAvoFerd51Xz7sFSIGtkcwIpB8Cge32Qmhx3RvO+ddQhJ8NmzKjegQrg76KVUBOkBCql3gLJjG
3fnDfv1L2yN1vKZFMzyfWn0KCydP69RJbpmRRX2zDbf7f7uyaXvrD6yWw4ARCNGK9Gau+Mxecjcb
ytXJaSRHoUqfsxBqnPriJ6lM44NZGVeQ4uwIVuIBWcCnMlnaumvAifOagpiI8NV8l6hvH3F/BrVS
x8E6GYONBizKeyDc0dOTpEtH2RpLbXXQiuObj4+J18VhnugHhcspifoVYbtXEzavkVBoFK+i+Eei
cf2fAs/7u+32Ck30x79CtHVYGFCRCm89lQeBjWw0Bjw492mCFuR5m7Safp5lQRBxD+OyRO/1EkMo
Nk2OuvRmMY3W0OO2OkIORyouFUzvs1qlRDlE8Ew7woOXCAiz6me9RTtRKsddzZRSLLwL1b+QhGfH
Zhj0urYYKVLqKSiiWaAgtQGgzxKva8O6lJWzjwaba2yFKrqAVDm//PpdtLa2qb9W5Gh5WXEk90mm
Enh7y5gpL9SH00ApG9DLZ6cuONtdQRZOmGpI0fQxemi9fV2I21HuLjClYdsmkqwtSjwMi5qVLFtk
qsFFfwozyg967LUnAxGvOBR9ZhI0Cr57XBeOs94aQ9LEkZkoroUe+qGeod3utzWUEiWBRNeEyzDs
1SdBKo+WgyLdlJixo6DGg5HJXEFborwU6ADOmriaojYXIT7hG0mKVg+vTUZn5rZR8501zx9sUGOk
Gc33CEouCGWyQK7B5YjLXxB1KfmoxHoEf0MfZvae64MZPzHVRSrMWLTRv4NiAC7g6IOyjNy0M0Iu
uicWP8BMkXJOXshrS6QLB+PDHaogdCuls1z/ZJTlDqm7SyjXXeZYB8mcu9/JLhscJi8drQloGw+e
gKVB4BALWt+GmlxJftaTpXr4e94TrddUl5lAv4j3CNIqvS0ZGta9kb8bAp7DeK+QvOeiFfi0cIL7
iSPmwfO5hql3/uXYQpYDs/ECz2Sjw5v/eXRtMvmIyLrDPksR7G+VsXC+8Li8v8bHSyFkmCz3TPIP
3wW7xrdPEt4DgbUPLQAsFt7C8I13c99HGyieExo80UdLzy0chBgKTQcoKIxi9dh3vn3nAlG3TJg0
B4CP2wja2VlPKHge0U4E26QOjrE25GWnnQah3G2ch+c9bFUinwjh/TyLxBJrI8nOfLAqb8rmXWP7
pGMOH4kprafLoLCh8vvSVgYTFuwtsZsrZ84SUzmvOOHAjKo1UMaOSMOUESq2qgwMvtf9jkwXvE+y
bUhzVUqyTCoeUmT1/30rg3Zad26BlIsISgCIR4QqHWSU7r0GfodgauDh96FBynv2Bo7NOP7w4qP4
yaj6wCZF3h07co2QS6Z3+po6DirWo83kBdcP/xV1MeKGTpD/eLF7L+yIm8Nspbxk1yjg/0sZgNTK
g7I+iL727Zjj5a3cf5gpV7tiERnEE1JU5RlXFblpYaUOKwNnJ9zRo+FV1tJpUb6LuCTGv2jC/OFm
1l4EBbxbD38mXRC5c/ZFQTG7fYaw4uYnXPaQn9zK6iLDWpof9mpxWUWM5mP6jWzvUSXwrUbMF7Vu
1bIiI2gU8mZM4EiH0zdjrR1s3NIqDu2qJ89/OUKtjRvQ8IDBr1jidxLy/hFYmmN1W5VX1JZA9Ywq
g45talpDlt+SXQJWoguru0w1+zWv3/nKd/JfOL/SgdQ8s7KgfBY6gTQenczYwNzIrO58JA9C7vq4
Z5UZIRuL7ZE3WRWAkXsjO83Stmk9hhuMSiy10H6Y7Qn7cSXALCX6eTFJx5jikhZSnK27aYp+xrvO
TabWnxu04h7mBye4PDc3C7CyAcbxRDIfjf4udW14vM+3A2kl9knS5khKbaRHseimkdWY4mZCsNW7
gz5PBaBnHv4sB5rYyBjKdGt90ZAQxQDbBoQp99hIAiq19RdXgmTrGZLXAQ3xmGr7d1dP7xRXevyI
DSblIcMrfkPBjHw62Uevh1euWFlKpDdaBX+uiGVLzrcQp23IhFEWxYEa0/+Fuf+1SdpQ2rpWBjUn
9xH+Q4rF8G8KAvgcR0sPT7j4NHqwg2iRm9hwkuSMPmL7zqp+dCABS58wbVwGTVB8wMCGwC1TRZa4
7orm98ao+53Zqw+91c+SUXvm3xAmWPzUANPxYPDsGO7UERf5EzpzF3Lmcc6cNxXesUJ1V9pUAiJk
gotuPo3ODvOTrkV5HEWwTSwtcECS8XpMeZkSUxNUDdKr0NYg1HZF6zYK49sBwGpMviN4wlpgEu4b
8HGLn7+r3T4GLM/xJN6fpRMs0iBMgM3lCD/xxd2kaL04ldl6Jfrt8+hPKo67vBty+T6VEUBtgfp0
RLxJACc4TaP/SnI88aiA3dWoPdb8kx7Tnel2UwLS8u3YcyIyXjwDeTl9bGKKPaFrWbPLemHpq5Gr
DaHMV7n4dcLobZoNM5ncUIeECpNfLebLN3MDDdj4eKB0nxHnJVofh+q27v1X7O5VXWE99Ic8CfUj
RMVyld4PDPPEXaNLyM4WEMh8Z3764cNo1fHXiJF3VTpHCLYb/Xhn4XvJPcWiN2LM+ijQc1Li+3lC
mPIk/PaksfxR9ornXj19n2J3FkGt/l8fBYuhKp7Yz1NUARcHK25fiVfqLj4TQh9uDuktcXe/C9IP
azZ1FR0dveL1dwGbNWcfICC+UmNycPmHUi//uONXuILRFP6xpbXCCr7YxeCB9cueEYQ+SImdf0Qh
tdEHGm+iXocbjt7Boy5XXB8HLzsC97SnGs/yHdgGHhsl32EvnlsvzLtloQSFuT7+6H1n/ajnutf1
DmSSemVNMODyFgbwIj9GUsmPTSpk9xQnGOax3jD1gAU6Axi2sT1Sq0E7KLcmYPgq7lHZz5AgFC3r
1osDECv8HwVPZ5bmaT4nSH79ytnCDo6/1dX7UnDlPX397eEUQA5WXAEgtYB4qjmURF+yKcH/XXiT
KfeXpigraz7zSQRkimHXZEZevqRh2maLK16m/5IXTzt6Urw6dkoczgV4bo2n84iQmlwP74knWnQE
CQ9REwGJ8TN0KRWEN9Dvsf40IypD+4GQUBDZQmhCJzfZXEBmaJmBr/QAHN3xoH6Na2p55AYr37uo
UuGU/MjHndgKqlSi6rRbOYhssF0CTHaJmkzsL/J4Hb8Vgpno4hM9q9Mz9Oe2RI5Jkhdm6VGVT4wS
dY3gQ/b1seMFkYmgjSTZ80YVl4qhRsuinyjqi//Elp3BMaO9VgZCQaojd0NLLUgCbf+RBT7GS2KD
AHEr+x4WlrGjbyBP6rtzw11dDnJek7A5tWurHyISbHtPXj++Zzo7C1ec9BMsuHiMobno9iz67Tok
WFCtaUYIPERkU2dxr4vHz3erRAraJf8uD3I0lFfZ6jGcC1l5WgrrqpxS8u35NS52sLvTmqztwIII
Waq0P5mNIPXsQBfZ15VBErYT7LahUrKnu64ON7tB0r4YinjCkEmJfkc1J0LfavdAIyQd4syjQyt3
qtH/Ug5WMUOfQ9fJR3wg/rwnfg4SubxvlCH2rO6r+mJ+AC8FC/QLNHwOelRCXfrMxmwl4hEVZAa+
RdEZqC7QGvDo3Mt1ofAymIPS1ccYjuTIug9V4umGzq8woj/fO2xfuCENL29TZOqEi7afmBjHc8qe
BCPdUBBJN16gsdGmkoqOVtSDl/34fTd7VO9w6KnfdtXP/mPjVFC4BakmVSn8NNHGpYPEmwQCTFzd
BnjSnOU7MBOYSXe3TuXMz5Daq7ou5MoSH5TUXRUp23mu6qn7mM/kbQBnJqp1HMPUG0fJsmNDR+KM
95d6lsAPbmEau9wODkc+cR3t7rmjg10loOv9EjAOxLUnd8McHiJMUDWponsllQHWx87gowIfirvm
6+biQkGR5Exbg2eZO/gKixJSO5tJnYvbQMsVwXgR1ssgDQwJxvUTsPddy1QEoK5V0+LiFPGyrPNW
zm42eoHHX+FWPqUmdsTCWDTQpwT4or9ZuNK3K1HPRpVenKophF1MboAiwCt1erGwO+Axm/CepT+g
boNHKisd3DeavSNg5v60qJTgIwaWbDImr5q2sOJYwdszhadBI3AEAqnyYttx0mMwL08Y1Qt3dZJ8
2gZsdqui+D5j+YWD4d+0vo9E38t2ui6lB96SJcq38UmNE/zdfstfx/lD+QDqytD7zOQ8wgFXKAEf
QTPvOUiLlYQ9gqCI5c+iO8xrjAJWpUcNfmqskoxHzk4RcOD2wW10C7TknYMQ0MgJCcIe0ncCFp/y
FEqSowP0caiNNmngi2cDQtZCk2hzGOhAuQzfPvs69Vid2Usd84+1TI91eTzkGqxYB/Ot8o+ZLedo
Uy+lOR88oXsyZHfK2NYO6Nx91QdVUbQuFColy1gG5ZliQVap6RF7KBqfkn64LrBXwUUPLjB6HkFP
JK/hfyaRVf32bmrZJIxAF/RGCM2ux2LhKBlajCa2AMa/UymJ0GcyWRxXIQpMzKaZji4uM7/0MQzI
E23bmVPKGBZ78t77hP2J5b8rjNRbIOZcTBB9EBITkg8K2w3SW7b3ZMrRvpEaKA5TNPDiiEH0/OcZ
QokIieRO48+QyavPDNgIhR+Eit29MGy70x8+ZCJ2Udzbei3cDkhLsa5jvRvO+C1v1Hi0Fy2rNCPL
kXlUh+5WrkXRdl32GRxckVJpE78sN4/SHgxwPx5QZ8bfIIvg6QelBMT5O39WXj/+bgGBcrmidHnv
h8lMSQ7iuWjLkZFX2bsCJSF2DytEyLM33NR8X0+I2aUmtqLPRSDOIBrCZCDBlrPFiiRxdNhlopyo
I9AT4uTalqFGW6IlybZiPcR8KzeXzJ+WMSekYR8BA208twJ46coW2AzdN1aMkHTLBLWd326ujJ4y
5QG+nIVzNQCp2VWlaTazirGGmFpwQ8DPzz4BlPGsbq2ur032sSNxHvN3/qA06e+QNdVjvkSEuHFh
Es+G6eL48dpbtU/wOVi4c88sWds5Oxnor6egtNQTkdfRWFsetv7D8+kIGwxVfZ+sUuLocIrWUv7J
T0aCLQi1+PkiqOKJbHkBsurXzN/UIO+05YQjJXJvhwpFj3Ezs03Q6w1Xf7zcYTYXnaDiIk7UriaL
O6FEsdyamiawwMqwP23rlgx+1Agnaag/RTaXnWhTaNQbLPTi38+7RgncFMPnEdNcBKCyRHkNtIrl
yGJi6JbIWkD3bgglEotPp9zJxADBJMpaErO6vbG/uvo11U+G2pJpDNy5XdpJq51OFxSfPLIufNAA
xUCiVAuLRcmKsSJjY0lTwJBoOEb2S719vm39gBQZNzGMHGu+G5Tzdg8geU0pUWEjceKjMsn1KrPW
5ozJQpzRz9RIK611rAe6YMFOICQ7RyFuX81qmeTBkaXtFirRjME6p0Mc9kcVn3D5zTM1k7saobSO
wHhbUoV8WHPrrxiQIg0mPhUNvaAX5ZzVst9FraSx8BGVaWripQiKrKbhVo/MSFa+5w2jC6G/TUgh
L1XngwS9OAHHxpplmi0twthXow3bHJCHtQkRebBvVzecYkJYzfxEYwkNPAQHclQVCEv4BZJuE1a3
JFDT1lbdDqByfdlLoTzADAuKqvRYNyiylMr9YgijjT2l3KD9TmXoo6Ie8ST8ZCuFimAu89mei4yh
vQ+CwkqnUUaByNowkBpIVdI+Y7X2he6vioxnNJAIMwy205I0B31cYdV4WNMYzdyuoKKYGxNv5hiI
YNECYm5DwFyCAWkPN7m69BauUUuTmRdMoyucKgJ9iHzA9t1/m1ViXvxqEF92g8Pii05q90EpmtuN
PTKeSDhF1uKTtknVWPfSdqBpEJdecRLh76DTfL37iuQ7cyX3NuJyEtF89HHLd3RD7tk998N97gY3
BopBGOlCoocBEJunO+ePFz9Gl/e+sgTMfU7KsNrRlnAIFjGRBC4JmohhmCE4RkRQKTn1jLBk1r9P
F8Najlc8wvvo5n+5+B2PQ5aukh55tco9o6lTmyB1G5nnvtmSMEm0Fm74luCR6R0CB7v107p/mwaI
A8/YZuAO3WBfVidQeWH7x56O+qjXIa75vj9MxySXcJEqkTWVuMjFPd5Lisjz81fn8uLX+pYfF1g8
1aJKj/SNk8IfWGyvLypu1aJ4g2KCA7zS7A3yr9i2eLqzZK9VqDAayJCOXfBjHBK/tTY16jQFOqmn
LdZDgihk3FqKX136Q5wdn0GDftlywexHVu2JVyHZ7p/jAXs9EDm4COj6UBKrGuaRsGtVIgaSlCeo
IBuxJNiS6FtfCaPqKKYHxbv0c0oBAKXzf5p3bQA1hOzOAOYUv9Oz/Ly73CZNFDghzavqt+5krvgF
2ZwEw+elCdTjQ+tW/sqfJCgVcrPhmggWsiJxuYOUFa902pCYxVG37KkltmcuR2veCyu9rzKMqAiY
c1WmprtsDkV+r6nAznr6i3yNt45xC1/INBHTN1ABsDu0+JDAmdRThyv9iWcsFiJsrD+Qv/JaKkim
MwiuQuZEhXzURIX/v6l8RBTdHOAzRpG6MHATA6KjEGLQ/ZLOSaVjB2Fw6Av77Yh+TlhoF/qjauGI
3BC0+lMQlxWijdtU8BaSTReQYtZADP+0kuiTkOGJDR1zdaLN3FAe19WLPAOm8qeoTH/U8EeUqyxB
41bAyMT9pbW6K4ll3G2Fdn9kBGIZROYjsRtA5/KlwkDF8m3nzbpzTXt447FXsdLXU/w9BvrxHt5/
eS8VMvwjt687TGtD62z/l0C5fs1pcOVR4lsxCLE11SCNHJbWhS+Orln4LpGWs5uRhlQ/2XNXrKx9
egqThn5JJsh2WRTYx2bF9sgKEnRzvmROxy5UgAhojrC2zPJyS0HWw36z9hSfV0JA+PWT9zZOccFr
que0d53q+4owjNerhT0X7n8w7iRR2oPx3emxPKYFKD8gtUgW69rrfJESLppyAJDHoqUUJUTGI/C4
BcdgJIHwq8eFt7Egvqj0fgJ8u032mhF1iSQSru7jDlwl05Wu8ZcsA3N+oiQHP2BttPE8oCEKG2KB
SHcdDPkI6WXXET0DdB1EXHN7UTFN47m1L9CDsQJ8khwAcy/TcdzFrVnDfyPf7W+Zn/X5tqsp5URe
botqeZX+bed/Ehjq5p7E7QuTgtnWZMqJjt8LsMfi27ryExcA+DIN3cjfEdbTsfMhhSpdUA88HI6I
ETAvXTb+lhdhAlf8XZ3SdNjJHJJ+U9iXsxCjIEnFrOxSndLzSOcLjD6yzmYpR1D+1OR1sW68LqHu
lWwWFt1iFCtYDH7BrU+FF4nGq0VVKHi8vZ/48emUlhcu1V0QvjNfNgGhQxe8uvIgcyjKCJZa55yd
HFXmPyccnxgI1eI0Wf0EaVigKLjaAeAuGi9nCX+JZ6cXh+RejWew/N3+oEeJUCIlImwoNQubpsk1
Rq9WSiBosP6NBCnl/PfbjOdeq4ilUYbcbsEs626s6LcPOPhLJZeQTs0zlKr2UELz4xhhEEgtf6S0
Z8pA2ltaCPceZyMkEjQqvO9ZQqcK/UGba+NZqnZd+Evd8ycojVoSosw1oeCKgxjUEPjO7adFeEel
DvPqTydlDAXCTcxExnEzZZNlcBoqms+auq4ZFJg2f2lxv3laBIh9IF4dLQOCVrPxigGMuhjd/YTk
0nYFvfikmUYoRFT3DL4m2W44IK1akQipfyPuIV1gPyjt88zR3qWcAWAAxbz9d+2q0FIy4VGBGbTK
QR2sWDtUOuJ+GzxJaJ/EbebQ89AlSnCcHsfbLtpLo0ZL6e7I6vMfPd0+U9gKTYXPaiqulryOz1i7
gxkYFgbfjtf3NpHXa4utCcB1vb4ILbKiScSue1F7lFcjaW0WqMDJYNVtecgD3aw+9GtR158CccpQ
cAFr7i4DWAjXwnLZz7+wUcEm5oMAhKuFkdWUSh9I24d20mHr1zNZFsEOgb3WZkhlQ5QNqjgqMucB
C+lYz6dUZiGFW9O3TIgPNNAAsBjykV4KfMzq9yH19isFvcgY6kILP8lJNYc8xpQKi//Zp8OygsZQ
ezOC+wayoOYejOCmtt0ycs0NQPABAJ6u5MfWOK5JLLSC69eKXp6GOq5nqrgo51rbfE74fPAkvkmX
sp+nAyxoEm9ZRuT4WdwpkhTaRUAIfN1TK4AYtQ+7CfUoBCXx93YUJtpGesZhbDl3irqJkFvMNCfr
LO7xX1OoL2lWRDbSnmtri0gvYEbV2kobaNsCHf1mHelMbJ49GEbNlP9HVG+C+1kP3Q+YllhZPuvC
vv646EmXlpiMp5fNhH32WSWEr5cjZfrmKb4yJKHHBm+U93R2nSCrWU2kJFuIKVqcoFfdXkXAsUVT
gnYIBHbEh27KygZSPzQd/IykKpv8DDFXECbbVx6TJ02gff4+wb2/CgS2PBFtoi+jlZPLM1Dan63k
qp3F7/fHY64C1Jz+t/leO941uNOG5fskGiFLyZG8zRqKnjKiiYFidW+k+6+PaoOPFiCZInBC+5MV
DVuH/JIwKPCQu7ZpZowe2nLGsuWiKMlDDagMbs13Oc3Uy5Tql7ojfX57JjHGZmav4vfcxYNIyfAy
LeAW8WDu/28jjA4vi9lw7B9RR0sxmAxFMDzu/mldsngC/ZmG47FP0W3uquD4zg719ytajCbEeDUa
Qj8qfj/sXUhLd3qWmF3W0m2EQ5GxnxH7nIGJlU/c6USchelg0eBPNHuiphcvtw0BtovRARx1zR+4
43l9fUxTfhwZorJZgGHL1W4EUFvELh8FqNWMOFFcMcT8kgJhg+DEQYNUk1J3lkfGJwy791pEtD1H
+/6jPTewChjVVEmixo2wg92jdc9cS0LQgRzI0WmRfLPnU9hba1QzyL8L/Bvj90CqR5/hKBvUuJ9d
ymj5GEcHIVYCO3ZAl9gWc4VtHYDDWO/lDaZWS23tvDRH3ReMx2k+eaDbIqTUxia4FkL5ZzhoLm4E
1amDlXztX/gYd1Jm6L6NsgxuoCizepW+1q3P/ArYsUs+hlA/m1LcLB559Fb9V7vcLh6sHmH2RvGR
V9052RPKKEvSjofCIfFaXu/oDGAf6FMOs71068qApxWouHmAsc3x9UiBKNHmXzUja4YVvvUEnQHW
lXUp+vj8K1VrZ1hwyywOStF/s3QlHsunTkNKV6EaXIKIqcT0Y+PpPISbWMGh8o3olEX1qaB3cBKW
BNwM1Hp6o10zxKJpeb2d2NFZw/tTTp8x1mrZxXzJeaDLavteJm2Gu7wqy7eFFMi+ybDDbyeZ6RhV
OhKSZJEuWjnp7MGgOrUAl+kfOa9lCSu+ExC6J+YGxINBfzCs78vxTLbumgO+tHIWs//++XPaJtsf
tLJFs6H6VlkwH1NXMNa50fUsODzwG5xXiNpTYRb9a154/lRoD6wPt6vzTcV09UHPVSfM/Ajzn3H9
PFjkw4GqFWb33izfaPe1UgdEvq2dUr4Q/lDQ0wcYcr0ma2ZMRZ5tMrjkNY13x1wbRPTOorn5uDLG
S39wYcxz0ayFuNazhN7rMCoxOtuN9EZeWqJDuV9HcSN3bXlF559jI5g0tAC16GvaR2imKAY/HXCW
Zu5nUsT20K2YxL7miHm4+lylFf9XRxWmNoWAbUkqmv89XrTXMP8BUXs1P4us6maImEjkbey2GE32
SAIaxpeRMIbo0KtT2jYPYHZVCUUsQcjEGyqpHo7i3Lx9ozoL5R7AmzB7Yx6qQRnUmnnA94TDaCXF
qft2ANLdDzzSSMao4AhbL87p4iBhDY3kYC/2CBzSWaklCTFMwGzu6Ojx5cx+tEQGVytomA2oV7Pt
CbynrA84lG8xUL7tL2vVr/kyprrM57mHVTpMBQfsiWcu+HU7ECTAQZRzlMZ6Eg4hyFUDga9g56hb
Kj9FVMl5Y1dkUDwPndpZ/hkevyhsRAuypAFr+V+atjRJyh37aRzCboBwdiThF1UIJatviOX74FFj
DF8S0qFL2gAVFN+HTdaVcwan7capsVv4vzfyDVmGqFnYSx41KvSYPZ9q0oPBlwKPPqoHTEm0gdYL
KlqM/eg+hViMl7TznLEopv1LtKcaXEBaAaHW+D+a6o/XV9lxzed4z+o/icLXKrbWfb2Hy4wqJdjx
AuAc7WI60moJ3nB+sVJPHBX6fid5/s9ZMIyHvodIdj0RIZRXlGCQfoDtwN3jjhdq/cTQjXh6XjwV
8vARIxGJd4UTE0PaS9/+6qnC+WB4zUC9R90qtVVKef/1UeIJTLzRl1zaLT1/WX4eQw3S4gJ+wDY5
De/L4pfV+rnm5whqe7yaodolg1AJdfoG0GbM4oKjR7/dy1p725+HshWE2MfHoD1qB4ZYdtzvX0ks
lICQdZ9oPiCdt/E+vyLBkf5DimxTbyJVV3RseN/LwMaa+Doo7Cqt6/PnPWCK5vPx6FBWflwkq5nd
ZPrQyILZfMavDZKbYbrpQjZxLTXHIc26G+oOwRI4egEXmcQz+bIKeTvuOxjdLIW+liqIVBtiSVdy
OJPS5XwhBU4aRBFKBCHNLYeHWiyXJzsP7KFbO8sw84IQ/yCQReoX48ezjS8BqmQG4vjrYQMfToQR
b1ScjW4HOm6m1ypw8dWJnjBLIGLLYIhd8LLPrcmxu3CM2QLee1Zke6aI5AEQOPCJk6fHrqZLu44Y
m5TeJUpUs5Y9nckW2oORzxT2GB/oD9Zax6wOBJzq1le5j1oZUgx3G0KGmi4GA6iRoDQwrsJhnWvJ
xov7mqdrE5ecShWuBOSbbw3JDEwwEGRZ81KLLbczz5EoRL2h4Umo/tRugXnSIdJlPBN7i3QlDz6Q
TXb7HhiFig4ZJEwo8nePWyBsT3UTvMhP85E150b0/hKqvtO4w5AW+OX1xCGQa4qEAyh/NjMhskPB
7Bji0DM6nZwHk/mMnbV8pnfzaVsSYv9YfnnF9DXb2eqdd9cpDafGi1FTbdizaq2i6vo9KkybFZOo
fdSQNutvu54gdRGuon7OKzzrUgulO7IeMHzO9YzOdWdyBq7PcLydm4teRiRzzQHBD2KqURtLaqvD
9VKFYCjCs8BwLkt61rRo+5UWBrMBjc7KSaj28v5Go2B39CeVZW/w4qzJfEQ5muu66xl8f81mSlrm
5DGwldhQBSVoLijC3I+wbwNnK3tYlvFwFnXshSn2vRF0nCA9onfMy1PhpZKQgS7RSQGCm56Pa8s8
pZP8A7PtlwuzUr1G93xft2HdzpniP/ejWg2Fj6KiHkiDhEcUQvVSDFg1CybWES6dqVstDhGudln7
CVav7P2hQhhyagWq5n7Upcb1Wp7n0zPlqffci9A5EV/pXhqb55bc7PcbriV7Dgit03kuP3Pf+8X/
B3LZTUQMbaIN0SGh2f3LYVvQ9AGEKhveOjoD3e5YKOBtqi3i2q4/HoBl75tiHBW5x5F3LVbw+dyn
vCS33+5/5VGck7/iYKPo15wfLm4Mh8MtCfR5bFeM7ID0lY6Sduse+G5t6cV4tLA+GXEplWun1NfE
AfvfxUqKS8jNs8ktk84EUAEh6r+VXMnB02L/88h3IPo3ceErtUwmSXdVEc2bSLK1dFx/69wINPdY
xRnyQbhBMJw0Z47UrMJnDV/qOG+qKo2fbJubsX3h4n9YVsQJak3168cOuDfo5nlbBGLvdC/3hDU6
KMf3f0JuJroZ50yNjWLrBnUq1mEEIKM3OpjkZZeJbdVW1mfbrMr8bZV1iLrty6TsVPmgLEcmCO1N
Rh2AbKKz1xjlDFEaxDnM6ky8ZF75/KqHQOa7ub/A2Q+g7sQJUyNziRqHNw+JRzjtcFMm9a2qngDk
myBxGB1HsiOSf+QjQeKGqberPvxlYNIySao9y9JMMiLhG05exeIM5ICOFZe3fslixchPpzgTYyAK
9uFYUrHO2M+Vz2UrEyJWV0rvMi1X9CHqQSacE9BEk1beKAdgJ6PmiRtTxbfknja8d6uVwBT4HYkS
ie0hdhbSAKX9YmY/0w9PAyULqwsEIxXl9cBJsArvKYg8+X0oyNsQITK28Mgig8/MBrkZlAahd8Ev
9b2IH1OqJ6vyjgD9N++EpHd/9E2CArj1e9l+5r04+B4MwqTm0TWgFdSfZwBqXpiPSRe0UW8c3reP
Rar/WhHYMSoCkXEMazO8rnoQ3GaXrmgY4HoVaRsIal0UANrcYuIrBtlwnFWSIVn5HY0Hjo/NoIKY
vv8ruYHQH1QGM6RI5AsghUjQmnMMOFje0M9uDShQZac0TcwIDTP/fiPbDxikIQ3JakTyZqnSyEY9
T/A+BxnrL/tAmp8437NUGyfFX+atsIOMSguGfkYfDWA3LHNINHsHOYDW3ZN4qBabyAwn6U15E/w8
MD7PE+W9iQt2bWfw5jxaniGo0DNSw+5S171neo9zxOdsUKNdMMI0iifORdX+evDRFVLdoyX7bK4N
56tM4RKeKBdxBHk2HXbou9W7+zaLCDDVhyPAAe6RRKokUSCXGls3voAetxhstlzJUwW+UNwm/iRO
8r+HXtn3Rbt3jdieKowNC3f1Fg1Rk0rx9F3ZbscMm4EFjTSN5zPYPySdAiliDGgjNzeKHl4bJJ6K
UuyL1WwQCBJffzfaGUJv7QMUwp0uOp5nJdMI15GiEfZ8nkQT01P7NGDlpVKz43rmImPDd2gyzdgv
+AP3WcwhWrW+qsC27WWzRRfKwNnr0JxdrbX7MXvO4jskCp7nLEtur4j8bm9/+UnnupLzBLZbu0+V
saMzH0Rn/gZeA2OKF8VG1BaqiUJzdIC+p3/3ISWt6TPpsn3I6yTjXJe3aVNSPj+cORrfqs6KIymz
jZhuUxdy4+VqndnRFADC0QVlneM+nrroy45UXQWEB6BNnkPo/zrzzs5wrAO4HUZVku3bEviZcrXm
aTuICzz5GDBmVdW4WADQtKJlVBhRSX/re72qIoDiTrC/0WvjVdMe9Sikq//HDVJadLyZzA6VXLxt
whRnh4fB1RbFbrewWSZmlDqa4l8lBZDE8SS5fClA8XEf7kQLESaRsuHHXY1Jr0TJE/RvS87+FESP
8VKkJqBe2RJ9hK0/R/XwdOJoLrdxzUOCIFchCJayMY7pQS/3WIhivD6u3H83Faeywxd2eMqQgTIG
ZMhk0Wdl/7QotVmgwEO38Ve+zRCKru0OtFfJHlZUVeZEyizIV7qsBGHDqnZEbxlTtmcQC3bmF/Tm
TeqDcr9usOOkkTEo6xGjngCvu6ht9507KyyjVDdERL0e4cSUTY27ouk/NXwp0OnGW2mE4mtIbqcW
0xnOJ3GEUXviDJVu9K5P2130jT34qP1CZGo51hbvvXlvgl7aC7R8n3hIlLI2Ff87uMNqwVO2uoNI
doLwlVEfCKgLexE31e1v/1V5ezZvYJaucdYQr2mCslu4OM2/rSYQOuFUK3n1uEXnoeGhmGZHnpmM
mOFaoACx+gvUim4ISLIcflzQxRkCOlD5xj4WQrL270JyGxDto3j6NUIoiUTX4ONF5YWh2ALDOkMb
HMKL9cUmDVFzgpwLpiyXErZHNg4yM7myxWUf/c6yWgTi9t642yOR8+hIW1MEiZsI2dzD2YK77Cny
4G4f1a16LGnv8YZ1h+3FR3kKvMRQH9dOpFoAzd5qo5Duc3M2eJqIvjmQtvJjAg8PRHxeDkLzdhCT
k/VUuBAyv4aQnNDTyG0nqGhNe4VvT5/NpHQZhLOnjRqq5RVmbY+TvhouEEuOcGW3LYA9pSKH1cKx
kqBrQlKinChsKa3+XQmZz23bHbvVgEwwNvwGSWecKJNYBgq/pm6EOxFlfQFHv/nZp84+vpJ5weWD
ZZigzyo6WU9Fi1sxiec3Ar4YZkiUJsS3uXjjg8VtPOaDVLU1ovqHnf4pRxrar+AgHfl7el4Qgwl6
TjrTcxIwBR5V4SlcprA0XHr2iaThsiLLXRsvf62gpHax/XuRnAh6Et75hJRrjsbrDBTyW3fVYZPY
6O0tHASki5lRjAagFjDFKNAM1tzgvcukYk+yr0dXfqaGzvD4/rgfYDfsbtkGS6wdgk0z+qEQpMKq
QSPrfYa7ft2BHB4YllldYvUUfBwJynGdx/lXaHGWJL6TNbvClPvPVCdS4JQ9XBtoMf7HH2mJTAct
gOlc9Xfs2nys5USTu8xZsP7LKBp8F9Ph48TZQijKWc3+p9GVdATVe/oTIiEgDo5bSDXnoL2DpBbW
jp21wu04PzaTQ13BKq4oXGbMIjeRbw7CxlV/nxqrTZfMvFBWefroWmIhsW9yO0wCeuvmCSGoBqs2
Tqox2X4f+AwlQWQsej/hLihRh+ugKBv5diMAWN49XhgzclF1E1B3jMWz7mbdxKAspbuZ2HlOavIb
p8n7pxlPWUfYGgv2mwsLjfY/LK7YZ1qXoG45wfVyu2OOCwu9W3SWkVHATMpJ6duJ0Qkp3JavAoq+
LwryIbUJsAZVTL1EU+uPzjBhuJ6PsBx27GdBv/4sDNsuP6KNnPmkRpb4VZqDiXRam/q1khDt999K
YqTBJeg6bQg3b80zELZTmUL5KPFy7vblj+H+W/W87bCoz/1JsfoyjL/q1EhzmRUcxTTZY2yyJT/s
MeoLPfZXk1fH2Osjv3TB816SmM3yXTJXFVJ8+uKzWPnhEn6JKVYr/GyXc0UruaawBPXjwj0+3ce5
8kL+gcByv2Jbj0bHwTxrCPGvX1vf3P/M4xqp+CqxIbP2F7e1G1VwcmF29N6aCwZPj/zpKI5uNB7x
HvV/9kqXICn8lMoV/gIi0xbnaIlSFGYbBI/qntStEC7dIOOM64NQlh4WLsm25j+xAN9SqqvUirNb
+Ro5z9iMMuKR9aSojB+yq60+7QKlkJakCgSjv4e22iSHuOTuUsstY5iQVp+moRqLuSkXf4kdu5gx
IvcWQQIo7hGc/uOfaEm+nZQ4PlxWtPW6bwCBrB1Slsgz9UwmVQ4fkiClMXgczBybpJAyvwJaDfXH
KDk2/WGAm5xatntN17i9FqceQcZk5A9O7IKFY5XLEbk92qhH/M2k2I3CsXw6JKw59SgZ5CYTTJKh
xhvHB0jA2TCIiDn7V/mwb9M6ybQI3qPeu9uVdDcq3nOOhutLggqPX1h1zTUr61RK/4unDKGWB/hl
THKVgVpczOYaM12IgDxEJDkor1NpBQSgerqTWCaMLlyBfRRHuliyxbcsZ1s/B2UOL2Dpi+xhx4My
5isGzmhesedDX3IttlRIQoxSu7ztFpRv91oBLheInVaBG0tGfzyV8gM+7Ml7c3aUhWxCOE8yG1Gw
rqGy5Kfdz1m+FLRB2XTvfTjUxjdOyTg2RUQkwN4/3vSfzLvskXxBwKO4DRNvsgGsT2lg1OyoPkrP
y0aVLlwstqUo55WVSIfpbl3ufm2ZQU8rTFKNgEXS2vSQhvjrKh5vAHoM+CcEURzx8tkWAIrEqkhy
FG0O7BXyPVQvN4/Wp58VxvcaqSgkMM8dpit2IoVmnP6YQ4Ol1lxxFoYCKYYDXxxjXHy1KD8uFk04
/WgQNTyrXYDVAdBp7h+HA247OVKrXU7tZZdRdUVid39MWKshf34zOR6J6AZ8KXDN5KZnvJgUaSZA
5c66OCTSEfkvaI77T+ssH1ojDMXTXdhPbrMhxBFEfRJqlG+ycV4LGf5vswZJlHtNDoZdJitfG4w1
4mxns1RUsXCgGLMha40Ten4qigJmpA0HTm+s9LVuN+4wdh1Oul8yt98GwAxxwbeq37JiYeAyR1Eg
VOUOlKd/ZJa8Z0jopVt3fQWT9sZPNXG3/F8mUhif6Dz7XvUq/7kJt0l7EWhKoAHfnoN4s1mKkqla
J/9jjaknRWkUuYkrgHZNli9jow28uZd5Yow2NPDStECHr8s0/FJiB24OTEO04YfV3zHLwAwQcVbZ
fdu+IDCAXk4HnI52PJEkrO9yY7PISGqGDMlNIgxv7HhHOHHGMZNzTAdQ159mdoqCZQ/7e9QyKkjK
iGF1mzxfXwM0n2WHdh6vL7AvLXMepqJ8seUiYq3nD0IHgDD93eHVabnWmB5eQznVxF077XAKw9FP
+cwdRXa7L4j6S+fXhlzWleNbDEh9ykK+ToupjNCMdIfanlMHmMJRmMJ4xCywx1pAG0e/kS+LhcjK
Kk1KSRZU/ybpLbLtdoNsZyGhKOY2deMUKQztry1wNKhCIaKe5p3tgX47kD1C+PRhk5VseNHMeatl
ARGdMoYymV/FLp5DNGwVDY+j0jXQx7bwF00BGmyeD7MaaaBOx4yTAjVo20cy1oaIzAw7a4U0j+0E
bYeFu/nLa9mcdFsvP9isKu9ts+2JeeKLrOvxcqCV1jezWeidkSLr/PaB0LPcYvJvIciCizUfsGYY
omgHBG8eyuAPTZnWkA8rUVz61CqZuOkaDOsrm3njuXglPgYSOcoAWevXQ2MfdE7FhqNqELAUgGK5
Qp4tYKYzSXNma0E5mWwZQvb9YJDJx3mbBnVQsDBzYkHvOdvuxsBKQFBSk8pbjs86Mk9rku3w507B
azXSnZJYzm8ihygB8N37BN4sFBPdb7M544sTcsdGMLYKjgxvt7D53vD4FfovnwYVoMWmws7NmnvF
7tBI64DfFTprj4qZ5MA4Lw7RddchUtSSONhnxybyZPAzzy8revvMbsN2TmRq5J+xMa0Zg0IPZV0s
5Um0mtD5536x1pFfe/mzr04lUE9z1u34/u4h3T09lwuBMmxO8ks+b5qJIjfvIQ7C4epRFpZGqwrG
jH+c8meZhegTlu7Mh1m8ZI84dWPHYD8FFycB8SsAyWQYFY62iHFdsUSCO5CmLj0oELpJI2Mgw/Yg
w6r5Pp6DCBF3KfL9w/DT1D3E1URz86dhl8mfRTtt+TKE9sGp3PoDqXD9JFen2wxxU/fQcjgXcbn3
yCebHKGc99/sjRe+9JR6xxnNcUH6bBJO5QaEED2G8LWTku/uVBos1TnTrFa7GI/2jWtTgyu9CRZq
kmE80LBERFhb3hrCDU3XhP30Tan9rK/IfWNjaLs38NBMtVt20nPA4UV1m3x/nYWRkIG9o+AY3K+7
jkXNYkOtPZA1avCImnGcmB6p2Rby9HFzxVfZZ+GGea81AKaLClKj3VMFvmTGhFBZ77LSF2Lho5Uj
VF2YEchEdkSBcBNqFX8BcM8RYFuYhOYOo5z8ilEsrkD2t6pANhOepbjevKZJJYzm2ImzQ3MOrnrF
rWXq2jH5A9op5TH0Y+jQ9HZUYUD2JnwOHBb/mE11ZUNIbAJzrVCGSL4XSaVsTynVFJNTb4960CdH
lJxJ/vldezf9hNLN3bEQ34643DqJOlmwNeAhJ8BlV5gibWrFkM+UtoG0DfU1rNYgvrwc5MidVYiu
iOcxwxXnExqiE/lE7SKrzvGwN7+Gss63DGfP9KQfbkj9bSdhvolbQw907KVE3SdQJfbY/SXpiBMq
KlpHfifHPGvu0+RX3L/CI8fg9WfSGiGV4oSyLN9uYjWf0KlrVKIx3KjQyoU+YtuFyS0IfekNYXni
glTJ3GIbeEGXuX1uTltaJrQVEajzQCZyF7qY2W6Ce0wOCjhDYrP6spjYOcJW6IrD3dJ1xFUO+gZ8
I3RZe0Vxzoc/M85ltnzxYe/3vXWKlTvbnFeTEZ2zXdj8L/b8eUzf3+gWceJplfk48hZV+z0yvdoj
kdCbJ0128wzoRmMyAbyGUgV+nbgQKeuFDrRhHdFTT/mZXKzAut8EEY6Xri4v+hrL886YxZZYq/7t
JrpM4PoHHr1eLVaWf5+fRqRor/6RLl8dXKPhNagPvmmU5QPbsTutQzOakSGisflTslw0FmFSUd4C
RBzOyWwrhWstdusEQIBWKdTXJMr/nbze2GC+54cvF6BGBfWKqT2gWZVU2LyGzpOBaYc9lhDlCHnj
Qh9EGuhDIPuUdSowlHEYZz22QU29HcxT0hZCvZIsL6f3JFBIgSq2Uy91p0/Uuk2QEthCTWGnZJcZ
yBbS4ouJOe2Atyr93Ll708nWeKAk+ZpcbJduV+OMrYMheaxbequYXL9s+HDYyQhxYl822ou2rr3F
bskuCj05U9QSWltbexF/6+a+MkgbMTHuV8df1Gz9CYwvLC8+pE4FURR1qTQ3oFXqc4k6JM1fK2gm
i2hoKaD1egxuaPIoqeEBQNF8KVLZvd0yU5tTZm5kae55ySqYtFSKSVQKslkQ9+pRKVK+yIDxUxxC
kpGsGryyCPmJvH8x6tNGzFMbTLHPtPHQQRgsM1f02wbL00nY7FkpekaKnkR3sHtntrXzNUOQyp4p
XD5r7ca35K7wgwWSq6ZOytHyVE4ETGTIyTfqmwSSBjs2xk7Ux0sIbMNL1xDtiDiatl5EjCZNgtXD
owiFVSu5VX8NK3bLpzRvyKIbmmBRclSPslgv1vGij/gOOo3g3gcyqzcDNMQo5QI0mQ8FvFRGk8/Z
6O+XEogqffqosb4CTXmqzl1UHFVYFwQSCI5ndBnLKM/qYm+PqqRFUiFrOzZU9GLREhtVqd7kQt0t
N1CdZBERo8Lp62dunZe+AxssLoF8bzpT0HcxetiZE9wawJy6ctMuZ2pYtqeAQctRKWBRH4/cuXOW
69qT6+1MwbhrBfdevnDhOdx4qZt6bC/Mgfhq7U5UHLmfa1yDkOqCfwOKbU9gpbhxBrAVW0mGq7uo
RtB/WRN/PBhsmJCSIghTQ4fpilXqH8HpRM5/SRSkGVYicoLz6lb/WEhkzanNI7u2CljHGt1sT0ql
BIKY1uid0pFxl82q7oDVTeByjL1PomPpTW1msXfzC6Z4wCt3oUtYwOCHE6rdIoD4D7Vu5uyuUlmP
NolMt9QSdMVsdCtvhZdxWHh8uK1Rw42jTu0FWrnQ8WQ8TKu77yRGyv2tUiib5sKFhOTbexZVnYjT
60pM44daSPvxr2oLjRZ6GLwIOAi+FiX01NI3es7qLFEURIDfkY/K/SB7EkXMog61AjV+7EcMk4Ry
U5R30PKA+Fy8YG+2OdR2EWzlehTKZMzwpT52ivij4jlYFf3/pGAofxn524C43j3zTFz8BXIueukZ
wtjF/4D2+4vi/n10X5tB04u8RbNmlHvPe/xEHw818raRio80GCHhh63mwYbr8hBTef9ab4z4A121
hj+q/1QGABZ8oI6meDmmAP1ALKVIM0kF7ACi1UUF4XRnKY1+sqQUBE781hlVsFDbRgUOH82TquHJ
gUuKOi+bK8DfityaAAKOkP58wKcaIKmzORIJzgd4I7vJN+9JrZRjunOd/sfXU3f50wqjJRFz5gwz
wLBG4pcpmplNMopSVL2OARYO6MsPmUcm1xsPVolQJ99UqppQ/wml5pPvES6fmlbaVJuPkROrfqUe
Ct1gCT338EIWx6nTrmQ5P9H82BrPEamcX+f6Y/GbQDlyrSi4PhDjIYK/UZK2S8zsrLZxfwIVrUJl
cEq0MKPv2Wj23N4AylacuOC8QrkTBdfxBmaKJKeZ3DHa1AYkXe0W3YFqiF6WpQYVZ3CwpXp3OTMz
y0jaIYoSsEdtABgVflC04fTA4sVySlGcLeiGxSbi/JIy+Vlf0vdzhqBdjTqy5l+gFApLaZdP+X8m
1oZ8ytgE3w1i41K44x7DGxs1UHDTuaJaJDn8TCmUwbw3OqBb19jAyIfukP6gNl3bSxaXmUe7Kzty
5eHROgMoHjok14/U2Lo8cHWrGlSDg16j2GgBNojx7AhZCeYaHA8C+SZ+MqtvsdeSjrDIVuxzpBq/
lddG2yFAmfCj0IIn3eTVfXgikUsuoup0q9ghPSwy26MNOoV+5Pnv7B/dSQ2HUvSvjmooJCh8EL4Z
kJ2Xm7jl7eOf7E5XXqGL/K3vlc/mywC7hQTb0dWPYkNDwPF1oiUFj3SrdUnAQqHlk+vHZmrrarb/
2BJXEicPIPrsdTE2gDEydJYVLqMd1uOH3XFLFHp6/0kDCLDxOSK6Bj0pU98kPqcJR/e4Fm+t0HMH
jxqyTTER8PbUqKGZZyuf5EDYexdMSmuqHyISpzbw8V3SconH7nJlmfG3BaLDx1eKERv3asJi+K/y
Lv7G4Kl1+3aaHka5z4U+GiodZz7n2d9lF+tPVNwkO2HcHKoYQEOSz0jUkt4XPYxUcJPiRft+8tk2
qXVE9KU4R9Z1y6RHXitpIpTZN35ThIDsN3Jf6uMOhoM0+zHOPkvNDDlj5I9DFSEBMgmQy+ozUrru
Hfv/OUvs8eb6zudL0SbCuS5cFcEjVvYkIv669Fyty8XRbFeBViX0ZLE7DFeNvtTy18vx+/SgAZVq
PnxCjHz0VJ+KNis6u2ITt6IGOlnjf2F53fPOfYRM7ReR8roeSuVrfUigiKFp+o14BYYIkS+h51Z/
St5qw2/Efyin3XDaC1Yl11jiPmW4gMGnW9MpUXvpfc0SK5+QwMKEmYF00SjNX64WeXmJjtylqUHa
CIELZ35+DKgYoibwxGKORJ3ZruKh5jUR4V8o2uq+aCKWM8V/NsBimmSfbswmsrpmuXrkhwy9OJ0C
wdCQHf7PokvYsmiTlZuAJ/MiScgvt8pe2//rMbxEZvLRrjIuAuWs+oczvXX44HKC4nvV4Qxkp+Zy
HqSWRD6zNIpJFFpu0ePvYBIZyNsVCbaPX+gPUjE/9gqeH8BbAiaebP2S+KIhbJu+Wtny5xI0Fe1H
S+TnkrS/qFtq6mG3mgJJrAN8pOEnSVdo3jn7fNh6+9h4Hgl7TEiIKe0wkhtkpikIuStDHLzqByIp
3lu+5MSpJZNJEOa5EntLL4mdNaEbOoL2VlobG/OBv9nT3nTIVBxCRzz2Hiu2gcZTdmSLoGXuWEh1
XplID62z2fZL2wOcX3IDgbRAKyzv8S9JG4pMjlhmZWA5f08p7s26nAgOWE/g4PwiDeRPRbydIUqt
skFa2WcPWAeNAKI1fGGNFj6qMUzQICP4FWRkxbnaNmXSuO15iKexjiSrg68YL5cfcuEQesi+Ct2z
ntDMsUamSFIcokd9ENhuDvNEBo+e65LJTGjrSXugyTI9tSJCvlfR6CSpkXMdO9mUJyvZze3h1PdT
yIFWj35A6wkx1DfjUObuJmOB0b5ZGOt8VyDuCvtWUFiq7LsylfxwxrUiaaVyBsmsb39avBKh5lG7
NRSOLN27xqXkb0cE3RrkRvp5BtZPblAIRzED0YkdRC7e6/UzUIv08iuuMzFo2JgqKTth/kyaEloA
J2yt16aS9ntR0FU06IurwzMeXCcPKjnlFWkZjXp25+5joYAVV9i52eUu51iZIDgDQYWQtuwQqTGD
PNB21GP2eWLz+ueBsdWSoTcSOGb4zXyWpgD1u2XFHPm2Cv1iYAmpL7WrF0wB137YT1gEJl8mE4Uh
WRQutmEIbdj5qq+dQIiZd3I8M78QdieiA5t7PKsgnQk00cmMyu511TY5cKtYNN0kha2S1reiXtM3
zlYKf2B8M9lpv8a7cFolbnxHTmWkyBP/9yU6GBYHJdSQ6u734g93MYvMh0isAuYWSsTYhW8k+NKf
YewABbdpZV/O04gxXsk1ryqBWh8fO0BxpoYC97qhsPxhqoYJOOVnFDYaHS7TmnPIEBTiYlXM+Fhj
JdmnpXufWr810o3Rbk/6E0Ejg9S7w8edzE9QJ4xUC5SXe2HxJDzAsdl5Jz8kWF70IkzNGT+iHiGc
HUPKRKUWPzR4jqFzWn5BJUrqYCT5PICKvyYa4YFVC5Gf2o6h+Op1+vD42PJrpWq4gApha1Xpc6pV
+xpRM6i1VOY9My8N12yVjqXdN8u48V3VeQDzd+zDN5XckphZ+HLhu/Wxs2Emd8LIdbjKwpdj0Xsv
6j9llqm+wb61jIsUMdizavqvNqj4m780PCXUewZ9frXlpYF23gEaI3YJqm1Olhd9vx9zbVkSiv0P
Zp+tAR0+5/ZnWOVf4GEub/xgjkFVFezwfgT2rDjfUMKXDe95c++w2uR2ZMNxSsO9n0duJHAUacya
9zPsHnTSCNCq3juLTVsPVVR489QDLQH0O+8gqKEd3DSDBoJPlmY9hX6J+RfQ9MswP1+TKaQyNJNZ
cEJbJwvXorspVr4z9EyNcRGzPn/oFxGm7Hk8MwqUMbykOkBMyyrmf4cqoD6lSgMBmSBuZwUHSAqM
SJ0RW/kGkvs1cfZrzvb+SKvdsb4LnB6bWYAr1bMpF9WLwEm4FEGZf459w9UvnREpAqcwVKgjxRbm
c+kIc8GmU9OSvpfz2yY8S91UOxtHOLq7X4U9B7VROOf2jF57nTRy+Q0fIYN7xBQoPNvwxGCAtxeQ
dAFQT7PF2D0xwOTDkIWaSFYihtc/ahFiQJdiag5j2h1iBlsXDTfntOzhc98lGMmW6+LTBcQWVi4O
S3xavN7MJtqx9jcl1leQQJcNeizChOldXeTXJQHlwUZ1lEcf3PXWKH1mXuqKwMbp/xpS2pzaIkiW
gntFfKg8gmOlPhmdjfNzcDCmp+6/CeiQSV8jy73vRGdEaD1tWCQIFQGGVXCJULe/vmWSugUJ/+5D
EfzBC6LSnXrQEep+o99RZE4+ZCE/WlHqNLUC1aMz1QQzjvLkvXRpauQZDuOEI3o7/04YntBGS6+C
K56TP6ZYBgNGOWN+T1P5qpdFHxk/3V0mJSf3eHzDbfQo0Hu6kPKyzU2NC95ssrQaLz2dSDZT3LQq
GIHDu+rjp1m6Uo98mVaiRJHoaFF5HCLwCoatCYMh5bwAiQlN58R5ACtwPaJrCiU3awg78J5V14WN
WRDo0qKUW7obEKPWxq2T2f4C9jmdRdy0TYcnK9SdW5k+MqaCeoFVpmIgvyC6sftrnWGFjrKbCdJt
3hSARMmcetVcMsHOljWUEADG0JP8fhg6g7uogy0BDjsBBefvzdnvY4NKiCQLaP1MTEgkNg8B9UYR
ZmVj6YHFVadwa/X8VmrXSLAPGdIkcaO6t14L5XvcRzAoLrFq4Zb9deqAA17FTCR3ymxlkGsG/bVh
wpSPh51JT881d7o/x+umAA6Wth5ULsoo1ah0Aznmikdbei/hEtq5QhabxQKtF8DoTAf8Y0gCc6Mf
kKC9RZITjn1x5GpmWcG2Xxk3vczaH/gOUg71s0CdflJ+CPIupaX8tJ43H0U9IWLFXzcxTBJ5kkeF
J0ao94MAYQA8nEJAFu29jDwIbQjjYPelnDV2ZSvOuKzqaIkv4s0of+ghBGT63x/JiqnkvKTvT0Ej
yNBThN+UCNGIi3GEE+e40La+7JOeh/duWbN7EtosFbAtY6hSxiZ3zeYUGt53iJEqbHLZ3GI786/l
zwU40J1EQ3B73mWwEK66JhSZQt3xLYXRW4ceDI4igoMNChSmcGD2zKNPkJNE0Pl7lwcIaB5NJkg2
o2g6qxadCAKMuEJJsWL5F2rWLzVCM0/eCRWOuSHmO1c6Iqy47DqSHaHZLuzc8SfeNLXVcXnw2/Gm
N8gS3CLPu3r3kMsVeywYjHxddzDgmE0SfsMlJcBGQlyZLAHPAmdB3HTnzeViUqsmUEJDQw1sPSXi
AYsHhuFrLiHS96vjH1a+betYEmNHQxtyeMcJiWdDYIqGQL6ery9J1G7qMCPx5CApIHZUGOM7oeUV
ITMvv/pLPfWY7KcTsbfbh0Ta3GNN44dmh3FODvbUYiS1eGc/orcMci/VZyM4WOJi3SFiFKqcJ4rD
wlYRlNdAYJPDgjN3tDh27Os0s6Q5703JyVj/eXRaApM5NSiiwyWyUVYitUdb5xW+QoVnod4o8OmH
eQV5Pk6RAk1lleS+OYmmAtYJHpL5auwtjQCP7Q4iTaIAoxUVVJC43UxsAgbu7Fiy8aKhSxd0xLSQ
cDjI3dYZ5UC1hELCdOvv7S6S+IUF96XjxXbG3mMiZJ6pRrFypslaD0zcTJtpcj8nE4N1+7G8CHWG
/EGmGxUX7KGnKfNGCLWDLz7uvN/W9uH6zlrRmOUp139WblBLQoP0aKJN8pF8UCYtqNYnb85zMS2l
zG+/2zsn6Pg5BhMPPIBgllNpAjVRLBPesHTF409QSBTkcKiR9ZPwK4ffqAo/vLNvislL16XlFv6V
kMDlzxM/yissYRQB9FpkOFoFo+3fIPJLUkoNVILeeKL8tgdBNR78p3/b7sfHmxPyicBuzCZL8KBb
Viq9hDBCUbAHGl/itJz8qRGlwGW0MD+2d99Md1Y9QghF+wiDlO6MSWaTkMq7K8flszVCNPX5oQtS
IjB8rQsh2EoXFgqWNt94nkSZFYx7Amct/yFR73k3/W9nqa/FttbH5QwJpVo76tjPBvc6nqiH1LhL
nWev+dBSmq69ArqtCHEAG9wd3fEiJwVgspHtCrhFothrr7dWACGamwXPefXqQWtwpr02sYeNzK8C
Z29tQi8ToSJ6FUEkiu8OOfxiT3b9ZPOqm1fDPVsGATiwWleKR+sx+XVvhr0e1Rxz/AEi299i4Qx9
Ss6Jik5RB5AoFFkTh9RiJRjjzsJRhUkSBhTXG/VciLzN1mohfO+v3zauvx1Pa0DxRw4lnPiwY463
CgB0aMqYlodqf0Oe6o/xJl8IES/hh2UAO8vlIWiBRTCi9IS9l0iFwJb9jPmKpk+EhL6RjLnyxfMF
gCrRhEgYxGU6dITn8buTkpfKwrrbO//blShb+C4sTOJmGBxeFFuOPgMJF7HUr/IO2c4yjIkhYRbj
DCVdujRQ6HkkAtUQVzYBbC7cWotVtOC0d4wff/lEqhqvJyK039I3p6Jiq/PwgfYWk0Why6veETzg
SHVoPWuX0cE7znMWAUSEuIB5lxhHfj5gZ+L411DoKLH0b6Jp7AAz0LVby7Hr0eBT9KogrCR/sbym
NLxOV2q34n64G+JARopetrpN/WHNKp+3L9Jb1ZDRkxQtb7WDW4ZATFq/bk1ou3xGc7WqaSr7b5jV
uWjyPFpXi9lYtFB3TI7ExeeQhBs5MtTLp8FU3Hk3PnTdKCskwmWFhTOOA98SK3RmOVfXtD0THpAL
+KQMdgTizyrM4DuNGvwmsQ4cKcPPublF2RMgtFypkezAR9V/ppkjfgobdDMDfFRxaZwgLr3Oy37s
BEC+SzWSMgjA2D6W1sNA7TTruAVr3WPv4wj3tHmC8SOXiSlraUIFIAorVCY6bmN/64qHinj3n63V
agdgq0Xpr8tLAQtKPRCdfjtzw58Kk8AX8K6IxoQoYkov0aGJ9vqICAa0N7zDcG4RBLLpo9U95GZk
Wk+a/855IKjb/WtMgipm77FZHpIFI80SgyDya2RAUXNwxuyNfnl748mWEbUoPI2V3nQwsJxP4m9f
rtAyMLDOmmxEkJWI8u5gT0s0F4yD9RGIg4mYZml/5cABZF7t8wuavZ6rKwV2hhC56AQZLVz1OrQd
OVXe9Z5Mp3dwped1jfLuPMJGIGytJ1ks5YeH8CoZ27G/7/W/9Q4ICxteqmNikiUHROKQ8DjkFU17
crZA4KcWAKz0CCwXieUysIV+XG2+ax1z8qtXQc0+3GctdnzBHZWQyg7d88/BPnTCes6x+IrKOzQ9
2CZT9+U6KmiYEai3v9yhapZ3tCokDc7fdVlpe1YAODj+X/aDIhTN4tmzKGjF/KxBC3cHIT9yROZj
TUC3qZd5QeeS3uVQhnFT4ehwDDqdAusbTELX2DkYEdbas15UhJssjJ4uDMi8JoWl/j/SmXA7txfb
88AXo8CFE9RT5oOrI4UnrEFElmfdo2Eb2sQyRmMeN9hDkBvmPNHMJRbPSAS6nungAnmUC9iT7MwE
POJ1h0fXTkX1WU6B2POKwmDfslZSOuQWecj4UJUfB5pX7qTz0Zuz1ug4XWL3DMP68ZAzegFDgg7b
o3tt3QUUDfrZK32A4G9aw/1EU7T/q2rn7dA0ib4wngliR2dKBCAuAKFXPuSh5oqocS1rwtdt9ZjE
ytm3C9vqGMFe3XcjTcd99R5mqdLvXbHswIacP4oegVynlxyKF5dIkoMkHMFB43VYdy1U5U6TOa6l
qWXoDVoZpmORBbUMZ4DAJ2S8sweeJ2asrCGYVcVCwtUoG3vjdw1ksnpjV65sfNywZg9R88lubKJ0
lmfpg8wi9ZAG/xJOphpL7NdH7f0zx4VlnwpwWO9UhmxWv0ADMJhvYcM8nUvB52OoJzIvg+YlgzXx
TfyGvZrl4/37pTD3YFdGFOXC1lmPMn1gQOMO9Snm7eh/8CnsaOYy9DEUtd0AWGdgUVIFH0Qt0VGD
Eg2oKoXut3WjWDN5exiLRSf9T75GrOLwBDLFngLxLV1P++pHh4qS1TxgXn0TdROLSMY+JWmbxxkx
3k2G1Ark2Vq0afXB2xDrKRAhBoN3JIXH+CCvH/+2SrTazBGaXcwXtR1KUGbABmqmiPW7XN7arXQc
6ZjAbF9olQJtBXe1u+tasC8UayPlwT/qErQ/3pjzbQYU/ClHh8YGCI5UXTrC0PlzyrghzjlGSzaf
2F5F2rwUXSJ2YFXhKNcCesHplXSAgAVFCiXI4dRnKcTRUI4wnAHBMemo4eEiXrnogkwV/+uOLI3d
CYnn8tv1PCvFVSnEZXNPVbwcojSETwyH89+FeOS0ZOTOacRAlBTzzlWHxci87x77IrUcjpQjbKIQ
45efYfX/3mxxPE1cHuaGne6hK6tUc+Z1VGVBufALrI9zuSBqLiD3oW8RpyFxWkuWvxWYZyW45UsG
auQ11tOHpNGzwIkgt6X+TO+copdwAG5e3zTochgrc3nlvt9k9pCm+ORB98UeXO/w3e6hA5naZdGf
zy9YyIDbjeDXMgGA+69n4iNuASAXkgxm9YPBKkMEHotVf1XQEzFela4vt/rK478J5NA5e/OTlHS7
ewzVPYL9srO4lOt7dxzcL2CX/HH88dPqQoyXHhhOUzvHfMTMuMbQX8Qi9w4ktog+Ailz46N/J/7U
dEoToobWuKvK3DZ+k/IWMS8lmL6AmDK+gE4LDSvwnKA9FYWx0PbUicBGj3mjsOHrapDUSTUbr89L
PKKRspXh/gzd4EmaNJqoJjdWuaHEaVqeWQv9JCPr5H3O1CLyqby1cQEfYUPc0mA9PDidxms0Rttp
UgPHG/cuaeu/AbicqFC2Jmq6c6GI+Y/7KXkEBbBRiIV+cOUpwSaARxx3zgUBZbeoQscXxSWoetgF
y4ksZo2FMkmG3iDFQwNpQWNW+AkYFz+wL2MnV7JIVKNMxl5F5AOMm3aD+rtcbsulh6TSDPYkvWZ+
emhkwjzgg9fIOaWR3Gnp1hpYnfHS/nbW0Hd7Wl8u8bfraQf4FGw2o3ZOegDtNoOilZbhwoAq8Lfb
THO9swMAdBHnS0PbnLwwIfC+cUt9xx+63BVxT/j+qy4twXtnv9LzEcJzRheF9mY/NVXrJ4LTTDOg
u/jrCS8XITgNnYJlbXJpN53ILXg45cvlthMkfnOToELuZmQf3Jz6YAmhiDLLxINB6uCpiw8BRkvq
Gjt48Az6TgopHpNOvaBgs2kcphOkce5FbBFsTW0sqz+kuyWq6JKFijoHjcvGCSvW72wJStRg4IY6
KV++mO3XssutNz6bum39iYGnoDPuWncsACE4EaW6TMmTuNvUynythOsp/snXSF/sZAK40gUgs2a5
FnZHTWnAKK3J0zvWRTQKnNzHuAhpRTdRjXy3thYKh/upsepPgK5QhKK0gn1vymemeujd7EspweB5
cbLooxGkoPPsy+ALEFBolXbqkL7YQGM9gqIjp7eOJ6L3bEDA4jhqYWb/+9+qyl7l6TKXwQkQPaqL
WbNkC4bKEktKczkmxwagBAVSYh9Y0YEiEwUDQN5Ll80+u2w1POJIi9JdZoNX3TZP+xLdC7NVJEUu
6/KSmthbZh/EzOjL7jmZ3goN8sRRyWv0/lcsX0E2ztU+gQeEma/KOMVAIC7UQ0Y/5S6GnGtZaQaa
4r8pYK2HeHaioteTLftgwerSX6bUbQbaAD8lp15A6jvGtE/safYpZMbk4JRovefj7Rgj5M1f6d1I
vnXAI/X8vUFYhp0ErDg7eN97iVGwBldzvlX9gqNll3zQP2WAZb7GO7scgF+bDlXb+rd9YyHLZO73
Hs15m68sC787I1KBKN+vVeNmbn36/LaCZekb+DM9GXv7by5cLrCy5LKMXuzK4kJRPzrMNt5TDxVm
rZ21h6MhEZLauRmxeLaczIHWwPBIWkbTuLN3UXJNeROWBM71q+Bq1fG1iVC7Cl8+mNsDRw0OUd3h
QmjTWe83DAZ1riFNl3TXH4WDxxmS05PkWOj8oTe6+kQF2hh8Fiy2Kdi92xhmV6JxJvH/jIYNazuM
d6aAmtEGNHoRrji+dFQC81eV4g/OG4Mi1Uk5ak+QnXRxNNk0y0s2DkZTAgkQ+6OOfYJbd/7u7zkM
8ZpYCQDdv7xpLWs1SXfCUQsyhE2b1TKmVFDDyFyBQuXL26hVq2M6N/jkoWcoK/PdmO/FJwYQPNHp
YBebEHXx/vDXQFaP1aMaiO3Upud1R7UZXFJ6mMqTjgKM2eXiW2/3XOjlW9udzBlPmiSFC7Ifl0Lb
KWSRV//GsdRc+SbzbuxNE/r27AUGQ5PtIL4RVk5HXaPa4EUGBGppMlbPw5QFAhc+4Og9Y6GMGmSJ
qTwFV46WKxqvUY7igs9m/TKpUejmAIIxgw4XGp2hk0QRKq3ZL5zfMWP7FoY/bMpAYHZMScIbUCuc
yzIQCQFXbs9jLpgryxW6fHcA7EInszXM4emJNvZ4LkuuhTubl/Q9DQbdGtBJ53lHa06ContwFzzF
QaL7M31pibBOMUCSz6f80rEfTCeR8SRa2ybxPjNFeiDXxvyNg/GQrIx9lO0szPlOQcsIOHYMI9tv
TTsoW5L5RF/AYqK9XQgrkL3vxJ8dbiGT/Ev4HtVid9ADESg/hmEFXizsMv3wGEqxvgwC+WHmxXm6
8v2ujQuwogQMEr/7IiP1kRJ0cFO1Y/gdEyds/3tSmZVhG8PyY1JYVattgnFAVaKIVhO3t2c2K7Rz
b+pMymke4h5JweJ6Nowk7eB7Z9McYjCn6CdfBeOtLUVN8vTfsY4YABKoQlgk1cnssYvGPf/Ex0yy
FF4Nr7kHxBOb1DTvt9nJbAB7KmyeE3oCT1tjnHoWY6bz2NBXZfiiegM+cUFxLmmWum8L4UZz8uxU
L1V6U5RTvhkpaQSTrckkao+elFDFl4DVqChFPXqO67KePgbLRIOqvx5OWzBh8arS4oGiHcm/UES+
upjcSw0D4fpJPutBHVoufwQsbCVAogPMyiCMcuYWLX7j9/MeFiPKVcAnCb5UCZnrmZNmXfEwObGM
bMjnRv4wr0SfyYVBcv84NVTVYAFRZ+gtV7PvvT/hMxqiOTvzFkI7UOkO5ePBfck/mT3G30iMucof
Gx+60qAkbzPdhyzCX1XZ6IYaCnIW10XOPmO8DhyjlGpTWLip8xx0HLGaHw/bzAe5qRqLxRpVcDzu
QxvABpljLcm6Vso/6KToATNHlD6GuJOt4j2eHh72La0U0TN+2gdmN5GmQbFa0Di4oNoP10aGYcar
I6wgqRe3qI+UcW3L4oJk01nbKYBaPFs8QUnS4OzGDnVWMHJ4Hz8IvQfuoU+8Buj0AATjzcMjdY67
xJZNLC+SrOZLpZ89pYCgFZVpA07PDs+v14Q3ZF3+OdcXHa+Sd/Ky1Ph2e++QbgRhzV8v2mOQPYno
OFp6XknLIVRVAisPjO4DF8hnlgVAb3q05mfTIbHQjuIQ2+tRwEE8Lbrp+SN5Hd3NiJfNQvja5PIC
C17YHaF9umYn7X8Z7ruCaLOfuNMSwWsrLDP7WdKc6zIj/hQdJSUc35467tMKFkHfPVKiLFwVT9a0
ah/QpbhIbri2QPW/VFU2Vw6pio7DTmZOq54uEttbr2T8QGCLOLG64a1Y/yy8dYVFrR5U7XFLVMDn
VxXMUt1kOtMT8jaUn5Nba47+nBV6bwUlEa1eROtcEDVaxFZPZxgSlnwTOPwhf3MxWskSekaQfPEA
Gd8aQXjlM1aqcSsdewNTJ1unwoZkdJWsFoEdgOSysXatjPlcMzp4bVnFvGsIF+lbLcf5XTEObh/g
XcnqeyD1njRAYxhitTYpQ9vYgWG9nnPbCiSvSSeDXi95VKPQMQ9JmVNfJpNcCgkzz79GiophLtBs
c4Ddo2WI3vRKIJF3RBHCH/FibXOfrnPphJP/07LkMSMolLlL90rJ6qX5c8LN5tRFXpTSfQDLwrBC
jF48EKE0wY8r2NrLyFoFpqtEKGRUxQ4+IFTYLS8e7T487HvqeTekfODdcxzQqB2k7vunZED4uDeR
joHD8OuUPcDJHghduMY/vEEyH8Pz34wIz02ZpcgCqnYPFGiQxmtuIYizmmBhCfDdLLoL5EDg/9g8
mPUOlMQRprCXUI8U9wYkbYHkKOCf9GTF57pyTTm320CfTcWjChM8QVuHQs2kAafDFHxVZu7gOLv5
KutPlPTGiStnrttaTd26iHqgm4rmFP2tRJEI5yLwNoD+23/iqAjOL5wPl3lSLAF7jdmloLoZRmmE
p1+FtBaUImlVe6DACdUS/HQDLMGlPki6Q2P7yHNRU8KitgcB7rpojkHYJbwqeOvA/oMTGnvGi/6b
qOAvhpTKwZRTgOCrsN1IvJD7vaExvqh+fjRvKT+EvyQnMiBeOyCaOu9ajzbiw1SQMFmqR4tfl0jp
DaXwkgsZawx5jKqkLD/zmjPzPt2mKn7HxQuFsBLEmtBpiTP+zpLqgK6HzMKHI5dd162wzDYlXIVP
dpMv7nNPIvzHtE81ybNIBc1AGO2VYAsAulj5xN81Q1DnMc+eL7aPavV7nowI7envWCEwEy9EGcOH
IqclMTmNg87d3WRICGoVlzZ6OJsrQcVkXSaFyVEsi6EX9F19BIbdVGZnG5sRTNXewCeCQRQDkM5G
ZOIoPs5vd83qGXewZh2VhAo0RqZDGyiHhm5FezoHIsSbWt40B7vsUIN39EPJukyIp8sJ8tU6zb7V
MR3ilQG+t40Plc3FSCYQ+SINKostgXvP+hPu/gMQj2JjMFJMVT+TS9TtQnTqwR7g5PnRfXTAyWKn
3eLBrRzQT2E10gqKBgSPBMJSdKS8XB+XhkuZPVAWh0suJa/gimLSz0SKXF7uBHfG2Uw93KYssIu6
FsP8xoxG0ucb/cifKxy1f3wYt+W0YkhalSy4fgYlIWad9xapsdpIySfGSvitmvpZ8v58Fy00wTD1
s/X+0DiHetgHXxXELnM5DB2XJmiHKUufvrnF646tjDw2cCAZkKf4JqBvVIFGL/iRd5OgqAS+Ucsv
uvgJtJIAAoLyolhSo9oJZikr8lImd04CVSf7hbcOLKWEjxvXQzKGEgeG2OEd3ESH0M80TqbeyUV0
7sgTTRxQ6IHgjUKDtKFkI8E3BB6/7b3u/XM+0FdX1v+6EoebRj+WRBFT3uJWnBoseahaIF9Wf5/A
tIgHWtO9QSKcp4LQDbinwkUfYwLaxfRCoZCl1NgAptyXElB6kdzFmzC6ROQZwY8DbRdBzof7nQge
fL1JUz9H2zqC3goTkyMdXZyzHC+70xo7R7FuNx71zSqr037mz244iwlxQn7JQn1V8T4Tc+v8eAQF
jIEOV/G63JHfjnDGGXN/vGg2AiZ+GSJdtQ5Fquwv2nwbGOG1MQF8OpUsLSu9rz20oygA0CdzvE6Y
7IX2jor/0jVbmgUoX/HI3NXMkHvzhfMh9+tN78jXCJ6CDuliBUIix6CQT4flcAkRQr0URzb8L0QP
pF09s3Q2H4EGaW0TU7YGJhP2q3bOP89tIEEZ3WsMNo6Z5Fv+CPOLmffYjdm0/KtxdWdXu6CxkR5o
yekxmtRH2BqN7y6LmTzYeiuLn5nPid7qBeez4RryelNUh5j6YOhv0Se5JBHj5PTa0lzpFLAECABt
jJvmC2QEuC8yGJWQuEC9HLJ9G8ZGX/YReSi9Qv6d9M3TH84Ws4Ue8OiOs0OI2nMyep+CsCFJDbrs
k/OlpI/GgtFC5/wDGy/Q42q25BqjoLH6xK664wis7/FuwkoSAqe3Jyxp3uP2tYw/7ti3pLSoVZuV
pvIdl+ENjX55Txd5N3FpLfKiVchBz+96JVJCRG7GAesF4IvCKhaVJ0ARxTUgSpsDmFZBWIfIenfB
bO+zTXvm+XBhGp2S7vUw1XxYlJOqXtQsMiWuc8dADMkh1wjw5yRfiNIAMfIvT7THlg4bUgtIil3y
gMsHxIhRDryUUiD3N9onRDaJfZx+WbR4k6XJZ/AEa3z79fuCiv4ojXvMM6XssombYrFUfQ/NlvdL
jnOawFc1mcs76vmyf3X8XwldMZRyO/mBIopixMx53iZKwah2J2Fas6aoQABVLfw1009C3rsSe4RI
zZGuYBu8SHVMCTSqlq4lBMNbBl24x3xSP/WcD8HKckOxAX7jQ4bVHQnoIfytNsS1tbkdk9pvGQLS
yLuayU1/p1axL3OHLhnSy6vHxbAqSZDB96C+9dQlqbYaM8Cke+c7j1CzmQ+xKH0KvZfL09myya7i
GTtbJNQOWE/aeOqM19dd8IgiI1nXelxOP8s47CJ5evLZnoUF5nST+bIl0ZhdwQvnOu5rXEi7asyt
xh17IuXuAscpBrhG5UWqVQpJjwN8LVLEFEkwI1GA+NmqVUOXMQ2YmDc38+ifcLMavg+6DGsKfmEC
QKMv27QG6M6L1i6PeXWrO9LJnWpZdS4/w3y2oZVsqxBEeRti86e0YQRmxe7zwbFw8YAGCZ72GqWT
DV42pI2sFKPcDEHPTITBfizKYnNtVbaIKvE+pK/wLNU3JHrywkAfeJ1ZiQ5hoPeip3mXYOFvmsCX
BlU+3QKz1NHGTp2yBYwewyGXxLYi6Qq1Lt2NU22V+LHsZrWuleN+A08qFQJP9TsSMosVG8NmuUCz
qVQ8L7vL3Ga1xiAyl4xhti2w2d2JhucTla793NWropAh9EAL+3frXkn6SBI6BNkg12giXpjNG1UH
sQ0sYCdZ37mK3WKPwMICulc4XR2OnUtjUiiKVdq+5ETR2ArIVXis0YHmoY8YFCk6hGXtfZVLKULX
ArPPNkF2TKIbyFdwKbHeymOVc0WrViRX/6TeCvu3mZm7VjdjQ72pyWngI5hQuaWbWo1HRwkb8WsN
O3TYPYwcCUXUrjgHAIk73KFvIh7+k0eAgg63id1TdvqzlBmaPfsJNZnHGdAaMKCH342AyhGrNY7P
jSBOwxoTQZnb3BJkG8YuwvbbyFGU9ktTX+cuyMczJ0sS7hFq9pJQIeyVmHvz09WklfLieLBUEf+S
vFRrsTQTmRq1rj50wEKwATwTJ8yi0Z/E3L97QOiwbLkWnkhJs2eW2YQgKyj1PnF7Gm0vt+IsZ1hD
IdhdNt+XbhuetzyT5fnCHDttvYVkaHTZLalqDefYMb3ykGa/6Mjfsho+ohXv8zu1+6lW9qRg0TzH
t2DtPYH90CAifi8NYktLdRMrU7RxxLnqIRZ9Ny9/lFj2oGih4CsNWRH8wVohhvF/DaSJH3T7IFHj
QCUMfo7T3NUgkwf7Ff54ROr7QMuW66aQppgldlXoGb/KiJVtEMg4G1ZSjabdppNW+rFiS7qMQ/Rh
rsps1/Wf2XpruWIhKiO7fBKJPlzBzSze+jHoDq8nQWSLwTPTiFHiZwxDHmIM0XB1Q9sUgpPzsKT6
B5/StEInVYfUDtrpYB1vJjTXWFd1z3uUiwW24y35m38H10q+LU/4/xKj+orAqgeYkSe75VFZV7rC
uqa6CncEA0kUsDlcZ3ePO11kgqFsmcQPHeTiVLgA+4fd5Otf07A2m0/lrjFit9/AorY3EdgGiEbB
mfixbimVNOvK9+wOtPWNPSj/D2pn6zGvkVBs5wLnKmKl0iP3Qmyv47G5Od8HJY9Cn+q7KPrerfKJ
blyTUB59ObTVgLi2osTZJtO3EsQo23Lzyc9PL68M38US0vDE3G6ooq8GkgEXOTjfGQudt8pgEKEV
tjA6eCJwoEf17f+wTAJdXOd8r94queXZJ9MVE4X+d50rGeL71SNIwyAE4x2e98579kICCUSXYDr7
UXMs7ZZPEhkJvX+Vh0RnXespaZK1Z4Ocn6gqMFrGPxp9GUGuJWmcloq99vaY3J7BaG4zAbA1o81B
pmAMFwl3lP3MFjp6J6LpjAdu1AN31sk0KeVzORZtUY/pyVDwXWjIAZ4aPmsaghKmtmrgLuoYoW87
V2WBEUIDWiOkBMsHmH0MeVMHDV4XS2Y312pHm3myHm/yi36UIjkxmwbyVwsKOle6/n8TUaKh2J49
UZw/naTJjx1dVcrtMXV6o/Ner13NT79WOU2VKHE5ctKE4bimxcAKBthOxNeskooGhXNUeS+pK49t
Yi3d3oXBmPHlKzuyGUFAY4ENIturspwyCxCcBV6W8I+yX8q6PweSmDg7HrPuDI068nuDKwQr8udh
H04HwYOBCspepyqLWukKO6ckbMSNCyRaUe+O4H2gh0YAe+qavSfMptSC4aO1hV+k/4Lv/xpUmAOD
TQsjpHplBcZHlMpU5QEi5HrU9T3BkiUHawVFTLugXorc5WJVOz2oEPhzlr418IwS6FwxwGEm6bef
EWqsQg5XAqr6Bl3wC7nwbGucmovqc3PDcgLk5zUdes26OyvO7xSc6DK23cew0UzQ6tDi0veDV3V3
14Qmu00b/PY5U5aowjiJBf9XKREuwaJMraQ1XLIiz7vaL5le8YdaXcYBUV6VZxdoc2AS/N/wmzDF
oDeY8VKc/BiU8MBvgwJqkkcB9uC9hxeMbwD9xhTZHecO9CQpqfA46nyZ9QqJxaZSgOsj4x1S+J79
17qkEimKpDyubImAhyUjENhDjQlFBESQ1kiTVWihrwpm16PdLiG6murLhQgEqW2T2/ZgSe3WO/L7
MXaarpwCkrcwvASIKMP14O5OCxz32RHca40/zNCI9gr2SBL8MYhQkM/AyjQIx+uuNzg3Rix/fkvW
Jmv3oQcW9A6I3wAT5BtYc2FVBedb/Q5VwwqNyNP0Aw6NLSRTR9wSe/b5lySslppnPtWrvwteaq+G
+KdjGTqoBsFJRCrreoNp5+SxkW7EflMvE39xDEOVaktEFFc8/eUKhBSnCGXuXemXqz/4xAsk1OeL
VCNEmoaSy+r3i/Qz+lV+IFTeYCj7EpMGEFQas1a2fjB8SGX/ZWf0EalKqBOW2VuTso3HeLUPPkeY
n773g5dWK1tYrPqZ0hTVUJ7urf84iaO+UnuLEZpLpKIE6Lq2JZVVUg/7JTSoE2eZ2eETI7PT4GJk
Chb1+4+mW+i5R4J0t7NVQyF3SizzSTu66Lg77SjPV53bC90QYAupODth1ZwbPYPoZLmrxPdQc8P2
8hp2PCm+RjW98/cFIb2emBABd4PCq3cpaZjKmcyIdQzW410v5E983c4+iCuX02lfV3zb79Za5ogR
cZpCzsIJ0LPFVd1D82rtRoatYbM5dgr95r72JsdvPHKkw75+YlCI0RdL0VbEijbh9AfxwHa/O5eR
7t97RnfpPu3Tp1tIR+/2ZUG3yyBIY8kNXHRstaeWUwtk2IimwUa6lhdOdyA4csff9AoLWZ/zJO6j
0u/xRWpue5IyiP7hDIczuhu7yIxezPOCTiib2RiJxT8ydcuAz9dc6lirgGUb5pQ7gTGOljr/Ffz4
UmPXI+CS6syICNilpVzH1tR80n8jnbLMthW4uBhsZfGfJRPnqhUcLqS/S1om10n5k+Jr2kPz/U77
JTRGRdidt2DdwtLysVaWFSBmL51X8+gSKqL50Y8qOn8k4JxFkFtw/rh6HofDergmfRsofoXvm0s0
e76U4X8xQFYNnWuH/LlpOhZ7ImMfHUgkE1oA1E187HD1/iSaoaSUwEAzkg0N+UxjJiqVigl6dbjM
mgRwgUADNqZ15IYStNfOZyiSPWxuSr3XeA7wKggJ7o2WS4ggyV0rsimbZjAyJh1BaQ8XqYDcHhwe
C+XJeIqlcV88KRlYOGsm8JHSt/YVvVp3fkNvwi4layLLbzwlFSzezdUGUMutw+QZOKltKM2LRkD1
P24GMMNWr5M/T8QPPyBwoiYThUFq4MyUtKLK32V/3MiOR5FaYHxAzyt8ZUCjqq2+FyFGmxXWP8gH
49g2UmpD+jlrWCZMXD0+96SEDkB0lvYvehhmDUDOZBDlYmbS1boUljSM/CKzjKdKR5TXbz8UqIbY
Eb6Th6O5f5AwKZ9p7STC7aIdlRn2zx17LHv1AR/FafZNTi1rjgR3po2oAAkZby4f5px/V//dkQ8T
62vnYSMN2hYjRLb/6vZs9+uAKy2Rn8IFJ9K81dT5VWz6BrnMV7EvEJjUFxix0AKs1Ox08J00IVmn
odrLlS5XGR1c96X4u4xK5UJ8nQVnxMPr2qCUTGT01YqOIhh8/bH5qNSfxWG4N7Fxo4B/HIDldeRD
A1HcE5sIqEfvvESzAoluYU4kdYNyJNKO5FLh+tw7XDIhClSrfGyQTiAEHql2niMEx4LQtWf+dI3t
Hnb18pn/2rclBZ8BvDkWFy9Z7tdtdw91bkmgfTbtONPHomIAg6CcxGm6zcPEt5XcJTgjKHN1j94f
OnQC86dHnsIdHWZNePsdObwbyLbbGArcAptbgUOw5FvUS0L0KieWbq+kFkpGfpFReMEP7fJTRU0E
YHwSVLvWQVomIyCgLxGAkZzCaqxEEk00ZgMdqWX8w5OvZychRI+mbXHojp58qGMlqpNCAyl8alfu
vI7AsJ+4LadFPQWidUCD4/UC4PR+5IIreB7MaLq9PQdxLU8jwTUJ4TralAFjG+Vcdqt68spJ+AAz
MLHEfCjiU4lLNrjX0otCm8rKmINr/0peDRN+qwVHyIEL7a7CUKLH9edTxrkedy8YL7+9gwg8Xnla
bygWoL3fZE7HvbTw1vWghECdrjj3cGbyOiESS95RGVXt2Q1CI/XkIkajuXPDG2+QP4/Vp1x/oPo8
0RJKcdZWFMGXjymXqLlBtONPhc21T1W1OFTSV7amOkRilUC5ZTJ6l82Zx9fW9WKru8amLeqGH2ut
K/FcsdnSMHW8SW1eGyta1i9mcPVpYuR8wzz5xRJt7iBjfO5XzXwIdKQtoMpPY6oURzKQUtPqd9HU
mz/7BeATuS7B15+uwXpGWwhPHMcm9yzMnZ9XvbOWkSUjRXLz1L207uJH+fU8j8plJvZzhLrhY0pR
ip2oPfwiOPa1JiLo5iqiZuxet7Tvzd0v0mxEDY9gFK5Y+U9GiMyr0imfpl+MCOGx4qX/NkqNSIuA
ByBKBaqwtGvoJcFuYksIJx6SrTkFu9+sCfIn5pMn63c6TiThDjt44tUGHlNfVjLN3CPSQQLUCkmg
WDu7NVry1UEnR6g+GrJJoqeEDQq1L6N2GjTvo4dLI5kmhgpqb6at9oFX5rtZAqBpmqBPvmRlfu3n
H+Qnj/EDcNv+JVDVqCNqLuiz9CyTRITG4gQzeleJ0wU9DKf6GFdoWkZwfWLuMWDK/jpuj0De7N9w
a9Vh0e7xK/aOzUxvIiNd1OvQpkfexkeP32q+/ujsNRkjC67yCHRj+mdNtv9+R/h8EQ4u/kCpY2GD
5XkdTEtc3YqZCF8Uz/P24YMOMz6aHVT3YNAcPT0R5806okFYQ4cGSqt+/ayyuUZ8bDuFXY99MbZE
u2giaoPuIXfVNcwbTAefrfoanEMe9NyfdeLqv6IlFBrm7OQvEeMl4dKqEdB9jad6zitt9tnuyny2
hllR2qM9E1vz/j/BOBw7mnsZpXNqUYgJJL1BRVPLVW7t2tA5et+KZFPW1Nh8xiauLrjkFx7kS9bb
IsbtCGttU5hGRqAvymdsIU67gY8T7wXDCcmvT05RlvniNEfQ4DcrDVWzliIs/AKA7ZNGF2eC84xu
9Jz/guDtkEH+srRn1uX82xF5h7mBqerMYV/tEy/ppgIC6T8iVCrTAHeuE7RcwNUYAW9EA6RpWW9y
1i2uDxRuz0eZYFFgBtzVJZf0txi5bnCgaCG6w8JpWj+gMOhsSMqAOl441TumWDz17e28YN9vTK+y
HMp+XOIwbObLZ1SLovEYWBcdvc1I9GqbxGH7gryfP0dfpVNtg2S7jJzKRD53VkLoDV5lsSCrfzhO
nUe+5JD9bmuQELMBacAutfDO0TWTOJ9h0iIntfoDo5MAZOssemuQpjCuhFlO9pymckaoquempY9T
v+uE3Iz/H0FvBH2fA7mz/pImSMd7zRx/pNoC1siLp/x9nQTWY+2f63cZTXv71JayhsswIWQpI5ia
H429OSEOhXhdNPUNBkT/+yg+XHurnYCLXzP2eQq4MQ59yev8tCgMCpSV2pk/8lZpiYvvhYU7NUIt
MnAonb9MxB04I7hLmECcj7s6vzVuNe0nhYihb+V8kSAVZTzcaWuM+Wz449krFRkg1GoywuwpznBk
w+6GYYmZHtV7/zeE1KOYD+1c7fgZU/EkFxZ9AK94bMAg+EKsBDZx7u9cLDHpioJ2OgN/knhVSjB2
LBWljrYxXu+Uee49iq8D1OYl7YfjGF7tfU9HIiU2yfDDWLDqDcDQQu1FXMKRbJoxTgV1DYx+smHw
vvamtzf8C0Pq2fszKmudE+Q9USd3mFKXeUCaK3DPptm/BPECnBk3iueSMxwMubUnZMW6SzqAmo7m
0ktdImZVTms9OqQP8yG7Rv+OMFN2MXIMv1egn7wfUgbdORVtx/qTfZxR3E7AzN+xVvQHHKLRMU8+
7bwfEaiWuYhgked4Z4BWII0Jeal+tGt1rk+24PGNeJJNtMg/Mvu5N3LgSNQrh6Nj5Whjxj3hojEj
vXzBsyaqorCzvVpJ8pSNDgQ8xEjKfNNKXbQJhag6ujcib88TZr/WjjrPgr2gGbyQeLvtIF/JZGS2
pkzzAR57epW8fCJ9FAswA8H6DO7OSI84YdwSK1Y1lFq1xQVW06lsvWG5jynmZkosfXrTFXtZz+Ny
Kl49J2cU2cIEoxXBXlDxZx7CIPuuZpLqJwTDFPH7z+TmdtjWTNjoUtanYgsdNBJyPpslax8ofkgt
2IUHYMuMG2mIFW/co3b7f1NMrnnqpyK17MRrW1jAuPoYOaFLrPCiwrbPU/2OZgwWAwOgEY8OrgZn
kude+KL+NdbOUDbRRskr+vQe+z/19rCWCt3baEykjBRa5zHjMGpepXinIxo6MBowNZNSYniSyJ4w
p3FOM/IzH8kSbyJt5alquRR62wt+9acWh1ZKWY1i65odEmeL9uJInUNjdtuzLaeseoDJ9xWmM3tm
yLLrg7z54/5HYj1Yb8o4zVg3GffrduZoxpFq1hnYvr0qRTPs+OVnArVOA5ANpEEamB4N1kjyMmuf
UlzWirImFcYRfPSNpS/8P5EmUTKDUbP4ECaBiu9wBewVLOadCdY94j+w23sjnCDJFqfkAMQ2d5xH
7lXETFCpjrM/bvrgZ0fWu0pYqwxLtDCV1lSUBV/C8P+1OlPHqJmETKWJtsEPnYkSfz10b3KASYz1
F39m7DXJFyQA5BHXfMTR8INZVHsTtjJZPlXOGbLKTP9vVZ5T36GhhM0+bszgjoqQUUQIbo3Dv6CM
SK9fxi1B2zT6EUW6V2c51oVwfeRq6oLrnAn9dcNx6KfID3NMfuQycIBmOkX8XGdNp8myjTyRRhz2
06WSHoBVVucRTFJfE7IQc0KB9kvvlxdpY+EZeWeXpNCaCijtB81mAJhHFQAOrm5dGuNiDY2/e7Uw
TuZ2Oh5pLbinElylgqJC92B/UCLOC8qJGSmQLYSvxOBUFWlwc/C8RiWeAjXkoO1GltjDRBb62kps
iW4KZ42BOpXBOHPWKeM/5gHDmhwJkaCj4mRToW4MoJfRhNhXGngByUoAcJ69WEqAWJWTik12WvPN
w2TNJoV741R9eSBlWkCWpD6Wk+aQCzAO7rmZWPdkIk2zjfjtAPkEnuNRoLaTCYE8dkxSLKkfYZur
lj9AhlOoasOgrPcp7Gz7ro3TPckeN9qUWdpPlzfuXCfWN9ZS8fpwBDDUnIpa53p2ciO4rKK53PQN
gEf1XWki3XtdkZjiZZKFsvA6E/D1WSIhi5N/ej3rD1z9KTh3phbI700LZ4FqiixHE2A1W1cUtsNF
sdjOlnDnb5f4l9Jf2+efmsEtLlbRj2bg+/o8XMFPR29KR5MGjV/cQIjft1nCqd1evfSfj4XNN13d
cY8keyUOvHq1JXCe6i5F7Ki1Zy4guZOzBo75kxQjQXiooeJhV1VZyNrwdW42p1UDeLwGagxj9tzH
47q59sAJP5ErXGkEuAsSILlONeUHkfHx3N43T+2wRHev0W19VOJ7DDRP6DtbVICJalC0OXv7sMtC
Vm2qnVKDI20LXjSbFIsVXRZb7R1OwePF+v035pH2alKKlO21Qtz6S8l+kbItG6cm0plO5HGFzl3V
k61ft4ZzrA5j0S09s6YJR0ifzoRoR4B52ZuNR1kQRFay24gQ0EO7UTI9Cw8ZLUVE0PGmSBCWeR2X
/vMYyWIm8caablDOeHVoSGkZw8MFYKtJCbUDDkfs/9r8UcTvcvLdQvjNsRE3Rd73H92tASqasjZJ
IwpAYG8RlojsJa/8X7A1Df758+oV/EEsypC5JCkUCPE4oVfVbqKyg33GJzTgYsFmEb7GO+h/376F
M3NhgPexVXPCTslByYN5j1wAAnePqKVZrCPFdcGV00LcE2EMg4Sq+sFE/PKslmo0mA8G/2IiOJ07
FQtZjKLiTgXxbVhjjhMpYW1bez4gYbg2CmXMgmxncazzKnxFgn8LnjEbs6FqUBMrXYl9F0TAuY17
+QSfAtoHMnieWMj1X2my7Q7vJJoWiCzeRoerm9tnKI1XPIqp7R5kewHrSbcFWwsCpbx6pfJlEdwN
vFbriRcdsUkHJZlXG10IsYMDssQ/Pg+7MblNwHaKqaT7vq97Yuc1k3cwm928lnBSNe0KT7gIGXAW
yMI9+Sq4XnPvbCHGs52IUV4jI8ImGPNt/Wjnp0NrBlQ/c60lXcwM+ydWNoudZSEFR4R+Omoss2VX
+CplEmrMlCGu6GRujSvdAAJ0eaF595YMF5mLbifm2YZwhvNqh0QcLW0zysQxeQ9TuYGIFEzO9NrA
jvRLorDbmZJhlQOkdneEyxSu7sxFszmrnNDWuSRTm0gG6G9DGhsdEYOBOcov4iP2EXhSauU+KIfg
kpwzr89G+LWDswmYBeANqcm2zo1caIBQMC5WmzvqTRYwJJMWpKWgN/m1OBjljHqlHOsWgGqDv27G
nqgW6q+RPy+ikOhxUCcuzBz+HqOOxIgB7mlSoh3NOWFk7FQdEfMSDP9OqcE5aXils5Y3deh5zA1H
OE+i1QmEdEugcWikBm8bqSPAeNCE5LZ8i1zPePUd6+i68tR2Q2/fnUVeO6N3uP7cgdJ66JkCSgBu
Ghref3Rqq33ZLwgFs1rebK52slYIVNE5/70XO4rXDAEcMlTvC2YwAt1sCD1A+gEQalJxv61NoNvf
Mvq7cHVqkCB1+oBFeSsVViiqExgtph2LkGXjFR6HI5g7K6kNiJqp8Mc5ZqiXXdhbOJ3qQcMfpOr9
8yJkfx6khrHC+K24EDV9mPaG3qk5Z/XTwFsUadt7z9XfnoZknfQSBuMHd1aSQyUJlllEq3tCELlX
cidsARVecRHX9loVpdupJdavqahDIjHigwH/yfiwDe5c3Tuisqn/NU/nqbemeH1x19MyI6jLGw+r
6+iESnhsZpUJzNAgGCcVC30V5MH0qp7c7sVpUnogxDZ3w1as2Q+ZaP//j2u9jVMyaEhKOwcS42IK
K34PakpM6/HB9H1vyTP1FWM/Xk6djhKy/3fj+KeKm8KudvXFmLVXNm+AYQBb9G15hexAtrB52SgN
5224r6Gvyu2+cjZR95WmSxwVhNffoQ+w//K04GKu3s3oYsoSnZiDc7w9PPZxPKdUFE1dfYMFiSSB
yNUFyzmEX7L8l8/XyVRP9pGxQ1dlIjgpLduA/Sy+ALgLrVlazYlpArVjriRpAQ2IREiQk2JTrkOb
QuNCTUVBUW5Ihu6DUhZqYGam0ZfPgv9dQsgSZ/R3v0H/ORTR0QjhyPXqGPCCqheW7wrGVstnfcmv
jmya2qIuj59l6DfN7EzzISTOLQpDapHgCZ86c8wQ8xbQgw7cRukyBl8u3HCjPxG5pmiYq8xmg3nh
YV83Dd95PzFHCyHjZcGlvXWJL0DUFHgwHjzkcXb9QlQ+3PfiemCrboYFjjStzGJgJp6BE17Qa+nw
/ydO63QDPIsp0E+Tpi3Z7/KAkyr4q03pt2D9bEfqnNMupnKSv6xt28njiLlWNO8VkwaY7v7AffU+
uGxWyEenjLLmNNYqqF6Qhzuo4mWN50KfwMN4/NELPHHcpIcq3rfOmkqQVQC5GMHIMcexJQpWQu0v
zcDhIHbRRvsFNTU7ZKkfvrNTxye1ez3O42uNtEavD5ICQIq7uvuoJzcPshTPnbg746KkTaFTqJJB
xmosX+oLPNmhl636fwq+NjlOv7uSYMZe6RjmtqKPjT+Gc5lZuilFXQB9+Kz8Z/5SMtnpQ8m24fCl
JWGKcZ1Ynwje+wzrdiv3zsHjKY9jo84TojEhfX/N0gtWIefbNF2jV5MdT2G+wtxY7jOR3/+tYf7j
NVJB4+n5KYKK9urTEKD3gHoixTyn4V265uJ71hpbqxvjiBAlbI89k3HvxlgJwydvgKqFwFslr/S3
h/24OTGpnuhzfnq5mzhJiUvWR/9/ZSifcGI7DUHn2sre+SO2KcYMiZtT9WxpPXvgzVFNjrDL1NHP
g4Xv3L5EnEvZi/ojWNmS6CDBArbfq8/HejB+Sa0HQp2L+A/fmCaKJpFQR6wpqzEVfq6oC9fuvYDP
v0p1mq40dG1dmJNBFgwPGAohUhHnQrx0owGMqLbYfRs58i+TmOzfC4aAxuJGaY4KlACo+5NRaNXz
PTSPgYgQuCkqiJHfD5yGTmebwyqqzlLOG91V/sHPXxkaW0kvREO/e0RYFOAp7DaCdEDMHDIHPkzq
cPwhP9FlEa4r4eEfC33EDG1vM2nNTJKlZo0vH8wnCwDlOP1mRubkiSy528EXjVW6oVnutU8KvZAP
FfN1U5VOcyFdTScz1I+OTpoOa0FsWz18526Wc0vmU3n3OqA21paOMNoBY1pa/6SUqD/6CAMXhkWS
jR6HA6khO1s4oAN4u0pqoIYIAHohxBx1RdhJOxSXpG+ag6IN1UTgOfceKEmEqwab4OJD/kNdPaJF
AI8oL/biI64IuyEIqp96m+0RI9D203A6Ocac5bDVbjWvZgc0dIn+SQO9wp1eL7L3Ma04qktnWOw4
/J5CKQGW2zxe+UyxFvrXyqO7sJ/ItvmaIetOOZb4C9HkTTGbDXtQa8eSWGV7EurYdQ99G3d6eEBy
cZeLihXL6R5MNYDXOm5AqvaI1+hAAsoSY1rQsFJmmVTRMSEppd+jSxxfwbbL/8zWNEJT5q3hbsmq
QolgMqAN0cPuJfv0GaIYlCtEoB7/BNfKSSlsFqspkHTNFfOfVseUxirq+D99CXfvr5blzw5DxXOZ
howboa/lxggoBxbausxdBRx03JepenYqCawtaVCsete7jYW9SmDm4n+4J+2/QfCegcRr+JV9aXlZ
7gbapn5N+zdXgf5pfQzUnXMym3E189TBEsGVqGgrx3cS78llsctfy1X7zTXZoDhU9QE0KGR0ZnBY
YLPG2JXJRJpcLN0HesXXrPuWje70J34HtpiaMLnPNHoqaivRAhYgZ5IsLgjHvie0b1uKCLVxEDQG
6jvsAvM8fvo7u8oX0CimedSaKoDtIbj401P5+VGHWM9j5/oigXSuNKdmRwCjzrd2DS3Aium5ebRZ
ajNkkiAOYT9exesVzkdr6QCpApU3vEJFiXw6c0ER6FhoqQk8+fI0g9BcJbybfg6drnL0JMpn4hw5
KnnwSXqiriX7kEcFS6cBB9pFiPwIovyKS1shicuanRNaFSx+DKK504tzHSvPjPj9HSvtrobzPC35
qOAYJbD/Ke5S94sxmeydUqgnSgqaQrX+oyurFi5zBIw0pFuqzgGY0lKszhXJLVSmWUCeWc+vD3tm
fgUEWl5PwyuDLcf7DMq1wmGRMb8dyURavF4k+WA+EsljN17sMd2debvp/eDAYNAbnCPKRcPb065+
loERcwQK7ZdARcAgSwoDIFUXAzORdYFkYPVdWx2ImFlL8/Ex3TYTSkG9q24XABXr5mEo/boJG5RZ
ylMyPsrOuhQNz3nKR8w3x9Gt7Yd2oKZG1d556R50LjVx8h46eAIgFyH68jkhYe8J8/ElM+RHWh4Q
3L66CpRwCD6G0WwUK3/5DVYhTnQ1FtwUdzTGhJXr7YxR06AP/iZA1k6FgGoURZ+dOSgkBB2nXAGF
TpN5KlaawOSc1J4GNkq5jQKgzzrrM6FOtMlVwzJxYodszGcmT2CPXO9uJh6JMQ6vd4dnz5oZbBQV
EbOiY9nU56gkaPWe4/OymGzE+RjlWodBQTYqUhBs8BCbBGHRtVhTvfnXTlCs6yEk+0a/9Aal4s2K
SAT8LQmc7zYGcSyvci619nyNp+HXPtxvtWpsdJkxY2sapX1+aw6GvFtg2PQaF7nXBQzIIIRvrumF
WRf8LPyCcZSmz9GbyqOddzMSJNvKnueI6jRTYrv7jLsaFjYlMZAydiC7InWE2pnVhs7FJ7lI/GTh
eS0JUGij0RtBg7WbkjNFJOA56lf9b+sAiYDpLfQ59lJJZyguC/paxB+MBYxNfRYb8GYuqA/iDLEL
BGC33/KO5aGr6hE5SAh5kFKdPKjh/0TEmwCTmeSaUum/SLFoCpqMTUAAnfFQfCwIgvTx3VEsIFXG
wHTbpj2h8yRk/WxZSJMQuJ2ActVNvKE0YkvnbRAZXPvEEl5W9bTgsFIXWkSLJu3h6em1gx3hWJ1l
7tB7aslovK5BHxmLoJesTfpZkK4jEn54+DhFORfQc/QpICwEj4FGJvXquxpWPZC5dPNFi1aruinN
BxFkh1JB7iawsTTgsylq0Pqo9blR5rvkA1Tbzx7oX/2/9QnliwCZcfX7G4lkrIvlMNgUkvpXMD6I
+mDwfz/5pXZQmF7CmeojAfG2PDBIfpdv01IM5ZssQ75PwMBDcTC0kil/hsn7XApydpIQ2YXkOAwW
iMRjZPyEBsCXBBns+boaAskdjVyY0/ivo3o4EIjRKa+c9mI6H3OHimhEydxUndAxSZV5R3VlIe+q
7CX9dbcP4qJU4A0LOHia9SebC8mzr6qBZzyEV+W/8u6CfV7uYLrecF+XFfAMROBZV93ajBoF7bOS
7/cPVraqvX726BBr41eggPv4ktJEKHBg+/flYT3P/0nO0awnAnaGEuWca46R/tBVHLQUQWAbEjJf
k/tuZKDMkZlysi4PvDvZWgSuPaKC19jQghtmhEC7tVgywwl1vRIpZnPQXxVHb46mkmtP8T7Pi4qt
prrTKCQ4McKyVMZ1y3g6aJ8v9V3ZZXLXKF7lCYNUvRb+DnL0neFEsusfvqjubZdW6gzwCo4jZrEe
kv0nL2to7L4IBFlri5K5IIhXOiHNDgZIRU4JQTAcdEo2Q4THaNf/ld7525wOeXkQyZqhlyPxNrdc
LV0aCznEFPV+bw2GFK6+1CZPdDh7XSSGcVh0ruOpx/yTsRRKFy7ekxdWRrkvpWE/29pRvce1r8D+
DFQI9ZZGUGC5kuil/11PBz1bf/FlPmLpY7OWfUxXMCZPSLmQf63WCO5WLNN3EWLZGIApTzXmqx74
XE/iWiMHiNgsTfIWMMnB0cJaU9n/ZYMdn41nf9TZyxH68JigCFq2Ew0Y1ilopA3yU80kbfdlvNGG
RsPiUEq6CsRTI8lXIdAPa0JWNt916wnr6LAOb+1kn3QW+5+ZGBJFAcMF9ZSY9EDoO9GovT4Mb6/F
OpTiAqVpjzSzXS8GjTnkl/ZiwpHALV7DI8RCT8p0RfXpGkLyOIq2YzvgpuBJ6uEFFXlGfb7lnkn5
XMkK5y36AP5Q9IA+W7gVYeBeuks9pfV6Ua2aAWzxJtpLazkVTzxVk3TyGiyEOeEt6cu0sgKW6LUb
KEI9ohzR5KHkE3FuV/lhfPAUDd3MrF6MZPzDJGu7j2Uc2zc9hPvZ5xiOvkuDSeYKcbJhkVGPm7BQ
+SHWY39Z//7UKD2EeImvz6PxLMwhIGs/Wn3DIUiqIoQJxBQOGsJRkEX1AsJtESFm4TZSE+5rLZT7
OYQuN5NHsEyhFu5YZX1I84+6fhIy6TJ+cpLIzCa91PSuQFkbg82qZ4qhtcts0T2ctauZDtQCvOaw
yC7B9zDHe7ChaI4+ilowp//O+54nbepETXiYzmOPW4NQfWQIZNXKSUN1La35ZT2qqRFozCgVa3dB
XEUGgaqmRrlr58lB1E5AFl6EI1ikpK2LhV1DukxFvp+M7v/hHTA2APKLowjgq3xpvr9+mCPtYN1B
4AG1MVkp3GExqfp8W2YnOm73VR34P12tVW1U3O2eGfxidiz5WboTGRe4NOEMINaZ1Q1Egyp+IXtm
bubUvgD777qtBKPJDHf74btGCKcSHb8w+LYlZOjvEUKNhw+H2igd77+oeY91VG9T6tz0qmAspis1
nC0+BqA0vkiR755vJKmgGK8UyhQftvV6oJc5kkwSYFoOHhL1/UlbLkI96O1/6HbcZ+aLCpQ0X1G/
k8kTs9wwb4m54ErQliwQ9cvBWYWNh/2iD6O3XfCT8KwjoKSd+EcZlKFNA0NK4U/VndNnmDSX4OLp
a0VOakdkgCk5iuRu8ok9PWnwLwLFiUpG44fcSpnI3uI0JKUxXXwgiDMy34O8G6I+CtgK6XYXs3fr
3hfQ4IME0IeHH3TBAxutQkjciMeTE9yVK8idi+9zYmenhZmg0ZO55z88ILRKZ181eVoZcz+Uo3Pj
twcLffdPelQHURF1JEGznFtAllHyF6eSfj1E0IEnFCa/lo8szlkWGCpiYSf75gP5Z0NQlyhFVmEY
PlQ6w4fQY+uXj9zB9EfOMdJEKSGo7/GktI8cTTJOLs+E1KJWoytGLjEYwbmeC4NgITfEyyc+1gaN
4RwjA+rYcAemsFH8gwU3M0YaZ0cxZbi5Qj3NkfC5rPjWA6iwzOfGoxnpCl0eunkSY8vNP7AjWDDi
ZBEUCVWaBN8Jx50waOU+eZPeYgVIZTAygwGQhOfWu40rVk5xWut7iumViiyjwlvfJalEdfboq471
KuAvQRL+Hi1rP+Z9Xvrj1FJFqjeGZNX0x5KEBIJoXdK4KEz5zx70i50ozS4c3C5Vv3cVNkdDPVHB
KgjKK8ijHq0pZCnr68rWCklxtlqCCxO0NTeUvB2+aDFnrF0JEtOKUUwM8jU0SWbPeB08G8kGMmZX
iTLazVSejVuUJCQgc5Es+lMhX6NU7ZGL0KD4AtFGwQF9I1ed04eK1/miy2guk/aX+cd4RdMSSarX
lSoB3hF8nwIratffg2DGlqqluBrRPwfoOb1+4EKdVg+F7v5WSHUfcN8O+LaEk9Nz7yVJIbNAOk7Q
oo6r7C9zr97XzbgPBVm31OonlN9LHhAavYhAQAvvM4VV+Mmu2Wp5bFgzCypfvu2B8VaK4gTlB216
CdCm3gS4VjLdAWpKHTRAyUHdSuVGKiKGbdEMnnV3YENo3ZrHdMwq6MN5ZoCnlmvSR+kZY9j46mhf
br+/m2vQeTDMMDBCd/1gCQcAdht7NwB0aFNARiCtxHocAFl5RvXs7rEgZnG84g2lZ58IlHqRgIa+
g/MQNWvs+uJoCqGLC6ga1z/Zu1rjJJ4o5te6/1iZCPx+ks9DZQg1rksp9d38xFgFBKJCBUInylWP
o8q0vOjaV/m/I5IZ1950eeUVISIGEdN9NWJ2uvgd2tAFc5Q6yAUioAUXoJzQDbCNt+u+BbdWND0f
GSenb2QB3S++EsEfoIzWq/KV/dgcRlyWGoEJ0+LF/jNzv9lF11w4+1QvnkRGkpbLeRzcf1KWP6uN
RnhYSpaRziDLtBks/nbWMCvgxAmsJ6lEzTEORgfxJsZmx/cbh6YnATgvtw5PWSu78NmRR43mYsxh
Ls+7jOmomXGS9gwwN4CesPh8ByP+SttrvUGwYSMg0Z3uzEQsDaCxSwDcoOo4dRv7hqoyJmLhIXB+
++PcEN2zcRRffUKioF7i1gXBLuZD22DrP8akJZWFDVM7et6mDUgz1hpUXvgfnVqb8nw7172ktI5d
x0ZkEzFy8LnmicBkZwbfpgrrIMc72iA7BdqkADCD+eZgwPnQ04oSBnHJsprkANqwvvvdROieU/sx
snLkiojbpOXsf696uTj4t2m2Wshi/XQTqC+XIaB3ZTCiiflWkzM/1BRjLAxBIkEhQZxAvwx6zMp5
GUn1dFGVhH/QzxiI16vrtGy0lPHE3Ic3+jobH+gK3yLdieQrjuCldZ8Shhzfuc9yBP4Hn7IIjG1H
05pRQJi4gBwBwVw0zVxlU2ZAfrPwu2DIY2x9S+MPE7YXedb+0riRFSHVcPeCb4/oYYISedeAwsVC
SuGrWs+q441nnZhyYvzB3eUzXohIIAt1zfNa3p5RbpkvdQ40NGGJopDIQnMhxZKLPMPUE+9Gm1SY
CpOab/FS3YpYOrshiq8EtSR/YGCM8YVp6Gfxv0t1TdMlpzIM3umf+UEylqMuLzqnNYB95r86OJQS
4NkSShn+KD0dJqVNOa0mXwxCTIN91Hrqs9qJOTbkvtd634vpMLi/Vdbaa88Ph3hM/SxU7nUH8Z6n
rSqrRAbXRBDQo1ynFstX+5w1LRsM5Zaz0X+ybkdquWsIcAeVjAyntlmR56A8iEr1t0vfyqO4k7Co
9ZmDd3zX4paCefhfIILzvQD51OmQCzX1ECCe0Zi9CXNhm+Du73WgxJyywbtB2enPvsOt+sB5Nz3w
fHO+nY+oED/4oq2QLsxw5heLwofgHsbzPzL8nwgHmf3vKZ4WOtn85wZo7h3xRGto6T2t/9GSpmH1
geNX3aghYxH30+6c2srdnopbCuaXz82iwhIdv3j0AcpV8WmgwCqo5s9JHvbg0KZzOYgVBa0ISOAh
Ysa7v8fE5HpqAm3tlGVSpUeV8pBwWgOS39czB17h4PJWLYa7tyhbxAN0iNNFKlku3gqz2EEiyReV
J41m02FOi+YZHCRAo1+yPW/+QXgnrq5gyqM460CJp4bgTrKnGY4onOIUm/w7iYJeMcAQ2cq4NjB4
FekrGOgQM1kqxTbwQ6Rs69OimBvPoXed3Q2opzSTcxQ6dt54YbQgMoc/OyDpFJHEUlCtvl4xYnKy
HtsUJ0MHcaI0JDBv/I/rhq61dpC1ArFRTrvj4Yzb1Z9j8gBrlLozHuIOpJsHOrGhieBR4h3XSD4X
Y/Q+8eZYO/RlcjafSVB9ALjy8Gp44z24sVrGcI+c6oWe3Nu/TS9K1zitHccgK4GB4UhiuWCsQtIj
kj90EiQS27ZFxGqOtCWI6WIMIpzk7cb1f7NFlPbivYm8xZOYcN5A9RDUzrgiWfg7/hYkzR5672Ju
YM5GHy1USnmvqbzI/zzAtZF4ZFW/GREXvPuP2+uMwiHQtdRAMjPG0QSefVeF/eb7cjJrcfCd8agp
fv0UF967At0tMmjdVyesOzxsfpBeQ/laRfMzLHJSlZEYxryJV+NHJpxUsSs9SFxpa2UlNM8a3ubP
phB6JPjnwbUyoJIbi+0QK8xmS/IRTBQ4HdPR2G7RdOQyyaLlnvEfBA8/mXpKGre9jQ+qoCdNocwj
EIRvE5UpJr/lY27h1CgGplkRGSpbaqvLKXozSBpWoR3jnmtMIp2ai7ClfZHuNKrgZmK7d2Rl14zU
mpbzBR2zqp0AzSnw+4eqNhgsUHDARXcRd8/1XlSv2drECtSDoC0xydXb++eLGNZ7DSEul1G4BC7z
hDsl4ZM3pb0kQLSD3izxHFYq0eeeuvGywDIBHJFTRG8y0hewATF4zfdCaZTj7kEtO6XC3AksXKUE
U2RlUz1kwH8Pzr+U9/7lqKKg1h6A43p3k07bVYvndX0DmVYh9jxhsS4xn5R+LT6R8zRzzuYrBiU2
ahSQQ3F52NT+nK8nxz677v23tzoGf86S4G/dqAHRNbD2XfZ2B2VnpmCueO4zXWLPCS1O3ChIUgFp
LVUpblnNw2AbuUy3g6dlzHIsvhNvJ4ukFChWIzizaeDhaNLWScxScK8aDWIJPOe0Fxq23p7EN/lb
d+SnrYbb4Yl2WLv7qZk7WIEGe4zjj+4Td/8Cfku4m+jY3W7Q31Az33SbVkIyH7+TR5L7H0DpT5pU
QfgQM533R3oW3xNBIgFsSsd9WTJ/2Db3w9BzE3znVfnsDjAagtpp71HgbK2Fwe9ypTS5tQooOhAo
oMVttevPXiYXtsUEMWB4n1JJ425rQTtHpYlv4c7Ec0WRH+2xkRpCaA5kZAeYJPTZf2AhXdVcYDF6
zTc2sr8TteJkUbF/c9C67TSHp4XcG286LQC1ylp0f1ThMfZ3j3d2TRnZNrw6cUPW4K6eFTXKzI0/
PQDePw25Dk5oKlhQ6j9mRxSW4AHmlc7u2xNXit35y3HXnk2l4G+vzTLUWonEOorDHJQcdE6OBuyC
rviEz7YA3TzRooBn6IX+cWjsqhDFIxURRKlXb8fiIM2u9hTWA3JiTsRShB8Z3FjKktugCQ2To0qj
5DCcz2sYauXSfYl8qmEJsuIxmC4sv1zVbe5gR8iY1k+5u4V5UlrATHeRRvkCBw4FliadBWNaZ23K
s28qYTna5CqmlUvTnrlLNz1jlCWTc9/1EptDXbTCOB5YEbVzgQosgzoalnHUH+eakwjRYqUzElXQ
dzloDu0nqe3sDrNH02zEZ7Q82lvdrRHT04stJubYFjN7kzg44OS4xBcbnvMEGr7JqXHcJtLbDmGC
SouA/lQ68k3L13dxTQGDHfviQ0QmxcEtv1dW6xrxuhPj6ATnLqWtXtfInzh3rKuYzHRZgXnSdyEw
ems6VCUFq/asZ1KAqG+eXbo5/T7B0jU51COHSIvD1pLzYASPR3Y1ofMj9DSRi/1TzlVuq8IOGq7P
+yqAv4iWw0Gpqw2kB5IA0den9HlvNSZnt7iN0T3HpyxeSRWiLusEE3OoNPqsrzvbMYnHmhMjYFah
zEHQt7ZxN7Q6Q+dezB110J7Jcge9umJQL2i6/0aW76Oo7MnlKNfG9TH+h8n+q6IKhTT7sYl0v9If
Wmpd+DypKCWtFnOBuwbdEmZw8J5ipM4JSq7oTDTdoIbMEQgPJrXs8dV9LlcyxRRtQEpNFMPu/0G5
75fZq5bnEhGSzVC1tW8cheEXuiY0mNQq7cnZd5ENyTQEbznXYR2/o7ujtGD2T95X/eBuxoXqy+3Z
HFdoYsCJq9fFxPqqmDie82yxoDp2vyOPjBpIEUpzZV44xF0KYbdB9XJZutWmO9E7WG/6SPQoJc4j
kdinIMeOGyQ4zRAw9E0Ajh0U4xnoR4Vd1Tzlv/c+LRtQNHRm3Ry6s67znhheqnloU957A25vLcSB
4bfPakXOjjGjv14PVIpwl1KK/nlvUvD4U4Q5fX3woVO6IuFgtNm+d3VhIjICZZ/Ucc2O3JhexIwB
GuuxRLzjcYKvydQ92JwtVOGPESO4CIquKZSsKBtMGxDM6GlihrJnNUveD+vjYs+YdH0iZRmr/Yj1
ghGfCmYwza38YCK07+JZBAVuLAM1Xn0WPn2hBjrQ/hkBwd8PulVpa12VaxOhcPHZrRktf/akIgQr
9Lfp2mADj2fJ3z2PfjuvgS+x8DFTEkivwo2KVqanLKCEP5L0pFOxh3xI2CSayhWDpGv9q9fCbpcY
aF68LrfcBlQQ/IBNrtCRHbewsusoOX0APp0OPLhyNZ+kE0iCofGOkmfvX6x3mxNQp01k7lzp2HU3
K7/M+vLTFPfZ4U4eOGsGCyk5MVa+EKCHCtn9E+jEzQDTk4TxEbrGIyop6qqkJT1LzGcxowJJlFkB
jH4uzAif0WpKdUJSbgClZ/t++NxWuISuwTve2WM6BlgIztHO4yuy9+nkEeKk9SFqLXGqnrl0+Q65
IcvCMjtjqjUk/tAoc3R1LFl8C9gH4PahSE/cYSWHUiMm+kbUEmfNzcaWO4pPIUGUF0QrbHljsSfE
shGlvEyaOF7164Pv7oGX/EskgOQfbZmjnveaJ11CcNGjV8weXd1NnN89Mj5iyxlzbW3SNgeCjUg5
40ITxrPYSYPkDBXBs+rjE9XhN4dBOLGcVeWveod26mOcS+HVPoigyLklmSvvXhSey3GS1uEr2wXe
WHtpTR6b/apSZVOZ6A1smDPWgWvAfcRUWtCJdDQU8QnazZ8GFzfHSOzWWBh+Ep41ifr0qIKFCOBf
1e3JD9afrZbmCIvrbiuagL/57z+lFS8aqmdHqDm98iwEI6eMqgCvWqkPUEB+i4iYvpOAR4y5wYEs
nfnAVgIDbDEHMi+De/zov6tJdu+A+D8RqA8eaAPCkWsrN7KG+Cwg/TOfk7POjX9YmYZP7pgKYqeE
zpNKlTErkU7NkzZVA1dAovnhFedcHdBkqBNxFroRwdJgG1e5RTcoeEFcl7WRNTEFu4e7uSIjWCvf
rb60Udgrs4lhuvc+NYQok4IIhMGMB2mmBm1vSl3jL+AyKQ6ARC06+zCHAi4vDV+mG1yRK/xeB1JC
4hxhi6JNmEK4ladFAgXRmXkn06xtN7SxxEK8EwR6qOElvwMc8go6b5xJ0Ry6olG/W7lAiYasqY3O
DpsQRpPN/Wyhd6mbh9tc1caj2BRUvZ2Xeg40PxLgYudnOvBU8P9mKruTJ9WhvcyZIUBfk3wqZaPs
fVhtwL5xEPi/u3NojrqOwxnAoURequTAhOc6jBSl1ZDYMFTUqI7LS007kLP4/26HUmI7wUk+HgLa
j5SZDyQk8mOJt9PiGc8EG6rTGc+krrRPvEC1cJ6rwBZIbQc56kU5tNKppqvFOSIlLjRLCR478x7u
ZdEsfQt8xwBCgAbz2EoD14eEn7A5+Hwl3tJqi/7fCXrUqV0VY1Hg3qpgLUG8SeibmVpMbImWIqSs
GhaYl6Dxc8J+0fJRGdKemEdSbkU2bro+ftEZnBdwWsDRjRFNifzWFrHf5bCYoGR50ZiSY62d+qr5
tCgxncM/RPw9g9QeJJH0NFQ7aby1cBKY3vpXvS2P0Uj41Hhb8eJXFhv00XSae28nZfYUxCk0Z9lb
QVj+LpBqlitl7EvvBRJG5utjBthk76mGShg6g2DZXg8qyzVMELWHZ9/y54hkMwEd51Qjt23M4SfV
R9Vcc3Gx7gsrneEoaraJO6lIz9ehssKT93+DLaDDelGUagb5gKBJL1ZpL9aJksrbwhs7eNj/tq64
zNeBP1FEUK8Mo4dDzOw7bTTHqGblFLZEBbORGtTu2Af0gejmMVjUN6yIrSaiJIRjYbK6kSBImMJu
HiENwTdV1Cw6lY60XRXPoiomIBkuDCBitox/Ph+qrk/bwGt4P4P7JvdR7EAANksrJJSUoclcJl4m
r3FTMzY7C5bRcSzHwO5kBGmLJaZxYMpKGm0ungPxk0kMk3II4MRwn2jkx9qBHb7Z5tFApqIdpe1F
PqAnnJyikbi3Sw8vHQ+SzKrihKcjOg4qfhnfrVJWI6ITP0c4CG2y6Y8UmOwx5F3CGWvOrT+GoK4T
DtXmtg+HXkWN2egZ854D9xcB5NP7us3FkFfx140W6nw2x0ah7dqI4VAmmsn3T4cMDYK0EElf4ZbR
j5UrNklP4VcN8+XbR9Vs1yMjP5q7fLbt5ncttIIV3KcT082TVcQJYKOZmjrHSs50Q6QREOS6FR0N
BQ7J0fFTZycuVofvicNaAVxOuf+WG4gCJASl+i+qd3Tc7hPxbFaPIFQwdENnl0knYKHrGs1SHoLO
sLAxbX0g6tzqlbI+a+IsQqXomj1tGAhdLhWf32KZAuceoxtBYbnx2TU2K1XnPoEv6n0OVzUx9l07
U1J3HjpI7hMno5qUXxEmq/67uUCTA9WiuKu+S5rTxJksOasEJjeZMCrMisC9Ih6JW+nmiBnwo7Mn
2GZQmBN7c9h6n2kkvqh5UxsHqW+FFXV6v5Wmt+zIUU1WGQQwlBfBY3zLNbPPLhgU3hafJyjNoJHI
VdDrVudPeRoz20NT8leFZ2WEjo4qyzHduO0jjb5c0kQja2cB3Ed/GJeChoEoqV+2JGzYrqZdYO9P
3smd/hr7MnuKoNzlKJxpRpUByNTpYwg/I8oC+vvZSA7jLTVwAQ1YGCTP8iv+yWPZy+hj7VozZ9vg
yZ9jo/nKiJj4UuMLeax3/SvfKBdLQlcHITYz179vIbfXSCbgyx1DpSXi22urpWsLvgbaOW8pJwMw
7bW3B+kJIlbzVFuv67yCf027mjQ/r6zYJz6Utnr1HMERZqdoHsQbXUVCvBBBoEVOt71KveeKb6hT
s7PSmSQ+1M9Xovbnr0fnBwweFRe1VvWwB19IPRIS5bCAMGgaUzUCLJghyVPDPLMJDXdmOQHsCF3D
nAldpSm/XPkn6D03++x6UIFteuTNdKkfQPsdZkEZpTGUoqOvMkdKraxGWGliuLKC2XXMAq/YlJgd
JzB22EF4E8xuK7rAwoIos2bzhDMqUU4wx3mHKbD+hVinGaWYyqGOlTVJOj28oj4o4oFxP1SeS1TI
Ncan0tgA3eJFdzdWYKGf6aWGAPEQtPZN6hgcmtQwAmQRh0uXawymzESPqwcqAzN7AE2I3RhAgacC
DX2H5mKgdNPy7uJxGv4M/JDZlhcYMTtux7o23Wu1j9rIDGGJgzzZSPqJSscsb2JsF2PUGm78DHMi
v2xLmhUSYSIoB+8KbsTCSDK5aIG2OY2IzqSfFl6HKKtLLKOqahioI/C4Ru1564bJqKtDG+R2trcy
8RvNFucy12Z+ENtwH8XO5kB2bCWkyGFFnTe1J2wcfxDEb75WgsF6grH/h1wIm2XQTmfz02P4lgXe
l5GXr64zEcc+e1nGv1veODNIOhDDAyyUzGxlj1Dpl4JXap2n7BL6A35IB1c7PrffbuSw2cyz7jHa
Nptk/Aw1XK67L4UNBZtJuF0yvZM58cauwVc1S0DJFu88u+hr1OGAGdelw2YWmiHQ/uc/Fg6RhOPs
nE9jgzTkxI/mpjz4Dq3UGsocKjcS2Ybt22j3mwEroBe/giug5fV2gERJVcvWxFiKOJ3qYnJBJTFY
vOeWd3BaLzHt8rDHh1JDxt0KWX2WvlLYPgC0RIDIxqDJ4+GzPJ/GVt6doZFdEJ8TI+3XQlWl0XfV
RgDkO4pY+GZoBXnJXp9L5IV2Tzv04TO3hKPfxY0occ2nseE18nY9hTMdMN9e2Cx4so1CLsRill66
wPBcMNrWvmZVs3e6eYY+ceR2Oi4gmnmuFPFI1KbvJVh3nrm1NHiv6aF5IJkvYKYUjjOw2azbUCA8
ucn2Rl5DlAJyvhJpUKG8xTLNjwASstJk4L8kKTtVbcWKeOgTdX0LrE4YZXDoSXupndjvwPeXW9bc
HmfaAb6xmE21z6v62ZjmjGv3XjRJBaTTZ/dRblPvrXT46xSIaFGTr5PEap6RDVAYbU6NgK4/vZq7
rudB+ZC6Yfcqe3jbHhUfNszYYEa7arAScEnJJzGON8QQy8VEQtN/tbtya7QGzZx5BwS6QmjCm8Ce
nAclyIfgAdcACu9QgqL1KDNOVxATbHW/gHpKPeDOHohBlF4VrexV3BUGC2mqxaukwxWImVGHMGbS
kbiD2Fm7hXELGTESDWS8NKSB0O5eGiYq9vvCHQ4+aMMIvhQYtCejiqt9k0F1C4yiVVBoyqjkOzqU
m2d42tjEwEOaDZdh3TR2SEyWwpB7cmInTSIpXkeE3v7S5It60xPgoExyISKyIAfOLI0+oFTcl0vc
kaTWTsXuNnPqv4z7p0qPmD/CiOS4nye4M6oNhqXmODPYCgcdC/STzQVOr3fxtOdxu05wkDgqqmdO
lBVAXnNY+6CDHzyUx9GtCXzq9bUkb4NXrD0IBkjvXjZkwmReO9XoHEvKWmJpGWi/jyKUC+gyf1en
ZYwlYd7GTrNPNCc4SV4z1CWzSyfSwXaHyCWISLlotKKiFH5OXEP2H0KFF4wouQcXAPqBFjtTfVbi
g7l+l9IO/QirNdAY1re05qE1dyJ4j4+mRyxQIqDqQ/FXqegm5SG/YaP3JSoh3PNKwfXmjwmSO619
HjV8fMPI7sUZ1N5tWFvcBLeskQV8ebpOd3FYE2wcWK2jdjGMe8n3zwhvhuAEtdmGEij8CyfhS3tI
+xcfi6kGLTTX+Ih12UDe59rQaggBIPIW4XbiJkrfupfo3naAn2X8RDSw0KFcnG22Ti/wl9QysvPt
dcXv1K0hdH2F6Yw8pFEAegMHECpOWoki2YGh2F/9CFVlVAZyhxWl2MT5h0sFFC+OxMDrVgJVznnU
y2qnonY5ohT262Ee852E60ntT0mCjJQ6eaweMJhG3PM81XTv1kR3coEfxyMwC5eY0VAupfVpJnTj
1mU1fgMeBmS0b8wdYAZm+44HOOKZkIKMFHyRdBJIjT7FTqsM3f5kOsAMOkquiDSlQ0CKKQhy+l0Y
nNTnY51CnAmWv30fVA9ylws2kVTSgx/OpMuK9braNrYp5Pze8ip7AF80kBjhpIlV+vEB6mev+gaW
QC0CEbCcfjR5Xzh0DGkBjdPeYdte1uJzSKN8jUEiIg1eGOpSMyEvOMgwfjtvxA28QgVlyixmFadP
m3bGGOzVklGwuewJWAK9OLPU7VPiQ+lPLgPFMX6zPaW8lAzT0+ku0yzmwLYUjgmmeCZqeeq3ajG5
X8oUuTUEJEhrSUX1WGao+WZJo0wYLVDm9qgMBw8wYdY5Wzg8l/emuK+AR+wPENk0cWV6H51COTrO
/8xgC1/z6E77uysso9um9yBr03UWEtuBmibswE2GZYSUT/vEwYznn/COz7dVxKoXbqRYFLI9NiUa
r67dsuR8wvjNlwddiwt34YuzoGa6PzeZ6MXt5gwqe7ioZxOx1nIpDtp7A2r2aPnNPS3xxkJz01yK
OcmqsnuOAtscGaZGheBI69vymIUuQh0v5HwQIGqUMvTS7iLbbDIll217WSmRoB5noBbrLi2AV7AB
XTXUHBNq1J52KJI/BGDIcJZTUaOFn6MqJOGsIcS+Wehfe3jn7N59vjTP6wT/d4gQUvzkfowlF3xx
e2865si2Tdyq25H/6FgoDK9loknq41ScdC2lEEdXgK262pG+dIZYxeXIrvj/tPnCGIFouEQrVfeq
CmkPiUKzp5LSHINB8ACLxfKZsm+K7/shJgoPtSt3b9yNUictWMMGgWKymj06xKtNW1Nzap7ZvNQC
qIUhVyQxmILeh2XwJ5AgE5CGij4vPYmzZOxdDIRXFGO/yeLeUsnxrdEiyWQyxRYrQfdeKlHpEXfK
hLWHvHdUiw5fYFz05k/sQBGAw8fuswr8bJ+Dw87m4aTZSzRrkRlPxyN18yvxg8a+DeQFa/Gq4TJc
mr8lS9BRd3IBbT2qk2T21NV747D7QMrVxo3H8Fc8s6aQJgEzBVt02TifmHLxVLijIZOgZXyLn8DQ
gn603n6Xvxfd9YFTB5IiD1qRIzSP7wWLGjzrC+aphB0Oyt/gOm19fvefPA4w5zHviHXX9VvXFR8T
F5oWeEq8wiuxYXj71ayo7VPSMjbR+TvhTJ+4mmZMUZNYyt2kksB43AjJKViG/S+Dd7Bys1NjiuRb
F1nf8DzRmCrzyFMt0cIGPIYvZJ4FMXV+LKc87FD/BiU6eN30tPKLr/T0mCqlNWFGH5FYcOV1S4Dz
X/3W2ps+niowDlrnkj8ilJ/f6Cs6FYRqvkKLqb42D8Ki9luJthIzhx5akSXXGE87jpMnbr61nJoU
035hiuaX9pEmt/5FXp3b2jGRoTyW1VczVVotu/WHVOrKha1d3UnGmAT5kkob9Vi42Bb8kYBNZgFM
oGaK/cHlSC8WgL7IyaQcvx0ek12jJzzg20BeG6t5AeXOwfIYp46c8NGKdxCYywtEob52tytJURl8
EPworwJgjIYPETSQ+nz5zr7OK1GdmnCwDX2YJFo9HwbpOutOfrvtEI1VziWI5wLx8gAyWLFMIz6N
dovk/KfJNGonDneQLNQF16Wg48wdgpmngWdaGfwzSclTazmLY3iAvk/wW8UYd+Bk9tFden/DAsJI
wqjRPwl1GY6dfNQKPG0DVCU5w1Na1hxKCH5KFEHCtsYQ4EprZllIvLO3skubJxfxDdZRJASGsybc
9mDpLC3j02NQJaUOGcx8P4frh97D9D2wxsG0TNTY+U+Y37P7Hb789lRcvPjz3CPPT/Jv2eDeUVq1
G4dcK61BUr+miLDb0vS2NtCYVjkJJOp4tje16QE57G+XmM8K7IpuvGa4Hvw/r6XKjuiTBWpAWuld
92tvB8K/Kgi7DsWJzxvAWrj/9O50Kkr0wxfNAy1CfYBnNgyyhMqraTwbyYLAHkIEgkyv4vrlxc8L
v0neoM3XXi8710Ap1YqaN6fsIICWolK5j0+LLVND1jqycQ8klpSr+RxeSBo/ZNIiIiSDUkbmmDC+
pcO26L+pkXcWogo3a9k3lKuor+XrGutSxwG3b4W7JOUFllAD8zzO7k70F8UOYhY6iGM5D5r7jPcY
hVUgqSm/folfHmxBuQboU65Nurp8sJgV765lS9aK1dNmvWtKhBFL+ApHT/9wbAd3UcAAr/kyFRTc
6o5zUFGLsD03QOiKekGEpO3Nm9Zf4bLx1Bgy0R6r4fl3FbzsTFpth+dSK7Mb3BjgU4rKozA+ogA4
MBNGTiJ51ipbleFhUs1R598A8cFvdZMAYVTG7ygWYH50fe0PDZtZqOw+3obCYpO9JJ5SwXv5HBaz
cTvYLS0DkdzN8dmiZQ/QedzC1nqP+Odn4JoV43omXB7spswPSREO8wA2d2+J7DP/bUdaAv5NdR7i
Xl4DVoAp+Ptx0AbRH8y4el5hb9RtRWpq/whRvikH+0YRxxemzmO3+cn2nssBHIWCXHoM7jhVSHmd
FiZqRMM0HVJwqbtpxpvSbLTSKA3kHIwTweQcEXdS0tWDi1A/KaJwbH6Y1iV+XIXO4lnzpAFZx64L
YF4Rbjuqxh7oCACQyENtdpEcWVbpRvW5dl917AG+9EkORD/BvKpK+32qdaomfhPC4oj6PW3KkSXe
euMLiKO6eYjY0gEnZ3HCLeFt7H9AlnStWycaZETiDU4fUbXlJIpWJbjEVgoILXlT8sc1kOa8ayAa
LfeOMNir9Bk5Sa8p769pS401anME2kIVw/3+Bs4Em8NDr3lSXlzgRMYTAPAzNbs7u1CrItnelb8a
ivEW3N4jBgmdBXpxw+gtIF+tWrZ2nJHUNtZ46jOTrybGpGn+zDIwARMxyJqhTYcyLvNiaAmSbbVC
H6vfr/Cin1PpI2e6fa3KEBmxaEyaj9N9P0I9Pav7Fax65WNmvAzsU5l5XAhm72PIL8P602szvnFd
lEq+U3FyxcabTENRzpyyg1KjjgNoXAUEH7jayPKNKLs9Ws20sdNSm/EtYfnAbOJ0H09ze9obLRPt
CgXXZGf0/Wo4BXYdg3BNlJy6dBL+RJdwarlIwWRS6Vdg6MH6RaitpC181tPqDEaquK36d/oucnJg
v2aU1mJ3lbHWS9PeRS9HLMhfDMprCdMSYkmy3g4zfSJEdp8sNFu2Ja19j0PnIxX+AFHImknmHGV1
WkIHvwLTFItddCBP6y2C614w1m3KUO8BjFvsyy3sYEXNXNK1Z6DSscZrxfdkutlgwV+fcpiIQDY3
kd2Ljmln05cvIoba5GEQXlikO8ssCJVrQ7RoYsPEbsYWD2LlkBRGoPUn8FsKNMegvtkLvNq+e2KA
0+xVg0bcE+5ixJ6AYL3vmTOofuMh2BewqB9HwQ3wL2HHmQfVsDbVLzsoFmcF6OzmF8ekbEKSqt0d
Ss4KWIuC6XzM6oZNZ+RIdchZ+2JFsBUy/GP2hNxkYhvwfV9zVas1vxT85/UwGogyJq/zXb8NKgK4
GzqeQOiYWABfDrFPrsp0jAowAxdPqrpKJghaznqOxOPDeUL+xZ9m2/Php3wgA7bAuiMH9Ty/v3eG
rTHKYncGHF8tE32AOe84de6jb4ICtgVS9rv/rokwuq8n4g+N7KpJsXQnvaDRbIH7nz7yfiASNkGj
B7j21wS9mdc2B3T/NTULBGHuAvSkX3w2MtupRrWB4/fmJ2OmrigAI+oyO3PtNnu/0QrWN1k9PZ3u
/+cjFI/8NAkYjOkVvhaoI9S2K8Fbv75al8XOBQDP2/DpL3oJfvGrVDlgVOW897L+erDw4xZ8mJK9
UpVl80JSndLVY6Y+WjVmVIqsmPHV3r8J0A1q/htsohJl6ekPfLpq7bwEPRxFPKmC1POFO+7dDPgT
9QH5p4qNQ1INEbo2Ov/O8ecSJHQ6gzZO3NrANeC7FAwDEknGDwXHjvWpu6K8do+91nX+36HdmH0f
HV6o2VObHhQq4DyAJukmWGuB+E/oVdqDvXJHMX+0sUwZGw1qzIujQqQ67uLWynfY03CWwfs78EHi
g9ZOGc+rG8jgd/TU0+tmofu30uU3azOozIdKCLKRuT6ILbEDCikXPdLetvxcTq5wuN+gcT0PhUWk
qJEN9k48jSFW9IY9b4iFeQyPSfREtGnD7UNlrRGtl0FDVY1hoI05oNL4CkJQ6qheKThKYOxTiMkp
K/UCIP6BUmj1DjjrZgCJYfjhLQgXnYOE+6k09YagNEXZgel6yAtlDYeJ3jqj9vFMJmUqKkwaN3HH
ZHT17BYX54GRY5s6hudgqRTxX0t/JsxAKD1E41eBwaF201ylJpJsilzcxBD6B0CM9t6S0STb7zsN
bNvqr1+qT6D+mk4bQaxhM175E8qm9hzcCJIqGM7H+N+ukUEXWqH41mtrCn/MqK6DECL8LxeYStN6
IavxWDZX8KjB8WewUEwZf9m2t7TjSI74mwwKEMLJFXYXFJJNcytJ86jkB0XtPMMPBqCNZP5J7Kdp
GIvXmI3LXhEGI/vYJO6W4tRLZW3OsnASP1++Mfd24mMyASPCMerIwCYE7aZX0oA3DCEFQ+9UUePD
sqE4dwsKBWtESO+8L1ddXYCRdaCKxASPd12I8DEO1t6ZZ5ibDv9iqSfYIT2SLBQAD5ThCaxryTIx
USRE4BWRmLreu9dI/qWqCbMaX687PMuru+im5aRCaDNRZ6mVwkL0LlDQK0i8VCdrBUSKO+vTFANX
wBjsqNuQXUH7ukkn/sBV4j/0C25XhMHIcXWUA8DYtmqQbCz5jVsO0u2lV2H7qHrowqoJBlpQ9Ma7
U3vJ7+fl6361Fp7HqPNctamQyYgZ+rTLnhrcxdhnW6TeFne1ZW8fQLr1R0kd41t2RxQROD//6JqU
5lo0ZB5dhmrYmzv/rUFHdMsCbXuwhn4ADrSTwOUjZ1i8/KQ0oRQCg+wS+Y77IVxgH7JYLaxkh5Lj
OgU1FOHgk34nAKmSCc8rMtS1lNzHppokBXZvp55swg+SH1N3herO3O3z3aaratSB9kGeGLvtP4hQ
jnRxelEk8+AVKCvFLy/ftTPTTF0uqx6NA/l7r/s7KfYEnmoCGi87zpQ8/ezbThnhmYy8a0JJnJO1
KnHFg8J4/LtfBwhtwLoc+JWSJzLJ5JzMIYVWCpMDM+tqdkW2x/G9prNh9CbndHjCgu8K56u+lTq2
yI0ruyxdY08AaefywSOL3QdEDUGSIYevvuN0pEXtGH3JySde+lMswrU23M3342ElEOA6EbSQ9yVs
ml0g0+XOXjJ7oBO0cVxtb5QG0wHcnv8LRtl3ExE0N13CIq7c0ba9xrt5sXFg4wac7ybDB0ZRWSXZ
3x2o8ghv7dHDOYuedeES/L9Vq9C5g0/t5zc4DlDUOPYoxBLu90/7BOsrh5XEXjKv9cO3tepguefE
Bz7kgE5HXw+bCBwtfTL8KtXIo3NjDp9EZ3+HRphQwyWt/qx+xpain/cEka654YSzbWA17WGBN5lD
5O3dKTbbMeCkPoQXEqYVi+yLLn7pa44RFyfnIFwpqDlqtiNOxa/e7ddJeibS3LfzGh/fKJez+yor
L+lS4bkB0PBFx5W/9izMuQ3mes2Hdh21evJBjSwUKX60jO6WJoCq8o3mXk2p43vK379DCFbTt/Hi
Np+G+4ts3+JZebnt2n5X85KBb7wPLhO0viTDsZ2xKSpgaRxSrHwpLp5G/hijn9ri9bHuESVqML+r
qKXOvfHK8d/gaV65N5CDW6FaZhFukpbPoQ7LOu3XAJp7coHD+d8f6pag5bAQZmNgOBSo8efgimYc
rYX39k/7rKapteAdngbVBW7PmLcyicK6qC6fpbs0sSsgV7LahvFAxju9/9NgELxcTZ0zODNe6yZB
6BkUcbz7iwnTR32X5U/xKxGhDTfJ8+k3Q8gz/fC8Qx660rVweD4ka8JiRQdRHyP5ACFm9NnMlznj
z9bH3aNTgjM+DtD/HubBKDNU73tQcoJITqJO40hVcWvM+LuPj2mePE1ZmAHrzI0WmyR07YxlY04E
3XdcwrbX6Rb91ghTkYWPgjZLhuftXXvHqMfC23DgLTioeRwU2V6AuEkKgEUQQ+6MJTkXwfnwzBwY
ycG30RGKCAeYIxHxLk0DPJgOjZvVF91qZgpDTviNkyW5wgdqH1A8nWfuji61gj0RILgz6oX1NFjd
u/R7bLSj7alMUJOZTJvgulV1Lw5tVgb5CzTKWeMRwk3RuihMVWEGNqrV3caJ1bN6Zp0Ub81Jlqv7
q2+13eci+42hs4OrLG4tH/ADzZTYj3ggHR9ijDoEDucWAYHH8LFJ1GIDbLc1X2lHd/QuKjsURvki
eYP4iyfLCzBhlZBTUF72HI4qU3ZYLn0FCixr7HmSI4sFhHg2vAsjA6rV2AITzExGqaOVzTNoIgVp
Lg8h+hgJDBP0v8eL8MBHP2L/gtVLY9ToyVLLjijOjojGuUmVgaVnLJ1RpICTMiFmQzJmxAFflQo5
7HxFr4pO2KfEjp4v4UiUk0fc+xU997ufPK7dTq2okI311c19Jme9TC2C0wRQtoL1rRNmiRxjbZk+
ZWMfl1Cp7Ops9DGSCoqcDzSn92qxPjodc8Qon0yDfqLeXFv34uhIF6CXX2cBorOsOdp4lj5uwkpu
HdBKFcwTlezbNfsMujxcYjvlncd0ADEVsUagLqVjvHZyPEX09jBCFrCfqb7iE1OD8o3ZiwH6Iqsc
TS1xsTadv4w+sqJPVrAxxst5pagVMC5bvzii3eepfsiQJQl0tXPKGSY4vCzwwkz9zJM3phXgcu8N
fmIj0cnFSRG162L/erlFuURAnfEazvQWe0AYlZAAlbTY14/g8k77v7kqO+fX6ZQnoW9CTSXnVZcv
bFLlKQa5Pmm2yyVxXDfvqpVkxjMIxTQKWm7jKOFNbcH2NntNN0BTsjKhopw7t9DrO7H3MOWsH9KL
N8hSPI9Xrf3NUkcjbBRG/njzy7EeON1B3YioIdCZLCyc7bNCJseKgr+rAJEX78ARJwqcKrTUOCsh
sllsbSs4QZyJ/msdYmag4tY4ue/dq/TGy8zowIHo97aeyutbyqZn+/3SfWq0mV90c/o4v86eq3mE
iWXrA/0vSLSCaDZta6RznWyFG7CNOryul+Ln84P8r8aXsov2b53+4ttpTnb8LFZaoBKEmnQ6V+F7
qIJ+G4Crvw0wcqL1k3qh7oxmKL0Fib9dQ/ZSVicO2MtMz8/2psmKlN1A5TqqHB/3rnTYmcT5H75u
qy7MDb2A2slaxko7cnOMwjfMPR++SJLXysNvMJiV/dlrDXU8v3M4XzdjP5NVMGz9bw0VkN+73bPc
L/ZHaxhojT18l5i7VNbH4ar2tEPut00WphGNou6I4rfEkZ3iExRtTRvhN7vFsBelu6ja/GyK+DQY
ssdEWma+XxwpDg+7G3Fzainp5KyEcq+sdNKcnsx+CcWlLGmswVWruOpASHX5Y5xhDksRDgYpKAW3
0XJxEkfQDDdiK++eM6m17UCb9IHU5yFRn+OSHeF+s/NI+J0RynEC3vOD3u3x07CA2MgXRBZCnJJS
0HKbBJm0CM5q3RHrowLLrHnlzadk4hNmkzfZcL+A52+jerxXe5VsKiJbjSK0TkzXE5CfKtFi2FAu
FmR+X06O4KC+/GtmgUNRK0AR0HcIAxB0QdjlzMpgqPwlQ4T+gGUvu+dBay9q6nrVP3OG1flMR7qE
w+x3emUPVAA4z4z+G8okJ21M5jtmunr6O0zD++rKcqwUbyZJOtloCu7dvRr5YUxcZybtk/x2B7Z3
K5V/pvlXNYKG8E+08O4KgG+Vu6XamKrWxOImHeqfZmNPGieZ3mWdbWvAtzoASW8uI4vazv5M/oVs
gDVsiEMqVCVUIt9soY956O+hEPbID73VjFsegBuAUUjXRzGoKHjQ3Sdx5ybNQgjNvUtWS/4tRt3r
qoacaMR7rlTDEJI4TyeeQBmSQM3rAgcWL0fx/ePBt3BTz59qltV2V9ANioGIZoZ4iXqLxUopXK1B
Nwlsm5cGJk/c2A+2bIjEQbLbS0HXz9zjeHFz2dTLnGMnVmlPMr7CvjskScZOAyRjPEg1EdXiJdSA
H0NqdUX7W23ds+fyloSayTGSnKIbcigsoUEQQqxUPlMF26ExV2N4oFFJkr8vm7VUsZAlJxJ77/vx
5+c8IVyR9kGY+TSzI7VckFTy32mXAqZaO3sTce/ECderjds7ha6WhQp7LaAbAcEowDSKbFkRysZ/
MQlAmCUvtS2kPxHADFWmVpbXYPJ3BP8JovgK2oQqU9b7epc3sMhjRTpvWkR/ceZm6kUFbiHH4+QI
MnonIqvTBmlJRU/Sk/lh/NRCaPlAkHuEn1utoAeS3+mgwwM5Z6FOnwHxkKJFDSuWB92XYWBpPEPk
+nQBBCnCfN8iZ1GLcAyPY7QtqEcnAFPET4LgT9Wp30qAMNtRtVb4tfvgcx/CE17lE1Ajpsm7aBpm
BjVZI1BvRFimUUsZeynngPnvBtKBaJrZcDM0DNRn6480WTGOVSTI+fQBZtCr6G32B3+m4Ab5rtC0
3VybNQkr5JZbdrko0fSOdzRjt0bKXyxopVW5LvftLYnnWp4bQNHuSVuZw6ebD4d7LK2TEYoRfFsa
zhDHRHuHxyeJSPmxxgoWjHXBMKYYfAaGEZDVP7szR6jp7ijumMLMuFcGBaFXPnGYIn8R1ZgXe2GN
wTq2bekT7Lbt0MqS8Q7jH61fy5+JbgpnPl2KWBxY8kDJiJZLjdoK5bry+zExMJ4GqT7mWJTW6nZP
hSN3nZZ/TLOGmqd0khMglLM8saSEEvu3GrTVN41zN5zCti34Y/ZO+Bhij5NJPvk+QBw1HKhuvVDf
LWsXC3sYAtdD3T4+iKLMyGiU260oay+LpwEL/og0FkqAnBJZZ7iHSQfvSRcrw/tR6joOJCTUfI9V
Hy1XneuHqP++uJVFqoUWa0LuXbrVr3JbBRhb4hiZIfVswl6+6aYnjaE+NIgnM7wNg+ylxYIdicvU
m7hzLfPQDfkDmRaNEKHdpnCRhXZ47W59woW1rf9MVLlLsxGIUx+hRAoC2QdjqlARE/Cx/SPRWacW
frx29NSsmaIxkN/OT2bYkyD6bc82y1tsYvKs6McKr94KoBKz/7JG4nNj9OBD/B6ebzC7HE89RoO3
cgAa+Xd8s45XI/npySUw9Znu8XuQygwgRSu6OO0v/2fcXvG8dJkN1Mbvkrmd8J0kUaaXVo43AqJ0
OfuKEQ5zQcQOys/CTsb+iNpHOVSDmk9Yh6LZQ+OmGUhnEN9snHnkqR9SABah1mDquGP8LkYjirkd
t70o5Pj5GdYKU9k7mnox9o5ycL9hwbnLisS4aN/aLlGeOeISZhgZX29BYMtnyXJn8fNWWlBDSTPa
tGhdhLPILv2HUIuOpl273piJXlsuZhRvKx06L31mexoDcQMPMpS0sfDn33EkW4CWtmjyoI2YQTu2
8XwP/B0Xfge+aXnre4kx2udxfyZYnF1zjwwpSnaPQpcd7HhHrH14n8gZulJ8fPYH83dnbG0yfzW0
Uh2yXjcL7iVPbluAOOnpcR9BPK13zbKEP/zu6ArikZrr5FGcD37CmB0EB8UQ1xRZ6u58y6HW/hlU
klH5mDSkpuZfxPA7vgwJsVeMY+fOYCVSItYpv6uzdkgqx7EaDzga5C5QfbLxntz4gwex2nHpak0w
45gmdC0th3No9ymH0PmBeUu6r8NTtv3rRIgSMDBBDTBqk+NiBBzx9kGweMjnx0dxuQhsoHgp7mKk
nxmxQmyJi7GOKSc/tgus3SozLcz86wToKAttvWGsFF6Iw4BePDvbd6CgfUghdJS0Y+hHmN2bZDrT
9lW0C38bEuDLbfkukQ6nbxP8nHXPuMH/yMV4YyFaSjziCx8iKKjsvbYJGOUFTqDe2DhAZiaoNB/u
4ubMlejjmWgxx73j4E0iChZfiRr5bdDDdS9UMhq9YojdUjol+PA2hPruER1U1hmWP/TaPsDyci45
aLMh9z4u8JJIZ78Zr5xcdwQlBF9QL32xOlf0b8WB18hQvCP54T4oP4n/vjw7kb+cVsGx5aupBfSQ
g76J7/FpAWu440qysXu0lbeV6gB8GEJgVItyKQsh2N+RSG6lFg9VquSaYVl84SMZXqoYJCAaGb9y
qHwzFqcP7HmyttiBoCgVIdKYtz+F9EZIkvQ+qD01XgGVhBWAGVjuG0CCpgbxQWKZ4sVjSGCYo0zR
lMFCtEc7NbwAqTfS4tAnTzunzKV2zkFd7kH9JbwRnOw/8N2wY7KcjR0UBzqaSYPCdfFawsLkRQ19
29y5Up/2r9u8FnqPmBYYUYDFcCs+3gCSDeGV3z2r+oEvNaFd0ARSmg53fsLvEph815gkFkHGjbYN
wkpndB6WKUnxrUMj/7GvIKSUF50nB1l05ryrGvsN629fVijv00I9y5ZARqU+0g7b7W1JybKM5fJg
lxgF44i8ZmlRLxtUBEOKmTuya1uEgnalCZwStupgqOcvQrYS+EhHk/9mdtjxDRxsZ0bognQmgbBP
Wzij6mCQDZL0sHfsNvnGrJWg8U4sjzNiiWlWdEZjlfPRJnc7UhIWR70auqfXmcSRA91QYIHmTyyS
bjWxShlS3JDYqGcM1t6Nl4wc6nm/0DDcVyPgys4dxYguj9jqnjI3qyLKcJtEGb1hZS9hoY+PTfep
iq08crU76X4ztKPZPNYly7AuGV8uclq7C0Lbehz7vwRXfmVdMUsRaeRjj7HnSnmCgseDDpzTZFAW
Bwjoq0KQ4AaGGQpgsWA4OoXw3QPnlUlVGIhnlrL17aLR6toCcFUfkWzUh+nwqIBoPvV9o4D8gQTi
kjEaHiTXFTF2d8hNBbWpOzA4Tvg0Iiw9rgFUo458jSCdF2l1NQ2cfN8rAEqFbDJOSRzeyL0+pUbn
nhuoqm/G91ugsLaXiO9yVnfcWLSusJVCa7oLJRmTaMadaSmPFTSKqMKs4+rGfYnX1G91XOA1zVwX
zWW5D5ztmq/CeoECTebINrJJnS7r0sn1sTI+XDyWW3IoK4CRBUVekrUXgWp4ZWOK8ml5rP8FHKVl
BGjpjf/7V70r70AQn/lsVFWswXxgg86gBb6LAyCeRI6a8RSXt8agf9KS4jdtQSjwBh1HqS0a4W3X
pgcfz1yg2UgpUfP/JdnRzBHuHWmOsyjZf2+JqdYneIXE53VxpGyzgKAmcGMlpcr8CcD6Y1NBDNYY
FFBFFD15J6cPZ00fGa3wnPi7GEiwswRUFOp+qC7C4IzL7yb65BzwO7dt8NJoA6tfT/10xvlwkUXu
b6ZDxMEY/E7gG0LC1ZM/b7J4Bqp2inanbp3GvJ7Rg2/050n2IapLvi/Zo+PVENow6YIPDK3KjaSe
4y9YvixkD3zf8GRzyEDslW628t4Ow2Gm7ximtkb9/ualh4C2Y6r7r4HHtbUNuHaJFvyLdvz7Fkf5
gj3s5hvtW2Hd/o4hPws0gLnDSXVwPvaZT43UGxzRv+RZVrxmUWIDRC04SI+7FW4gnOl0gX25zf6K
S3IMIIHRvA79Ky0CpFcKUDuI1PUvWhkc5K8wf4czXWSsTJLKraXzuD9LD90yY9jQYkl+PlzQYYxh
xLz+I4O8H88mFy6DpwKilHEe+5+FzGdRMIzYdPVvBb/azCEf8xzpb1VZ4CV6nRWUfBs4VP+sqzq4
wFlRznpiDwumjip1HzBXfAFwyuDxF9tQPTHRk+EsJOGbAiYgMO+DQ7wyqlCscXX5tyVsfalLZM6l
lCT/K3WpBSZB3PBqpvqUUgg5Agr/fvFnYGGJF3UsrmbKJBfsoRYgjt8BqwyjIVdZhVnYRFDa5aO7
4FNiE4lOgQfQDgQp9mvehVdKl/mJS3uJnGbORlr9Ptcbe90c1a7t9cdpmH9uKibIVoQ8ur4Ihnfw
yDKfmaDsZ7e5UcvOpLVti3idFTrV5L4QJqjZ6nXjfD9jn9pazZpMmG9tNVi9TA8mNmlgBWZTTwai
CkyL0oLAsfYxg8551cXKTBFvt/YN+3L5MzbyBLckty2PBEDv3TTCFpmRxSSJxnLCaVzY+MSUNAm2
7PFOC2hbRiFjH3NY1s6fAZ4J1f4vjHJ6/8Jn/Ij9A6l6kkm86r7/92nqKzVjgkFVo2UAocS0K0EH
ngHc5X6AntM2cAUL3WKt0XCS2VpSaUGNgk+4rDicldMXiA47WJav4r2GoUYQyTBWWkz8P39L/fB2
RKBsQ6vxT7I1vG0h5aXYbARa1RVxcO3UGFf+nGuHPLguPjLa+z5yUUrZoJTRGtpJUomDAPscT+F1
3LPqXtEHyUIRL4c1N78Oo97+wOf/cJ5l5To3dcwOm+OfNI3tF5oWiYVVHdn8KylXG50RAntlChzJ
HrLOGPNS291EztOyW531nH7H6HLZLL6RFl2pGPshyPaojZWGuPw9F/DVMUXAXKZBf6ZnjCWeOOEG
h12vHN61aaIFDX7z6Kmgn8LILeDyOSAcHBmSfwZrFqvFGv+b+kPr4KXCEos5+15yCpTX5DIvGlR2
feVmVatY9y+eAZreuaoslK/35pHPCQA9FY6IKAoBOpuZhiuLds8y2We5b+3suD1lh1+SO9dHreCq
gCidj8VzygW1KWqP38B0BHBtWanhfogiVzXPpyat+MtC4iVVX8F4XbgPyOH2UFZC5AA26PuVvq1c
NfttZ9kQRFLyLvUVjdJWYaRsRjSSlOhlRA3nnNtLKPuPx2gpbl/MkcasHCmbYLNbwG2zw3kx4F0M
wBUayfYLw28rYg0CE90ILNsuvrjyCk5UItDRGI22UOU3oVApmsfg7lW7ckkbB84IcNamOq9tmEnL
Ttaz59DDHSAiDJ2wSTWLwVgFVE4LfuYwEQYjak8+0Fz2UPDe3uaAThnumbGzWQfTi7h+O3pInYiM
XvyIohLnBj2fGuFztHSueGbAqdo+1LwYBd7ooEk2g+Du56Ch1rscdf34+9ixCzhJ4hxXmRN8h/BQ
xAZxLn9tOlXJOuHU3zjFD4YUdTlW32xBKBZsI0KX6Jn5/rq+WAwQ+aAS2M/Dd1YLQSoRCDN9n3dz
2V5ccXXDxQbVpWvuNMPwttXs5A6J1wBvBT7sqLH1iDHtVtNWrmdAMnSVLR01jDSDvIU24FCxXP9/
MiIcpdT/Kd7rWX7ROSOvxWUC1MJhbjwm4rNOysu7sjcuml5vT13U0EhLdfuWUQ/JXZ1PhExUa+TU
yvF7DaVGsZnUeddZVpS+QAZfKbA1RZxPnkOx8zLRxOq4g+GVZkkmMhagqZ+jmTL2/OW1NOLjJDoD
HxvFncsiGmInnOKJSypCDLR66WCbgdBQHI3jC1UUI/SOqIjDlkWsBGNwKHSdTsXMMAjujNOi5NgC
CCZQnHXzrajpgC68uY1gpDY0isSH2IaofTmNe41eDBql751AMuH9QimMvg+JSzOBiDk/OKK6+cI5
FA14+L6gdjW8cIQVmJfDKvPnq3IyalL/7VhkSzl/CVmZcSwDYlpjOnWzGWL/7Ty6mDaETaCS2kMe
kg3JQmTC9JBWWwUIesQW1T/DcLITjPlUlNSwQWWMIlXTUZbbvSdW3Xo73gxysPeEG0aIlq4ewVSN
/FB6NWBK+h4YhlcpkYFOwYwpvRq4W4eTIk5BuFVc5N3V3dA7JaWxadepo7wv/TBV1tMlxfQLUa0p
Os9qhy+YP46I14TcUfhO9DRZ+P5VcxvKAMJIX0fazt2Ae/72bKclMREqfhdkTTWdfbGvcgYw4E93
nVJ4/4tkz5BPnhhcu51/ivJdn5K+bAdC9x0w/GfJqe7Jx/m1p+avTH87Zy0jpvXOTQQZqC9ICiEz
NU0oi3jwSD8IOvaY+tlh3wywibxBnED8Ur0rXwRvfN8Gv3GXcMBhATPHJcTIk8FVHxZ1xurouX3r
Xy/DtU5Al26eAFjWFrj80vegeO0mOvo87rW8F++0cjZYstGrSiiXpz9MZ31H+5KNvdxT2r46QhTd
kHAXFyHnKMAWTVxQyXqumnknpF+ZS+yhpUlzykbWvtSlGzlOoNpVWdkGBp2ZTB/+ZGep+FWgEyrW
gcdHqHl6zK/wDj+Ro+NA7nH7jG9xu1fWVt3vdTDuLwdJw7F8sDdv9qoKMUHS18w07/YmxYnz2MfT
BZ+5inJKtk4pracAxO5Wl+6sWzhgn4k+ykxsdL+In8kIdWHBUUIiVgYvKXmMMe7LejjD8Dp84zys
ptjYvkWpMDmgqC80qb8pbOh99cFjipGdbijBz/ZJrBVUNCr4hwn5ng5u+n6Lzs3R/DExwexA6dlM
V1/PVjO08vXfCGev6oiAQELvu7Ne+6tSpff7A29VaJoPRwZkQQ6xTzZyJln2BC/f3FVYkJZ+B+Rx
d5WX2XGE1W4xHQNPHIW51bmjpo4zZ2+/p0V6hXy2zo4WXDqris/DxGnr16ufzGQ2ZFGgbzlnVQcN
H/8Ssr0og2gXL3m+g7qQp+aTxr35tZraQEzi+c+MxAC6VSILDTsvcVmWllaIleBAlOLn9KOGeIbI
3pixbwYPBS5ahsQqYSt3S2PgTZRijNt+TBhDGRoGaRUlq5nTJxsmUvYaH1Qu3xxXw6weiqXgFSx+
UFwezgS2bXbTfOsWFULKdVEGyFviXkfTtd6NnaowDD4GsmANil1TXba9dKX8oBksrQA4p7Z20Ucn
wdkBYydnGiUTLdbEuggnzXuRTSt0lQ0zpou2/FR7+mohJB0dU3HXWxPceLb/BpGw+/aclR+Vt1Pi
74fHsHpD1Qktsp6lQG3kPOSpgKSiBd3/5DfBic6/pz6K5xoUxqpg3L/YDWiewWPus9y1nVsPA3ei
Fi+I+sZT3kRtwy0avyuqjwF3tIAX+HASm6sQq1nptGc2PPgMfU7m9CpePO3+01i9esvXEQcm5Y7t
QRXTA5xTUzzSVIbqzimTboJmDlmd01IYwu+rd+x19MmuvmUZn11wMXP227myk+vAMm6TdR4pVOZS
J4NUqwMItZRzSxl11tiGEbStFlu6KnQBlG9Vo6ggNASR7TR5c/+IqaUMGyvEfxDFxA789cM6Eo+R
Ki4cfBKW43uFJispMiU9BdnWkNpjX9hZX0mBwaUPS5n3l2Y2+iaTwa81n1ZwkJH8LTOqCq2qxOtm
hgkH3nJbQLKWSTEdEMw56BFQ4PuNorpgPVHeq4oD8KlEW6E+T7aAY2hkRgNpeUE1pfEN37ljR2Ok
asBYu/bcAkqE+UcMEf3AFKsc4vU+tvtiaLJX3Z5TFugHzwwwv66m2i+qn4Nn2DHOH0C4+FtMnt78
bSgZAnKydIkCDbyVxQqJFBO9MHOZn2FyS178/XWFW7ycjZMgPK06+NA1V38IaYWjqjQxUVG14HHs
uOSL1/sQXg7UL9DSe3vN3s+KAciVm1U2HWjzC/AZyD9wnoHnprs1rXt6xOK2bKnOapT/kLlDc+BN
FVfOi+GKGQ6sktmdRvq/RONp1cqp3Iwq3M5qskZfbr842jE6HIAIc635V9hPsxF0Xp9xSBM+m+qg
7gMe94e1iXW7Qj6suWQB0ZUNhcJcFP7szs5CPZZw9JnND9krJWGFEQjp9XiIRGg1PCxIQOmrf3Y8
uIHy6R+JBiDj0bClTWHpsArMlUR5ASzLnvp8EProzG0/MW/tYwiJX3k22NhPaa/nvI8Qgdzy4asM
x+JVuV3x7Xmd5qW2LUB0cvkV5wsC3DWDEBaxCH3xWuC5yAF3ezBXT4tYBT+zFQZlFCT/sapEcu9d
bezB/1znBI+hOY6WnX4aLwxTV4UQHdzzFgWF2rq4WWpllYb89ebHNYrg0IGkbRgjeaNM09U/rgnz
Sr3cL2V5frUMpvlXC2h9pfHHp8Mfxz53jy4bsFT8/Qgc5Z1DOUwYYV4ep7mu2aTzRCQKh0IROi32
LfqSG15c6O/4w4Cd4cbGIFM8kccC5bBUNKR4HJp61eSDdelWA6Pup/x27H2IdS3G63I0hTX1Br6X
Ta1y/WNfvSUWx0+DICdhzWhB9i58tWVZbQTWcAcSrJOdiJg52sDxXPGamYqSEXiQr4/LFvloDrx1
N2+tqQEIOL3ZBLWEUWrRj3i7zf9j4C/lfERt23/d8TntO8p8lHYw5UjuZHt85W/CSeE4bA6wrQA7
XiNQb7kup/BU+eoty4lLur5YrC0vtRq01ZeSsMfBbjkPLI5w/pQVNQb7X8ndfTtIHgRrYykXmwul
NkSM+uVN7b6WvNrjYEmT8FSaK/RennRAFMYE/Sq0/csFqdAS672SbXoXJ20llKvlTzcae3cWG7uS
wcyQX1plMxFMdP/6B1fpEfCORPeh8Y4DyIIoVnsu3jy7nLlV+dxn5tXzSjz9et/SI1Ua6+QIWp9M
bO8c1BV+ShtjLbatUaxA1wvjb+Jn1WiFJUALC2JWMgDNJzqhS6ulLg6IarTxkr+BpsIPbmqjLfT9
KZnENGNBczhgt6llyCsvFE/fapFFQCydx1jXMqHDl3q5nEnxnXyIikju5ThYRqF4cbfUmL1oihWA
KueeEI2OINUmVP/McAS7x7n+Hk/qeV1IS7C1I+sutN4fYYiTyuuf8BjrBh8Oqt/ZbKySVGAPiBHy
Iq+0HVeSgbv5sG/9wMZ/XUg1WCh/bPmPJunFcwWvVuD+a4vOtL4ctC8VdtYo6n+1DEVHQV1O2/z9
TeH9AiXiayQknY6aAwWwi32ILFmaNw0/QSSniyCyoRt6fK+yzmzkPivKE03eIEsPszlt+ETsmZmW
xvYWMANt3fovrdH+dMtp4ty1554osnn7DbVxhKhdvYwPaf+VHFn37AZTz+fl8DjJ1IFN6WiVB9k2
T7YNGUwqi10DquI7neft2sfW98lhl6B2ZFnWaI3I+fQoeXdO+sBKYFajZXrQBBdQdmuy7CCobIil
EYzci0YrWQR2CgTfuSUvfkcxKQ+ciVP3T5Srt/hv2UdxSCkDgZQa6RfHDgfAeIWxRutSF8lPzlmu
c6u1X3UZdr3UXyQJQBoBOi0FW4hNY0No3fuYS/OgfJzcovrnGyf3rWI0lB3LHIeCi76WgVj2XIsH
ch0BSdb0ntpx5WpyB5jliYKKumd1Z2xA07LBqIryT+RaxS8adlAOUVTOV0L5urU6GkhaUk5g0yXW
JyUHxaJtcXI6/nKOQjelbW3qxvURKGZzTyrcaCFuYlN76Uw8IthxtNGHlmwvrflndcfCgfGYTnXR
JVgtPtesUWK/vN/7whYRbzR6ePdu6VPToATLGwPuZXtdczNd8MURuQFynUCgfJXNWLPMXq4DKy8d
LTZRsDHrfMLVD2c1iy2DgR0SY5kgBM7F6BB4d3TMrondONm1dXaQGijMcvAZX21kVEugYcEs6XdR
17rGCXRgTUXqTTj6XUybPlPpEMyGg4MdBr0CKwkdAqzXBcOhnlHcNyDTPngATbRUvrfYgoynutGV
g0BTfeGx+w8GYi0tVntBBj2SGw3aYxM6xtbkVfSYvfI47QzctKvfa7eBDTba53CarPyfqiHTC6fT
bEp7zaj2OYfVF/1N0HZqLskobR6GTR6wSz3+judx+1x+yDa5OzYtX47EE5NaAszHMEnT6okSsT7k
vBFFqkQnXd9zZX5SBAVulllaOiWJuhrcqCaGR1ZLZdCPuCmIfJWlnJhaUA5GzZVT67LPirm+3qzz
mg0Jn1GIWs0N5Z9lhFd/6roixnWqthHBNbnnyLZKpNMrqRdGPhJ1O6VKF8cfZjjvcJAP8vKdx6m6
gjZKlXsEkiZMsIL6gRImT/LW1apmAahDpQKIWjDsVVQ2buW2MCXelFO1dt0yMh8z8UeaPJCsPOwG
PH22ig/ffsnX0MNpzA+oxKVKyHEbf3VucgSkW8tweGs3RnCvNWNYF8kyL57hfa9MgH6MCcR0wxVL
nHMO2JgmHvY8zdtNYbqi8xei4DacZAhASByH9AjYtJdKWTJwgJVrrB3vjE5CPzB+H0LlRucWVH9I
mL78uE8M/WJLldIrpxtECPNK9pNsj+PZWmzxTzfmga8ItbxgHTeYARXliigkDj5kdlF7xUPUVG/C
cDhJll9jC6HQ2Phg9qRHU9vzkggAiV4J0OjMFhV1sfq4Ml3GHfsiIZLOuWxc5ea/Qb8HiPrcR32m
QgwfUXWB2v2SDohvaMe4hJ4RtkEaQcRh9pcf5XH3ehesvUu5i5vXHIfrRegp8780DfWCErAcBo/z
TgKkAxq/1UgtopB+BtWinbGsSbN0ra7R66Gplpwv3XQihgBD3+LRAXObY6J8rvYPmAJMEVTouqWD
iHi56GwI9qiF4ePy8qqGASEXLHyWJOh/NUNBK5hmINTrWfk0Fm+l2+FdqmH+TeuKbuTc5iVLB7oO
EuBS5FOkdrn0UVDu+yFRaBTuG7pCQDFCvE/v6Hmt7p0oNtqQQsdjaD8aREqQpInwbMf7U+viMfWo
ht40EyHeatsak9KPu0gLRTJValMJQL6yLX74QWaOuQkvRAFIdl1LGnFTcZCLutH/yMlfp1Gkve8c
Hn4MCBV9CHE/BRFK6gPQXulz3O3P9pgz1CRU0e7KsCAV+QsglGsEwwXEE8AQA0fxdLFWJAU0L8dR
ScoGO7wEVpFe6T9HKvtRF0b42SzgWpUhRGU7zefOpHu6g0Ck9VvQx4da3aCa8b2nsFwLdwXnwNYb
oAblnnKG6oS1i2WgVIPBGa27BMNCbzLetTJgOa4zxnGILkYdOx0uV1oRKL7rDQru4mZWGaBZ+NRT
vj3kIYRlNi5XwwaMHv1FznOFbV3rAwrjC0c/AM2N7GIbSAE9rnKJo9VAUkw5/M5KzX3SgKw6/6ba
9JWBgCJMODqbrR2bSZg7axz1oVV4wYcWVZElyzgvTz87mVBkFViMuxIPbz4DIL7ad5EPCu5GUYH9
ytHCFonOk5wD1Y0wfloxs8KK6FosPPt6EqCU4GFz5CQNMG1sy+DalxeQb+0SzNVxLATZNAZk5o0+
vx+2FcX9K6dyFgmQApum75P5ubW6Qsz0IPJvP4KkAQenPD6oa8HIxMxmI1/bJDpiAsr3urF6m5pM
gjp2Zr4H4aNzmw8r7euUJSorGb5tSOs8QKQvgLPDP4VkF/1dEJF1fODZN+QuTdRfH/TeWuUGSCao
2mWfepTekVfx1h1qYGMmz+l9cWYBahAkn3z8Untr/l2Hgkjo9Ip2+vWtNwHjNJ2gE4WMgwl//Pb1
D9+77p/BLc9MOn/lPyaS2tDhDsv3motLnSZNCPew+HXY4ET3quIEsmrh1DLGaheIt4B55NbS6MeT
s7Em0JO9RpTilctD19gl4nQOxm++2icvGHKvgyeKHvpq+fMDCd9suejFnt+3xP8CscMT1xh8uYon
l/K8zmBpS1twBPzC9jDDS3JizK6yD/n1EnWZenBLXmNlHGk3yzG+YMd+0KfW7LFj3XyMUzhABQwI
VcKL1sBPIZFjJ5G1vR7Kkoswdtxt7M0fsA6zy33tZEhbvotxFVaphNePrLmP9QLwsaTCYoc6vkBl
YsMskUux4J6+2C71+rPPHEPjztzh/5OE7jS5VbRriGOnb6yajLU6iSVQ1Vh9n1PzSSDnLtFwvODp
a6lBxOWBG9O/5vZiRN7SBZFrOV1MPloKoK4w4I3pk/Q8hSxO96eV32LgaWtDgdRecNvyS9Iy1pX9
O97uggqSI4/Mel10/zAGhfsNfYrXFKXXji5Cps5UBu1ku+/RPsgz+f12S1zTyq2c6L4dJPM2SMly
wxBHyWhpQ0bcKW85uTcWMfzKnVFlwnstMGjmRuZNSs/wpGQG82lceuwTKtZszp6jV3XKJ+tOfWXS
X7/BfFSjhaUFUC2SYOarbxEh72OhuNeHwwzgfbb19ZKyHAWNM8F3/hhOJKKPFC47x5P28tzC6g5r
8E8kEHJ1LbqLoYcgXKyumlvl1+4zOOtGOZO0PsFo1tCYv8hu6bdBBoDy0a+hHKk4C/L8uDdYAGJ9
+CNvyE9CJjvbAUNW8BmTYU+8XVll57nXTn1eBlYv+V4Y3OaNcZOulKG20blC4fULEMYcRYZtXoSY
3xn+/RvRZ/a8GKtMHsZBqwcqFPwjPjmRBvpbc5bOYmgur2QXgxvmMxibZAmE4YGRb+fwh9yqupfS
yeCHLZWm+LKVJtqfMa0f1chhyDT/gJqdIGyUtoFk4aygZpX9Qcz8bAOxFTdUzfO2Y/wNOcFMeNv7
0ojoLwZIHSkaEfEsfIjaxSuKBrrU0KeYaRpKQLr6C1JUubhcVn8V9nNMAXUUGDNltqbVWuEwa1Hd
lXvDJpVCJSYXFupCAS+/bGZA7TVk0MdEdX7pGFIC/Io3i3AnPBbWqAfPhkU/dOzg6zrgakkVVLJd
1gT/Ak+65tsXoVQJRloqwVX/a6MiMbdq2sE92pkE3Hv7WVbNNqphIsPTOg7ckXdmCmkryYknJpDR
BqTpyRwXrNW3iM/4vl0AuGXfol1Y7bpjetVaI8zg4gQ05Q2pGMLAbyLht7ih1uMjxIWIShe0coic
u9I0lGJfCyZWoGWgycV8c7EJ/5G2jhWzUoU/PBt90ggnbRLwTa/3u+6rOq0bz6K2uArpwdoNEgPI
SCtPJjE4fLHac66uB0u48rmhgsLYzSy++bnUanCYXCpHs5qbk4TuKPYIzcvccAvCDm1G4w0R5VOa
BsG1HYG6jci9a68gKmqdQ8ExnDOIpRiDJva0Afs+M7DwB1uHN0F5PUaPXx29BDEt3BFJI/Omj/8G
TkXg3ZdB9+hM3KgWBscyjNXDsj4oiYbSWUcsh2AzgnyxxBxf4DPKNvkeaIA06IpDsOgC9cafKiA8
EWH6QnOwFJQ4+QqhFNAlBR6GOWMrn498i4+sRdPT2F5sg2DSqLcn16NFHLZ6ZL0MvobJV04uNZIW
LfxjTmrMdaxUsBuEuRAN4MxHvxxMjX18PDJUqLq7A6M53oP1kHJtj6IUroRKbSoDrNLr2cY6nKTi
qlT5YjmGkCybPGme2l512FCHFx7v2jO5kBCq6QHcsuCj9wAcZ1KZxeQ9wOGzNy+D73QUOTRlkTOM
tsjqzj1bP61BTuetpfWXRlCWEDtWnF/N6EPnuxgO686K1G9S0qS4GWf/lgq/y8x5Kxogdj8XkihX
fmY7A3NxAOsjqTL11j26282i/oodwKpZZPpKEMDF3XQQMUD82d7iiSyyLzXGg37LvrNuxe0xL9Vr
k8RFpgoTVkFsoam+2Z2JwNcDn27YKNbrFhdFzG7cMf1VTf7v4bP5sXRBO+jwRsSswSRSvld9EmBF
aguYTk0FPJts4uO0Xl6RAnYT9jOyQNP152DIgEU4h9cqApGUk0E1NAP9qsCQa8hA7HIqW8jnscu6
7YLhX1Y0cM/z0c5GpALBbduVk97QlgWk1MduNex30ctjRpKnoawcsIyV7BoSxBasSyWf/7I85IOg
SQndnkki94JCGfRLMNxDG57X0Av0gxcrRc9vU8Mk8x6LZlluxWMhdNXOyKvASXnM/NLcw7Br5E2B
HzY8SY+2Rnon6rj7NuwhVLw11zbldRFjs8Nr0Q1OCRfLFeD8vAF4py4K4AdwRWhK//o0g/nBhjQy
064YgbdOL1dynoY406sEDZg6iPfdS+DE6AJkmSiIA6Y0iI7rLSZ97HgD4v/MPym07qirHQdlP8Wh
rX1H2LyRHSD5lG8yqvmOkBQ+3zRi0f9FtF95pbYtEUJjmkoj0JaNczdLCq3y31qSJxQ/ChieZ3eg
48gDYUs6q5cZwk4pAnfzhXDHihN3BIg6qPHjlYAcRc/cR7RvlE3uh2B0ph/vzIpp/2TBlY+cNpWl
QU1SjNu59W2GX82fSVg44KSoNxUD6EpMVb0HWIZ2Oi9F97LLpJS/entNCBSB48u/i4tlVbPISXev
QEK4o3mbW17QEZrUj/EmOQyqf12S5Rev/89VLJP01IL8Nwf4Dmfn+Npu10WC68Qj85JFiuQnmLTt
oarXJ4n1y7bHdqzUOszijaFM8zk9LfXTDR6PcrQesVHVlQWIPkFpj1nhW6buBqhlOZdB/gMCePN5
u/RAsNjOeSY/Pq632GJpCoSkvOH8EuoQdu2JHFnrtjfj4I3RmY3eKegpHczoBup+qhmteZy1BjH9
BpuFqCDqiZO0fUZFJ6mAcTcg/TsDQUQ+x1A3K+KHCWOi5PkhuT1d7q6gr8xJTp23voOxOq5rioSH
VIMcC3jMK45Dz5nUvaKGOVFolu0b+Lz3MNEGh4ASvmrREmaqE9d24SDE2AFCSrm7LEgVUhudcjzj
/uCbeMWBFW3HJpy/VGgMBXnf9KK6A0KHgaGlyAIG38j0Eh24YXn8oITP6mAIqnsfNEnlHXht7S3o
3O5WrA5w5rgLE2aCUzljxBOQsxzd3T11pT1GzxyPgGFP44DzS21oQNyJUZU2O9dH8zWbbhxRl7Im
1cFX21rFcDdUkKNdgssUWs+UI5oPbiHBS/BfLEZpyap+w41BaH2yHLj5oNUKRkES/m9R2YHMPlM8
n5CPa0fb/uhZ6vb5Y0UG51059PK8+aBA1KWIlFG4ZTL7FfiFLyXOR+hVDLrP3jP6U/ARM7qCKN8T
UC9HLi9Ka99VjRM8MsQec+1Tifc6F2nsYbGi+OjNX6H0XZ70ntV2k/SpebFMQd+0UCq7jUBpPbBk
w14s49ox/TjXQNnNJJxnpZIdcvwK8BTnZSgr9fLbVLfgDDdbYjkWc/yyV7Bs3fGln/Q9cyUHzJ+L
zBogrWREzxSrIL9rxKgG+NjuNaP0dCHMBh+vnl00I3ppcGQUvk+57v+vkP7NYrfEpOcT1wgACUh2
CFaXRo5vBLB+3yOO8PlKPxF8d5NUSLa/S+a0vfSNKNOs+rc+akNra2OruIwfp2Qol31QLDqUWurx
h0cyyeuXJpfY8cqeCk9ho7BZh3dvF3gcSDfRJ7TbZi+SDlxI/hFPiwK15aeL7wSCW1mNIvRWJ6jk
ssqyYZQaZm8XWJzpCPSbuSKHt1U/Z03ZjATMtPN4VrfpPKnqVaWRyoy6stmBrczNbWSGhl3ZGUeZ
Hy2VJDWbYyDLtwIEO16XYqUw8kb++C9ktMTCQ0kTvELPucoZ6oW1zp1qxqzlgT+cZy1a1xinGOEX
2z+oGMdDPKFJQDN5rxthnv6TK1jKmdYDJIddIXtu+ca/tsGBofxz/lpyVXz/oz1if3xhi//5DTB0
lFxOFdieWFItpWlqBHmwbsCRVyXiCY4Tb2GK2fi85Nyjngt4UP0XNv2Ccr0H/6UU6kTUyDX/ooZC
6uLWXueA49fRoXi1Ayz3KlWzxb2tPavPlCFC7d20XD2t76t59PwdU838ot8dNY0xGNTNrHOZZLFN
0doEmPYTnyYt6M0tqFoO44T1zUJGAUCBozgDfiJ+hbXemQ3wsjgLPzfjET3KDF8VIb4N4zTkaCzT
81jJpvimHqtKtfiYMVIuM0gHe+EAPW60+yWUa1T0LVVEeR3b6X6h1cNmuSUixYgqibjxfmho/05r
dt0D0RiIpugYER/WM/NEC8ttRwn3p9a25guOYjuLfaBU1nL8i74oTNt4M7Tj8YGiuA8BRt/eetTs
Jd+ujXdwJkO1fPJYUqffrxsjesxbg7k1SwFdyeXYtqZ8j8QBwr8dPwo2bp6JtEgfMPkhA5C9ZIQE
p4gfifd0ynpByymTm/eKsrmsEE0+pjM/LpcHJ1opH4giTiVKZo1MBKY7X4g9/TYPDtXQnKFUX1tC
nbeXuyzUR9JGKptZ7Prpcw5eVte3/kZdKS4JK0xQN/XFE6ncwfDEM0vcT46fmwnvxz4cDcwqapZp
5EfDWYwJGD4LCs8KyjjOHh6ZcFmMb8AcFj/+v36L646Pm/PbJxIVGOt/kgq4dqyVi0Z3Y8A01Odr
3c8DgDJM3gdxbhImZz6mWrVZj3NjP46zEk58aocB4QPc6RZ9DO1o3GFPwHCEXT4BUSvXoFd2iGnH
Y/AM39k5tgWVTe0k5iUzNSr3Blmbf+e+y9DGrKiQHFluQZDU4QsgKix/cxqfgwFP2zB1EZK0e+C2
zz5abzWPk+EMWZidzdSqY0EmpH3N6HMdzPjVn+XX9xsZML+oEf2y/xZSHTb8Co6vpL9rKuVeH6j0
6ZrLsnb38Gkqo57iRw4nvOXG7OJxgpWTu7TY1y3HeDjl4Rl5gOMUnf1tAbQ1tl1W8wg18V+Fv0z1
XERSfQ9YWfBQD1Rr6W4cPj36atrv2YRGPgZUIt+FRSRmwbhpnfW9C4ZDbVgKfKiT/vS25nFfh3Wk
Hi/M95+evNpft0ZPNgxahCevfjD+XwrPoISdxq4e35POvFJSZDcdzlW/oCvboky1OKAIOXcdlZJk
F7JsNdTBnuHa7lop7VoRXmTmaxLo8KJaL6U2L35w8vqN4QY6Jm/rDJ+kNvrzhxMEzHl+Jb+G+yj8
NYwNozfIJjCAcoM0tNxB1jfVplGJ9QHDaLfTCLuvpjeVbMdni0gYPNmWjvKj7qjHf71Cvemb9ZJ8
TBbSh6g79B+1DWn817KXG2JhuoeCKAXqLcIVbYs3/Gx/nsc46tgxIcSCAgFq95z0ZIrT1v5AjS+u
pyyN5mK44YYw6y/GFC4B2NacZEU9kN9jOl9+kgtrd3uuCgYK0dxuv7UrsCfXeD7VUHkJujztlx5x
Y5wVomTXkp02Fe546jE8MnQOEL9rYtYf1Nt8qWfqUqV02GuY3kEiByQhTqCGJBpOqOlHWWxzsmEH
M5mbxH5NDMccElm49UC7H+EciHemyCjEjVw+o4HrDAro+IyN4FwVaX1IsaMBNtY5T1cuF4Xt5eYH
xIBYwITWYVGJ5HQhFn+mSWiyEWB7yA/8cegvKFzyHG+jqvqb+rX+tdrwkENtJ3tzMgdx/aWV6Vay
31/ajVbHlCuf2XD+99T1uB+AFm4D0AQGtujaDzF2w99pfo4QJ4ETMN3Y9hg/bo1EVsbODHrWBblv
DIqr/fYjnjlIBH8JXdSfkftR2f4YudZx0Gv75UF5CisfZ0vjQLF2rEwSUX1pZMCQj8SfeRNIVowj
nDx+bGAjgwINE3puyWDIjqA6TYRtdbh3hxAKLiAXsSAbSRuP0pfpjYt30GXdfD2WnS7kS8bOId2f
/3u7iai7yGY+P17rUhxHi1+04Xrf3+nbly3XLSrHOY+QB/D5EK7U6ntRJi8G+JttJ30tT3pO656E
Uy54YYKHsuveZeW7aA7mkiTRPsmDQncjSY0uDnCsajUYJd26wFUBZpCFJ8PECeN3EO2cf0QXE5Mm
P9jJSRzPT9dFz0QJB1pfCvaVkvvaH6G39V0dPFcSmPkgG9q+QtNBOlyScJJiIQoJfGrFjsXQ4hDF
0L38VnFkgSi/GFcYgW4OrejEf4CtZEetswFCjNDyJLiLPH0J0BiUNweiLph3z6NktFt1YmoBfd+2
u+5ghIyoDnccx60/Nw5cZmn3TYnEDa2MKsF7Sdd8RNyXkcTh8FeJJXdkvDaBsMvB1er4tfgpFOYp
1g/GOffCw84v4diozyZhS5tDUSgMxOKndh2hpVofFpwI3b7qBHrNaz78Sri01wWiVgA7B1vMSaHB
nK1OJ+RMhKHnZV4FAWo59PuAFfOjYSYR9eSu9XnpW0hBmRT0eXjSkdmVrqV7norz2A8mcmx+emQR
BVJ5xqGUmWE4OIE80lQVdEotPDUdqMU51Yjr44pMkVCrHcgSB5KTt98WpZZKVvCPAWcayGt6gb22
HVM4UMhufrrih1kjTBoZl9/N/Ao6s64F62mX5rbLV5nE2UD6PQnxJ2IWeDryvqq3bUvjNYQauXeu
vzg6KXf+A/K6O9U6gvPBiXYw2vuvgVeQRmEMTwogNaw2OJZQqMbwRKk9CsTztm3nrKQRU6xwHePa
KSrN7mti2TAEyi7YW95DnsMXxsjWxFdCRLMTpaMt/L6+Gxdq1OIjYgxITxuMO4Gq1eBRpIMT3Q+u
NnG8mNHZLWBL2vTXYZvQ7LDN5psj6HhiHxhtTyfOnKozdhE7YA73zp8f7dMkxGn4nISmBpmFgell
mg+G8D9zqdzA9NX9vjeqwIBvcpEDuBJubA1dyWPQRWmXbwbP5OOnV3+0gwNlBcTVh5nUk4W8BJH5
7Tdh+EhTqkru+k2GoZr9jtoHK5AKJu+CrgzoStLm1/nwOUdkSM8/9dft9Kp/OuSIo0GvD41OYOrW
0GF6fbiVKX+SJY8V3M8e2zOL6z4dJLq74KiANAkaOhXodSQIc6v/tnGcb7rBs42AExBdwLZ71z5t
BN5Q7AhzQwjgZrRoqQ1seQ7KZGACcZiU3Hz1bZNQZHYDcn9Z/DL00evZECZ7mMrfNGLTyDtV60cI
mEPnwY/46n2YobPfMjV82FmDWTUC0WrWyUCKzR/ekCNjFoQpBAt9KPTJzsBeGAE+6iiQSG5JZms5
y2E2oml0R7Hriku5Y6iG3OZ1QtYZPBHJy0Kn9gM2DQQ7PtqeeF/+5wW6LDsTDJ6fcqZtjN6b8eRw
sXQjMRdLJNtWychm1hnZ0MZAbJExh4k8O3wYRyDL27Yp1lzQb6l0HvKWI8jMJFblCluVL9kwOUhz
hlvU3mbTmYH7TvtGBoMG9l6v3D6HrbJm6urT02v4PbO0/w0GLptiyajfYkwpuHjf42dNMnUYnsY8
MdtrJO8xf2qplVrgafjwmxdNAsjBf6It1zTkx/RPrbCMji3jkrxr8x/Oi0RyiH2hyNJDwxFmqVv0
+9ecjVWSD0Fb+gtWpZg1+q8ZYWmAJKLVQgiKhqBOC7/JZmGTogoYMNHAvNg8kQ9zKpaE/ENtHE5+
89MZpwd/x6nbXFsK/iXzKnhyqpSwNhvjWvJqMUzmTj8OgpEEpR/D1CiL/6VXbM6VKSEFGENtWil8
T7EM35qNdFs7FJMw1cU7uq2PKbOvQexD8lWcXP3O6vG1C4nAHdQLvT/6/8AKRSs3s/ABQKVHQ2Yr
89SNEsJvNz43RULsyKlD9ntiir+t0PhoG4FmLyQnrtbwYjgdUUAtGxDotjhNfpk4dq/YQvlkCFPP
s4esYRAeInUH4NNBnprNmjCqDYfvnn+fsKC48ylgvvkzBHT+mZ9Xtmk2gQBp9GDPq13A+NhXuAmm
u9QzhIDl49cb25M9RUiZet3HcgEzgqAQpiQyTzQGyYSvACXQ2kaN4fqNg7mxnjS86iyFpr7vxn1H
tVedejpGO+iMSb4P0lINh4FcSFudw/+oUbJEkbq7tUt8u7kkqZ8f1p3IHsdJVWwAvWCTcAVUpMYo
jqRw94XmaPOS3skfDtvovOOJryJQfC3sAPbB3vITCvcZ/XxzYLfG6E+gaddCQG5Hq5qjBSLVgyMf
TLMCEuo6AfzJexTpuTThhB/AyJq+AGuW0mkP4XatlaBUBJWaVSQ5HkgTVGeFFbbXsSUTvgPjoc3B
2cG0wjghXo8ztT7OgaGmu8CoQgqptmmwaarI7l5AodtjRXqhoEHQMLC6auub1JPMq3DZtHGl791Y
GnVDollE/kQ9Z3N4sxNaejwpJbVmnNVs8qjRimcf/KnTOSZpIg2/y6SWf2AeZqtSHrpxFtnlUm6e
BjxoamGHyk6Ek8jkVP4jUjyvtBSx9tcyKycVLb8eIYRo7W0M6PC1oLKldqXkb2HSMmRpBtBFlaNm
Be9PvUqHmCtIwXG3cQHCzy0xQQEBy+PQJIPBNLeVsMTLCSZ0KT2RSHK0scHIzqFWooebCsuE9hu7
ZmRZD2OlCfcG/wjFXNLbkwIi3bFylYJ0q/l1fy+2iWK0GOJ/aZcCys5rRhnGxFQWPwRdjoxRnEsq
iYqR+he3qQqvgozB3V3+4B1oeGvdxtX358gXHuNfprK9pzQ85UDEFmrB3fSQdG4HWh0B6i51QDLw
VVD9Rcmj5F33MbAOVUtDXQBiwMcaJOvbCoUdHt0Q/g1jM9OwIZ4FjnCn/tz/l0oWB6o4J4CLfFKx
66adSHpGH0CGC4QOGrTRkgG8nxQ50MGC4TnVL8QSQqFqRcsckhBZE3LiUgORECHZkr0n+FfMozUZ
Vw7uVvVsNtPlAspu4fHvbo8iCq4n+9sFmOmbaGQaubWXwjc45GjKLwRVPN5WoYo/eMMPbeGth314
KmobEbOjZaL1/j3bbWMngUaXnKSY8ThIKJftMgAmT2T01QjwfljDUZoIyF/EQvi1u/SIu8+2bhWL
nfpwbipfcCqx5rofA5tynRQpsk2H8++yXyL+liSF/BwyrRFvN1UPo9rWTwLzZX+fodUJwYHn81pw
2b0XJSVu7njfgRB4Isa7sj3iJHzm0o7o4yiG4fjNdCVnOVmQ4g8iL49s86wZHsVxkT9WNktU9tct
qtLLkpfbSsMW00xGNqA5oLtdBThlfEfuhrDgq1oz2okSB7JzqrtFck2VeiPDGwQ/Ue7hifH8pmYj
GuTeSnQ/To2Lf6liSCio67mttmXddnVeWzEhrw2dMx2xuuTAedUDRfHQMFdrwTK8yy3Hv4+3RqTp
cfkhUeNNPZYbXz7RrCTpQpSCfRkiSFBp5TRp9culettiTLX95YpXnVu8KrYX1Lj8Eix5+DBOS/2x
ffL4+dcxsADC/Q1sQTroKkujn4uPLR9j1XOjMJMBYETcYBIK8k6cXh3Qj6vxFvT/pByLdWm4CotO
xkuCBwLG70esmngaNHWQtKP9eBNu6jNHEOxOuZQOordBrAXrB0SbzS+ARTsQoMifw614jJ7O2GBG
Jq+11BfjpCwgioqytqr0N3r3+gxe68LGe6DJaN9Dts/eWjckReQQB4BmwKY+Cs2tV1czY1j+E/IE
tEeBIaFS64zh/r90qbVA67GMjXpF7j+KjG9Zx1S5FnIoccqWVpDjjJz/Ibqpolu/qImvqyv92rq3
HBI8bepgsS+1dcZg9mYVhj+YEubFdKBTUkcvsULBgaAjZmyIKUCoNQmmhH+Mn88LhLyhqgEHwcOQ
SvnWwqsUnb66tfmtapSFcB4oknXn9DzfuuEl+xD45/NfeST62AJqMEjR7aALTgtAfKNhlkWvlPPJ
fr/8IO5zCkRR0vnJZhukuYv5xoe3Kr++5xNHyKALCVwTKAzYihfJ1MjggSUGUnzJ4xyEwM1yKNU1
/5D/3d3vQTFpflExO83661JH3NlioVGbn2znSxLzRwJ1ELdw+MdTXU1EQKzAWR/e3lYOykNaHj6q
dB48tgX6EzfydoXQkiigA1zaPpVxJGTfm8UT+rBz7s46F9Bxof8CigZsW5sIVJkNza3o5oniAq2p
jFtKwYsV/dXJCXDYCNk7qYw0FtLhLYapjO9PgCgxyKK7hIwYnf2gh8D38kKTx7Ixdk+289TxruLw
Frc5jMlfIwlZvekvwJzyha+/050i3fYFWVxnQlu9n0dkPk/rWqrl+VApvwE+JobjcXOLnXcHx4Ch
/mNTm02YMl6qzZ7kEL2exeRCXDy5hREizStRmLvMoEHl9B2atyakl9cEG4Wqa9uMhhNhpG9veaqu
W2YVYp1qtSa+UbOuEOj94Eu8iVzxK9g8u1Y3ukNn2LcQImj7dESXiNm7+lO2u+eKHiMZZpUges3T
46C9U51KRRp6Nltky1Z/+wp2LYEqHSBs0Lo3LULYXNaFfRlO6BgdVHAUs3c/tUyGsza0RKf5IoW2
QIIewTBAZeYmqqGHmykwhvHofrdQt/+qnbqD1+bgWNgi11xY+ubiJEJNAgFDaSBYqK98Lys/t6RL
CivtUk9LmOdSszpNqlgCkxL4LQs7/h4mKLCyRdJM40ak3f8OzDa1NahNBYikd34vMphQNibrykTr
RYw4i30mrxH838rUkk3WQdHjTCmTL5DEda6dv70LDZZ7BWjNiTgmJcHp++neyL6QhGEzkZUJrRDm
Z3s7OMm8X4mHK1sPhrP4SQcYF8AEKk6Op/OGl74TBoOsgOhwXkUTG0DhEbsECmSDx8yWiYiP81V7
YNMAN2KjBhwpFEAE0cP79mOm3wCTtILiJHAuQpvWeI+uSGmfVXcOfcqhljrBSa0KmH+3hJIEbrP5
sge8w6klXlmZJg+z9iOh3+hMTkQ+UlSpQBnXaiSSYOKlcaBpkbFTLh95ADJtD3j2hV22/c7DPsPC
sdr2/K6PQRhyf9ppkgPzNs36PJJCoHCyKwVVuOK/ERW6FYBQxRWGTF4qoLjVMGnVRCkWNJsCFn/o
Dv9LFiMYUOPlv3xXsWacfatnUvo/3g78JtKwP118gw/8XiCl37p2623XCzH7xuyzHtsbpL/ITbRv
DqlrGTLbHHd/TIHl+tzgirLl3XKRbJoQSVAHfIhKwZ+uLtJd2RafZriw1A+6k8cYwUT+fTAGtA0+
yOQNw9ZL6Rm1URXckb85sPVfikjArGe+MSAxmZ/nuzQRpI+DCFizgPA887kI5BEFsUYwiZnNcy+T
N7lFt3UyuM/ngFh0pNbaKsqwPg3e9WziL07tJwdFCajPXBrT4w+yySCd9eWp2Hu8VbcNYX7cv566
MokGJJxP3oFiewxONSg4SWABHK3KSSPYB4tZcVyE6V4XBnlObg0lomfyqm75ntBliPnXolFn7dyO
YPn8Hw7NLT6oMArF4u3Ak2M985tbdHN5SwsoSpIfBZGB1FFh+hPdBQYWnjeMmdYwEsjd/rINnwUg
Jy1t0R53o3xWJz5SbqrW6cnpKQUk1FV6U9WMPrEWlI/dJyr9ugxfM8rET50dLFoHfTBnqostAMkc
yXXZl8GigvfmtnHGJ4dihGnjM+n3SeyciYpWERRxrb+iOrqS9BJsVWJX0m9ORpX/gxKd8HlBYTof
66+bFhOmCJ0YPquthWGyDEk/YYZQSYWxTtmCUCB/P3RP5Uj9OG5/WGr/cwO1SHS1Vzdm2ETwRdpe
bDxaUb+MEAeCqCqes2ECUie7BjPRXpRXCR+KRVZJPuyvffDYkj8NMlVXgXdDm6eX1mhmWmIFkgVB
3V49H3CVeJMs1PZMDp6k+/LpQuprWn0z/jtj3RURgG+Jjnz3qAaWVQmTSpltf9t0QYLje+Q5vM7d
u0tUDIy/g/BU2JS8XTPCskghk+tq4kVVfg28m/ov8wbai0FpE/E8R98/Fvagg4lOu4RPMo7RL5CN
+K5U4o2naFUUlFklMYHPvNxT5bV6U3cFc9kqssilFoG5cLa4c6JMPYSjgfgTuh6qzQMaxKfGC7qH
TElMKZRpRw+sTCMZv6veRkAmplJVPkOr177vG200ptnURo7d57SfGimXWe9zg3+FtB78s8PufVUd
LvMCf9vIwumycs3OOyVoBSdsbimc/BlSC7x44iMir45tA6xL2W8zyqW5Bp2Wa9fzgcwDB1/wFg6e
8gOKRbOgIVcvWfvPnOcYTDcZWzgg6KJtwatG++hHTzcmVoRxdsmbMi73VUUX929ImeqWSRmwqXZ0
okNfdwK2r2APdfEulopeO6D1gfKbWcD2ETR98PHzjUQERa2fLy+CK9ms9J9BIlgc7yr+n/yLgLn/
YUiYrUvYw9rPqLyHFj8sByJCU260hgAtTAXcsG/zNs9tzT/QtSvlWZujweEYTQBNAvcEBQqD3M0k
jD1B9hGqwV0Uvxw2u/Qa1FHbhZRLM8VYH/kEMVBvNKEOvlkGJEd98mEAbwRLgv7tB02cZFJvjm9m
HmFguMgfTy299AcR2iYXSDgGeMkKB53iIl0IdeiXr9TUxyFkrkKaAl9y6udUy1+wxbf1nZPgvqAK
tnpSAGJ095oGUHGhHLAJZwXaqjhLp2rrCMaj/7hjPq3BlZpNFGxhZfa4pzylMk9CYTGd2LpQYDnv
IVBZne7MFmGFDS9PxyA01zPMPM0yP7x+kr7e3/zq6jV7y7LtCHBVZdQY/fTUKpThTdKVieuNPL6G
Q7kP32n56F3yR5kewFdu98f4HTXe/YwbGPF5biqYYBFf+K6U1T+PKyoAv+XxJGCqbt/ReD+eenHE
xNrZSlCw6Bof9NNa/rqwGQ0AQaW7g8kbrybS/yxVgAvt9s/OjHEs8Y5PD0p+2lXBsTC0p18jbsX6
D6Y9FEg31JD5Ubg9tybEoXdmM2rvCg4hynmnEzGNwbtbtXdfQd6e3twV3/stNTnOtZQpIGhC0RdP
OkLm4OcDQk9DPgaE9ZFKyW6SuMRbDB6KnYQtTnUUgiWeX1SCF4u4IBR9wngw0vUMGCqoLPq2LL33
ZHnV1ZY1hZVjIXtUWeIE0MHCVV4tD1kKQeZMv56YJCO5h1QsrmoJ7/LJ2rQF+HopGovwgSlTZ8JQ
taDZyFTriEsi4NWAjVbgw9iWweFE6G7fIQbwydkssURVzCeq1w3F/GpK9mmAxCr+kfsTT8bOaUSw
2l+ribhcGo0kSUBhS+23v6PAWPc3VSRaA0i1Bc9VN2DVGhSClgMay4CYI8VGYjfIRFVGmipv//3s
WiUKL8jGH3gKToXBgZwxKvO/693kSkPCslXAyk4PrLSchW29mxkijDUUfUdkF+yED2DgFmcgGdaY
40lfMVWYuK7CU6/02jjXTM/touyUwwmrc9ye1aX2el+oJRPXGSmHha3jH+HhQHDv5NV1ICI9t7Ia
feeDrvUXB8Dx2M7EPhSvPT2IOYVmcPYjW9sW9wIo1iH2Wg96sGTVZHoR1Lnu2pPNo+K3vd5HGSeB
h8KruregkReWwwI1Foqp7GKn9v56wCdLx8/VyBcZL/b9EOddYYeNoQOIbI+rvKBw7bZaptU0Wlzh
CxUMaQEmwhprdB/LHYQ6KwJ6sCCPY1AT3nUECxdHbLci8eQerv1jWZHdBKzKWxWmNI7MJ3YFenFz
U8WLt2vuIsJ/wDyXM6eJxjHFGPpQn1jI/Ith4jV7bx7LftD5HPpVlkshOt5Xwig3uy2ax9HOhQAL
iBRJlilKeP3pB/WcFWufZCjg8l3xet5g5CVZjJRxd5Cn5l80pm7Q/UPoNmQ1LUU3Gm+nX01xGLqi
ZPm3hdJ5g0igGLQ6xH2pDNuFBR5JIAHkKhVsxNwpWQFs8eoWI3USacpH9/r4nUCE5G/qXaDzU8yf
+WiEZcmQo58+Zsnac6Bcj+Ayu7VVilz8fFldsL35OEXflPO/gs+gL0YGGiCwfa+vVSP51JofqOQU
xReghh57r7niVjtSp2XCwp6z6zkdb2sdRJ3IUg5gyvxmZUx1wo/gpP8hkp8mny0P1F0++fjlmVXE
EP+k5v+PcjkCLC2Ne8JBCKntTKmWdcO7Sti+piaXqyAQOVv4nu/ovYWRDZbCX1zpyPQCFPGAGhQT
gdAsxq/VDwC9Pb+cMg/XfvgcutKUFLZQmK+8gPRLsfcTKJ0lCRv5mdsgpjwLbQ1ggd/82GIHfBHP
Q9ZFSQU7kHkyT6j02NHGcy9T9GAArcw1cX5Y7Sc/mq7xbzL9kaIn89oXZV9cc3AtZPZFzDya1T68
OiWOW9oKkd3YEmvhBwx2SS8Oxj5sPUAlz4WtO7AWF5kwi7pCTah4DgNGEXekRZxxgl72nvMhnk31
IeOYLplOCIRLiRsjVKCy1mkFf+s+uFQhPxiGZiY5YAYTeyQe5tWPYLQTeLkhUjjXyZrHymPVbd3+
4yC07uN/T3udRvHY4bA9XTIL3q0f3nxOUa9UbNokXVl/PARFkcUWtssXFmU6Bi2issh3tTR2YwwT
TQLaAL/Cv4unjFlSfwHqYLHPhLHvzx2IMctRzj+oXg+EutCx2qw7eUhlOsbNxYpEYUu3IuskT4cx
pJtkLHfUWQJX0qBZ6WHaf3zUdIrNoH07zPUJ4PEwm2lkCiAbhDyjbiO657wkqNXgCZvtyVzQYhmD
h5F3ssewoXaLBIaw55F0ndp6jiipK8TVQ6/PeTZVxlGljW1HR3JzEF9tEb4DhnvI0OFgKJF69ugf
ChjTCrJaVZsugrkwEMui+RKmFjMEh2PKxfZ0emPIkWokJ7W+jffLPYeJLAog6I6uajLvOah3DYL7
A4qeD93dfaFdFeFU9rzT/d96/n8o9aVbVFnhT2km+i3uLhOFg4+3v2Jjk4rUdoxGx21YGEGfiBTu
WvPu5dqYYZjf+je5ueZzgw95z4vs9Qch141OyFWlSr/UYIxMPSDzm2WwTgPp0JaTzyXbwgsfZhvG
j8DjekXqkU0RQhWl1Bp/P+9kitTeH3yYYx0KlMbRMBqGSi38XzK/3uZNXssm7mxjRxYClswBdChN
0VyygykEh2/eMy4tTX0NIJ1HO3l8MRNxBwlEE6erLb/PNY7vSlvSp+UBKJvl/AF3R1K6/VOablfX
DAm4b8RzcrUIKYEuyUBr7HVKamB04SnzrTmj7GyRtEtQn891YkVXQG0TzTtDdfIzFNPr+qsB1H+b
YHohPxMb+Yuid2WTx5XbFB4yYRbQyeeAZyWrDYBZIGVdR8KjIeyYbLOdiWB5b+hU5ngJQQ5IzyMu
yxj8Agbrw2BkxmCMPfyhVklsnX5m4MzajpT5ZD902ZwhPN5xbCz0/v7HPXBUXfACnkjVdNjpl2lP
EE1RgmX02bBtRmbWL2MBZ8C3sc+TMpwzTFbTMDUGBH0sKspJc87ER+hl7iBnlPKG0vMl8m/xOfjZ
X0Bd+9f9jQW+3K7bKGUs1VxtukuWFytffaeqZ/Ioe12Ds3QnFm8XodZ9yZSKXMsWm6PavbTRlZje
gP+mSSQ4HcuBY2gA+pb+/HXC9varzu39dI57GWV2CMUfkB9fnHO9C0YR9F8Zj2upPHWgZ/8HpAYi
i+ywKqL8BQ4vofYlyqozcpHaoGfnRYA1soXRe7UujrOXZsi4StFbc/yb8Ozx2KCO4cKdFpnzOj/i
d/MnPR24TlgUiXr7kSAdGGc6OBst3PEXpZ3d7VmhGVmW4ddCo6Jfuj+fTSJ02y3Kyx8Teab8ZzpR
YDsCljsqQiXNQJ+cBeOxfTXm6bCNz4KhQS6S0fWKHewZeAUDzfN4BGbQM3lywmqvEIGOs6MZ8TIL
0ZVPqLsQVAHuL0gGXayjxrWBlfkZ6I7F7g6P0AtPf2pcNAjxk8Hjy5+6bWzGV7+32zZ7f55V88qu
G2UPm0ia3m79LRtkXY/FAiXwzUbBDLLM4IZAIEg+jvtjkqbuU9KnpjwJNAHvSYQpA+KeNzHMNh/q
02glVjF+ImvbOPxbPwAcfxYxDWetXJi3rk6KgbcvH6XVDCJBxQPu+uBITbC/SrD+0LeAI0wH2UA+
2X8IQ4VHZpNV/3PfmHEiePZFkx/fYtKDy9bW+rlKiH8Cggl7g6U1n2I7oEh+bzJSxMchS369VTXo
pzlTIp3FLaCaSnEthi/aDDCv4D/pbpCtqUMKxV5dMMummCPN+xvo4cA3BOBQUB9uk59cU6OnXcD/
d0bomVYxDPhfnYQQQ8ied7AEZa0/KBW7RzeCK4K0ebsBdsc5mQx+4JMfnlyxML/HoXMJ0RAdf4NV
vJwGBjqUzuUWcxNXu6yhdZ5ZLo//ZzhNi77ml3qUFsLDFBtdnA8+TEhJ/hbxFCXWvMpGOjkRr0o7
h6qHStsHE9HyejZtQrZgDYvKi4eHlYwKiAz9wdkTptlSpwZjGVrSIKuzXfQrXAEpf7d/HQgvAzuQ
u27wRH1rZrEx4dh5uj5c2IjkrXq6691EIQExvFexIBapaEUiPUEt9O5XvtjBqnccPsdyIt8gzg9+
1B37kHkcix6GRRgORja0EjlWYbyl4HwGuVRpnqFON7YqC+DQSQasrD/DGNyirQCgBdj7qFECs9VI
bt59HXFa/1eHzG7XfQrOoulGvfQnhzd7Lk/iIJ97BRloRtix2629lzI8dtoKffb8Hg5FEGW8d8F9
RaHEM/ILjtCHA+HjBk268dQ74w92JkmLj8IvsHyinJTuiTUoupluALoWwRKF9FUEWx19/zeyTeZN
WlXHcSzLmel0ETSundkEltMJbO/X9h94jdoJ+p/b/phU7QK2P5rnFdsuInMSuMDHIZxRO2xg69h7
lMu0gcLGYRxurhFXDkD1cG5+AGYJBIMX9Itctb8eFC+e884rM8+z2b5b9hxdlLH6OtWukjrFttxe
XOqwq8ymSSf24pzSHoPJK6YjzsYfGDpyf5TyMSWZwKK297/httkhku/IIDsRA6eMcA3hRCdN+d5s
ykJ7O3Q6OmgRQMwF7mTEmbTQkF1kmuJUlEimKz8MBfxV7pmxxZIx5STMKw6IZuDUpunHin5thJYC
De6WaCN9SyNhAIzr5O9q3UgbvcAk0y3/Jcvj8gwQJuI6iQwmgmA9jh3syELfoXxdD44P0ck/EmGW
QU8YglJobFXx0QXgy4Abj/3rKCJayKzk40Of+CaCYMz7zEQaiMZfjg8rVG4Q2KXVmLl3CAsI7zGG
ZzrzwUMkyMnJBtOi2clH99fNMB1XEs+0OG+8XvUHXGGFLhE+Cf9iUH5QsXMyN9COPmFv3U5vS6yO
7o4twAksSVBDaI2ev73SEyyRhS61Nwaz4ywALsCGnD/vJoCRGsJOtGzBE+12n1wa6tvvabkpdO8h
baO9TAxbNyGcjU28qUKp1buUZIipTgNtAuj3mDmiPUYU7V5ax7svQwYKwR3kIDebhIC8beQw9Eyt
ZeefO09hTSVvWctAooxVs6TI9bB0DCPEupHLewGRm7K9jp+UYGIh9YjQR4MWBXryz+F9MyWAfb6Y
ckbFH7K6y5aqMHZimoHBxSRLi5tgnkwaGe1RdeLqaUA1771897hp7R+cLjxjr27UrDwikxb4PO2X
2qYt9jV/Eumrxg8xVjl+GbdoVnU11GKECJg1jBtb3gJEZUzr/bM2CnKMOl25M4NvkZMdZkWU4v8t
8W7ZofwIZtcuw0KpsFU9yPsZz3R26VphBZyLBxy2txB5T1HcEiBuBNMdVIq5Y1aoOCoJOeZV6/RS
futDZv5BLMdobq/nZj3hskWX3fEi87sMmF2SGoDjGA/+t7X9sdP1dj6fxT3GIzvdGTz/dpmiB6Lu
fi9BIoRlCdRF2n6A9iL3y02/JZapo5knXLgymDoJl1d95l1In4A+24f86nneXWEkhRHRhvpZ27Ad
44ZpmdwT9BXYsikSxwUCSUca2GjzDjtXd0oaMjwwZEzSdUMfuvwDh68mEdqwtqaN3SsM+G45ff9H
76pHEYs19heR+PNBAg6xiJrMwKuEmm6v+XISGFM3+M0Glb0gGya2Ecf4lHclwC5iTm+5AJaVzPwf
z8Qal/9+30kZdJ4ax6FUX1TteXVkHGwgxNTXD/QGN/AocNVsy6s5StJ0nRu5885qETPYL6h9jnSD
r8vel8M4PfodcX0kmilUtvma2//szNdRcbb9w/092X0qGTUumep1SZMl4odmjm4H5Txi1qgyLhCT
rOxBdEAVQhObjAEfm0wKtTv/hCkC89Z8WYacCyewjkCG2VqjR+JI8BH7d0e2iyGtSi8DPOFQqHNI
BEJWwDYfduAAzEgZLo+eNUrtZzfp34cv2Q7ASGY7gYKPKCGpkoi36k/5uozu2ttEDPZgFm+WXfbT
fN/8xzmCbY7jA+5rKsqxYS4s/gUjhVh8Lzi4qvterULO54NcMZHOD6Ul0satiBDNGIrS2WSDlmiA
WB3Vtnqdd5DUcPrFFwveJbwBzatZB6xtoKLlI/8tFBE5e5L5KcookALxxJdEWcMYT9FyjBA8cobH
acdTTYcpyNlXKz9Ew1HlZbRTRjXrzcY33jNX9al1aEDgrpIO/xuQhJ0eabvdIaHEc0L2hC1zJmB1
rhL3QRG42fWcnVhiDKFcKFcPkwSrYctksbxgd/NTonv9shdRHSupH/sTk6MqNR5n5xI4VcorpebK
Q6IbsOflEas9404Jallu+1zmknu8178kvOa5LHkxEi5B2I7/3+VJjskAEBHTvu6GwvNaIix0cAQ6
Y/DHdR/QgMgnPieK6PpErtIEtV4gAbJz/jT0ZqcRKz96FbZHQ1BxxIne+IwTZ24d6WCQRia6Udkp
aZ9ZSCy+b5VdMby/PJmdbk/uxzRf7qiykj+8uMhVZR0nSd2zJghthWMOd94hzOxc/rg2bDCNFUYK
KhXscLnnoqjjAhDZbI06vsuwGGJluOtbXdWN/JqfNbTWdO8Qu7pcRQtM2TFelKosYuw7kq1LnMVX
rmDu3GW4vX3h3jO1Hi9ZHWeIcU0qRz7XPlL2GHgGODa5gMdrnVV4CQxq6oouj0U2m9+ewwM1egva
9bupyB5yp7HU4roD3xZ6hf/dY+cw7JyuXnxsg3UscpFSjsm7+jDK+VaLlQXlFwmvvdNow8IpEa9y
YrCMyaG08o2imjTAXBRdowKpbj0AonrEkjAHxTLp7wuqx19iapzYp520M4pxmgTsO3e99v37NjEe
Ke9X2mDgNkIPhMTp6nKQqEEKDI28HoUKW8mLpRsG/PbtVSCrgIGM2Qsh+7V63axe5AtNOAUv9m/I
KXX/8sr0nhOwkALIH+IhbZwelpXrmySgEToF3D108hkJ0P+XTg4A2AxYUwemcYYBT+0KHj3b7tCO
h9zjpSWtZv/1iLTTy1Ic9Td4Ii0nco7hc6QvMSEhilDEnrHfsnU5LIE9hX5SEILFoFuXppK89tbQ
mBBaKZMBSCFQ3zP2NPyBLFhr8JzAf3lWuhV+XJ6GmnOz8glS/+bUD3M3WxUxcpNE2Jpfej1gVNKE
2SzYHYIGGyzDksbFMb1ulnJP9G3v0pLvq+bWWNGH5ChLOISvLiCx/9Hih/pBaa7H+0+1mwGjbwD/
oS9yQt82QqGdTlyRna0jNkCIRRLcCVaFGjFhhdraZYDjTE5OKou2FxhwlWavuPcJ1j1CHiZjjQcF
abfPabMmdG/13vrO6fOMjS4uniiR+iZCQ9RKzS4v7tAhaplZlNu0P7pUgbQRERinI2ySjvBq71Pn
fOTmGjehI7Bob6WPU8vsEW/Y0pd0ol0+58VdiMouRhvQQgK5ZHTsH79WD3PILe6S+UfPPj4WUqjJ
xDmK9F72KtyNdxJDyCW5oPybnqgahARXWIzcHG3oi7xsD/i7FgrGumc830FqX37cpKVKAx0dsEjq
Tse9uJmf+7y6a4bG2uxXT2gkJqUDRewCar0AGLWinVnCM/334crOMa4LLhxibKXvX8Moc87vCHTn
r5rhWzee3z616pbNYDbPNg/PE2lVz5S9bENfeDRHsBJy/6kBnm/vo+POjbT0DXTI0x1doQUTVzyi
83uv9m5t0csATXo2wZgu7MC+UkHvcLJjcBV5M5U452Khk/jO00jMDl78k2IEtGeTY22T9Pj9EeOL
WFJDQi32cpdBpm79vQhco7vDc9JCkGbCSS9eXSIQX1bZKWjjdWgeTHk5LAyL05bOyq9o+M8mBgvG
pWYLmOeCe+2VdNdbTXgp4zkHlU74zNgGdJYdXi1y47UJABdjrQ2ZqIsroH2azlwSHGViffAWyzs4
GA/C0TuZDRTWYcQOxXe6wtjis7RfyjKQMvGburJd6J8CjWrwUEYb2BHYiaitpJJIW/DcDQw9MVh5
7r3C2SWIm9ccjEyrq/LCKRXspehE8nEVPYsEui37Hng5judo51/XJx5sjb5D01DSGidvMlLphTbi
dFyaqwyz4vGZyWm3+PGUCGCSBaS9KJdvLWV3EwCV6PlTfejatOiMsYyGlJ6GWG5mQP+i6r4EWyno
46qP6BxjIoi2hEBwlyYX5x0o4VXwAdAgwXeuUUlV7tHMnh+DKXBSy0L5rnJfmGQPEyfVKSfnWCt8
H0iSrytVhJlXRVR6S0h4PNnsYxk6zD/QUZRxDKpR3YAT5kMwGg1BhMsbAWIIKxUHMiJXe5+sPf+N
PuVstbMTpOwlBHK73dKbnDdn0ykJL8rOIi4kToio3HITjvwMve8z9W5v0uL9kBArT4L+fCznEMoF
MGeSnS9B1gpFEjNYqLcXickf6c3Av05h/JMn09eHJkkc20H3EZB6NnWToYXA1o0LCIKN+s0p4PVW
GKLkQQT6CRFhOp/b94NeG99TKzkEhXSllf+KtmWumFkLhXjzavrUo/8sbq90wtNOoR/zDZXsV8O+
dbWrsnDwqosKOPB1L6uFat5GK0k1QBcIg8HUfh5rh1ujKxXEHr+qow4vtNqYSewT+Osvb0eedkAD
IxUdStzSuQO5MZBpfGhNmx1QjpleA1fOSKj8tZkirxMBR+6jzqqQB236eUiF4GrUsvdc1v5+kUxy
5O6wrlknL5pPaqBDU5cFHi6q9BvvzgTCPhL1vVtK7I+i1J3j2XJHzXVcr2msq9jnIa9Ko5nIeGMI
C5oNF/IOGxCIuBc0UoRUDBfh0FJCpHbUBS8/apf8yr1he0m+RFAr0ByaeNoTpDiUMkzLdZwrk8er
dhqy1WQhLTrlrIL9Sa6TQmQWsCeinM1h8/JOACxsclfo7xoLQMgkXw/AJCcOkMViQiz7b+9yngLn
59sk52SsCq5bICfBvWl1mMJXwrtckQc6PiHO2L+PICeTQn84qGBJpreHM+UFnUP615wPOYIAB4lo
5kO95y6oywnlbsV+ASm+gyu3MvmWAG8vSXuBZbgmEtMMQn/2E8J3teS1BG16j3PUlG8diooTvqEr
CfMGMD+vI9Eg51XT4BJqSP6Iv0jLfCVcaBuwbWOXzEJPaJIeHpMTn6R2x+ywLx8ldlJml1aJFesx
QA2ByGs9ufYddqlTax8MwqBimKrYXo89jI+vTFaGRtL8KPTkOiyCHMB9r7TOLkhxIpGiRJnafgiU
r9O1LUreFfts+GZl2os5DLbEoqDSlqypeTDXw+wE2RC0ZOh5jugEF+lnz99Fv/gBMLJWe+DeeKhn
RUyJn7LUd+q8XqRhMRR2ZWuv/OlgD8YIrf6J2VB0rftO2CXoj0t8PfCPnG7KG7xV4bArWlnFjsb7
tHcNRGaC9Y/Dmx1oyuZkDKUYIIKpNK5TSUFzgP/RgM8/vS89YVnUOiRODjppDt8uT7GbD8onQBP2
AE9/m6DEYPP8HFbvHOAc4RUq/Xqp5L4kmYTVDJLRhP/OFBjBt9gmpfQyJvWM1hpl8TxVJ9w4iQvY
gTVoHPZEsvjNq3dv15jiSxZO2LtYrkfU6Rfc6tvugEx44aUwK/57bSuJY7/BXlA7sqKzbhs0ttZZ
hySyqICobOSkeip6HX+YhklcMsxUcmJWH5C1lrSMCwsbP5uCfZ+OfP+LOTGS/l2yeWWoBLt+/i7i
jsFztL7jRpzKF9Zl4lrKXP0Lh0zru+ditY3z30rhslVGl3PwIJiBv2I0kJY0x0Ui8JAbNf/u/ElB
hGp6dml6SDODtyqapTGQXTfA7Fkja+yTAz1AYjx+63BoRBSusWuYyTvNUFuEag5Rv3dB2wrXOTnE
a+oIcyF4NZIF/HgkydjdyFlcqRbF9DzZhU12lZDQrhs9fuvxfQo5nqCyMFFgSYM+czcm8N+HgQP4
XkHe80mhLixkaNFHoWhkofCVkDlP2DyVrld2mF4tCV4OCMEGF/31ZoiqklWkTRxk84xOouSVqaoW
Kc8QLflpIW8C8mo0oapow46tQJWaqyKbR1Ek5p22OwzKva6xkdls3p7d06VKO3azwlU08DZYqmg8
3qPB1Mp9DPxYdh7xduMOXBuQrFm1Mohz4IxiH7c8m+GI/3eMofnuRxE8PJOzCEw0eFPY5ijfpwTj
0s6T35/oWIESn5XNhlTGhLVdqhU610JqVxJ/gBjIVvSoVxNtrJ9WDSsxjtq8j23QHq7eleIXDQS3
Y/ZbSejPElRYP44uwqUhy0WU27Qq9BsVNWsQoEM6pMeOX8j/V0kBL3HaIzJusRsRF4yrDIz3os9M
CCMNjUdFBbS4CqlOMOdzW3ESpNim/6EVr/N7dciUnuqFbfTuhHKQC9oz/tsihc2HGdGi+KaHlsrS
1ZtT4NxSOTnXlHajTIv88qqwdATgLc4ao9uIaY6573kfxPyLcoMCS+iq/5xX28Y5lzO6EEwCqCez
j47xfcdaWl0UTGoVaEopJNe0a1/7zglvWEUvRl0XRNZUYCMo+UgwRX8AY4N/uJ/jbWlKWLSJG94R
hOaUxy4pW4dRjxKLhj+Xl4NRtMagNlnFnD9EQBDS9p7DdUvX8Q9Yor2VnOVJShp1Y1QjdTnk0CU/
A79TlguRiBLA01XctDDY8KN6wUqeoZl7Hb2aGmJEzvohP3ZmRwU0XSTppBs5JQqe+NswB5+/Wblf
iEHN/zUhbQ1FXDt98SiZ3NNKGyAJkSPqCPkc8A3QjGsnBKmANEz7OONIq/j30H+3L3bN0j6zggUU
V/O/gB1KTdFBekg4M+RTgJR2YbuMTJQXMMIpWXH/oTxRMGJmNwlL16jpPO6jT6sXjvnj9lxsyvTT
TebB3MHOpp8NhRek6cGRmXu/+kBBzRIK1Wn06KwXJodsT+KSE97d8RVqfVqy0ZJ5DmqBL9TyF5db
r/aKcsk3B0Oqqw7KR0FTQVSl2GjfNo4IL+pJZ/QygbCin3aTvI8s73Zq14q99A7b+yiCX2/V8Tfy
ctQc21VeYxM7qwi64XfvkFzz32vzDbNoMctfFqWeTil45iVfpDYEeKMACtsubhH9vIy7JzwN/MDB
6JhRGx5xsLaVKdHjGry6VecMStRqWsTvBtGee8s1dIqdgfX8vWGqUtFWxyOsM21pJZyq2A0uVA+B
FFz3c4Ft5mcdly51zDn4FQb7BmQ1XCvp71hCH+Nyem+LcECjNrqaF0PYXZvR9qS9mK4+lk79NdMb
2Kwl+kHKXwNdgPTos1LeU7Vl34XZkdkEtVAX8WTaMPzbmVNvAf8lNTlUGOgppqpWL9Ql1u3pHODp
XHXtm0IzVmXQ9kfwqMnRipgMrox5OrUv+VnReWoIi7ZvlXZV9S8JPJfQJMXR93orPqCPZP8SUxKZ
OmN2dDVHl82/byeo0ZayUv3EPiQ3qre9X6nR4Op0kvORNmxVLECNURhcR9PnUOTfrKepbNNlukJ3
1T9SXqVmSnPgFWoNcgue5ttpGrELl0+THbaAxIjdxTtUkgffsBD8jJNH7d+4/0LvJ0tuYHZSFpFy
TN51sMQzhd/LH4Nw1z6dS4aVWbffHj74BOnM4gV0+54yvgn0xzeWwcK6gszGum3wzGxtJbEWuji8
pUJvj531C8RdLLGzkM3+P3JK8nP3KV33m5LxPRbAxrHRYjPHNIncLnUmDhZrN5+PoPqBxbk9hXq3
zU3CedPgL7nPVDX5ERRGlG7RP3ZRFdvszmF/wSsKVPWgmIPdKfKmN3HPzE+0dT+PeirFAO0gbysY
dzyDt3cZGVXrsKLAayqGqWy6B/kuOpb1z2ii6TKrdbVQA2KSG7szjcp7fFZqiKWG9nRSIBVUUext
OyIvxVIRQi03YGF6BgdmlLAXHL9OfvDAfb787ZEb5a6kSoEHRmSoZ092BKbqVssuEIiVTs6Se+UG
pCGeJpy0lRpksMikMs9b3yIw6HI19woRhwNe2a5tUgyNq4zYzLhybQFRkLdM7LWXasPzI7zVcwi/
80xzpL09VrKApxzINvhTEcRZtAHtt+86OOFZA1629LsMte2d3XsHVskos2mua3tYZOtYfsKTuXhv
/cBri6aT70c8C6hL1OvHWN3gCYbajNmHAPqkRNQhXDmbOqX3oTZwUPk1aAt3r6u0mBjErX17L9xr
w7fTJG9X+fMFqIuB918hB44jr7OsGLci6hBQuvt4+8SxzSQDjLQm1pIpJKOOO2SMVE0uCm1161FG
ZNKw+33t7R5NFtFamOLwFuiAm79o6aBinZkn2DnRSIQPrv6NtvciDPlHvoCVvznVZ+q5I+wIrePb
wRNRnz2qS6Dv1AyFKDsHupFGU+aGdWFSLWtlBvI1gf+AxtKzWlVpR7PheTJyg48L+rx0tTxZ5g+4
iRILOMRMT7jDiMzkm1RPMckg4GdK4F+IytnAA32JvEYPh8VUyCvyukRzK4V2uYJLC3YVTrfkCeC6
L6iQpAF70AD3IKqK2kyJY2jBJpoj2gtNSHjeTPOHtlb2rkMMyG5EOPM6jdI4Tf/MqyvE49SEDj+/
uy1Oy+XpE7vn36kZ69gSjHuo0uUZAutCb0OK8QacJVQuGIKiP6Z/fLza2x93LftwSjFlkh1K8Zsv
8fxVt2sqfGIZ5bkau87HXy4O7yx6tDumr2uy8R295qLj94OSJ5eYHE/P2599MFK1PDfjAQyVIZzm
6sB606TaAzoFRbig4U3XauchFYuPy1DEe9F5tqyfJ4rEd4XwX3gBNgE2v16IldmG6kJaMVc0sNZD
7SFZcTSK/6z272E3lcuNCg9n58ZfR584ndqi+xWz3fh9bgLQuoMzwJTzKhni7SLaGDXrV/ul21js
bNd30gEXS7qfJiWrHwT2Zfw/MpfkirPpcKFyscbq5kv28PU70/iMn3aFpFWJGldEb5RxPDaB3flB
v+Y0I/8FS2xp0ZQdISFNTpTjbNBvZwcwrCnvfQeihS6zm+xJLH5ucnP1/kiB0Bu9OhdU3HrrDyOv
X48pxHO3Ro6m1wpRuTbhZksC/f+DFNp2VE2xGL3RTL1uM6yqJuUpwJ/f8IuGAGgxtD97ff1Adcc9
gWdFufIUQCgRyEJbmSQwUaVlJmEuBCUoO7pX111aFSH4bsuKvk7f+mLl1dNqbrAwLiERChaLbpZU
r8MgyMf7Usf12tpaqwKbJKW7mYFDIAs47GRTQfGTqaiEVKUENLbnXHKEvrTKhg3WJN/YenW2u/Cm
TyRWSPxvOdQj3u/ImsSoFmMcaTJOtVrU8EPkH7MK8D2lJVKcWQVFMzanHGoAkYg7RhNt/N3uFNuw
lqMzhQdEQ757Ao4+9eau3IEVEc8CiqdzQHAC6iCr4vFWhtndVwloSTGPUMLnCGOXxsVdPYq5eTPk
lHv8v8AptEsIb/sI1Cxyj3Lb60TaajaZm9PjHsQrRLPN+SYEv7RIJKh1/pbMvKK4oDDMlCIm0JFu
brNnMmImI5UM8M4kX/CxlJ1qZ+ooQmG7RwmhyIyeEXeN3J56fFobZGlLcDWIqt5PT7howGkR9wwr
RDG0F3heg1b985+FJ6r4Ozjiw7zJGNhLVV4rmT7DWRVilBQvLGZoDZGbWGZZXkCMCOap3nEbCVCx
lRy+0sp4mUZYBTmx9uvcYe7auXAtrkNWnRtLmA7mFxmKyYcBiNQr/t9kT/8z0sOPqVmt0SJbAlm5
QN/bWT7CZQZMJgirXKsNNKqP6KaVUhOCQk7nehj3pntZmvptcYQvUhtYO0IqhDiSbcWFgk8YU+h1
7u6wbE0WLaC7f1hzq+SQsaTpFFYQ/AAlJIStJcnl4S+lWaEb5hro3+GDg3bvIOalBEpwtWxLht7s
YtHFwJdzG5K+6Cr+Z0zMrvr+1L2q36LFHSuFwNsWvvTNNFNgBzQlXDD2wQyMoPDbEnzdPZZ1WdNI
KJpVH5FsU5DJ8m4xITHcWhlcqW3HtrE4mGCx5/EuqTyS/CAekFP+9HekXPIJzIA8hHKRPUX5VHVG
WOURTWYyE9bcfietVIWg97ctd/uM/MwyiK8FL8a3oEfT2YusR0N9Cq8TKrKyrpJTVKqVgnZnV7Jz
IEpCFVAGqiCyV2TPxL6mENNf5nKqAal410Pjx7nI1BG5SgTqroh2Q7SHqBkCPU4Sj3h+6JJwo5hW
92iLqZ8LNqz//IpQ6RZSulJbcoqmljvs4HtrgnTQ1+I6Avf8z8Rho8fGRlS25l/MnDazj8z+UZaq
mRuHhcLaLnKblrDOlO6ErliHdvq/Zb6RnvqfvNYqF3ly2waS4UXo6h+Z58CMXiR0Ei9x6pn1v9u3
yIr4CLa5f8OVs7p4RpS867p4JvWv/eWBGUo9jUpJNBJAuY729mUZ7+6sfMY6XS29/C+D4VDCuKiF
NfHNtt2xjqUcIOqH6mqdiCz0AF7me2eXjG9gWmUNLnOyI4ACwwCgxWBDmZ+2jrO17SMGVwOpydfV
pJ03AqtJIOLs6B1O/E/KLAT4Cv5imjgyOVBUQcLYUPw+VEigu+f+rAb2/lC0R3E6BBW3YTBO2qWL
yLAvNVctzBfcwR3Y/2D6V4HEnoYX7ESmh78pa2K8Su2HIqbcS1Q+/LiwjFczECKwrZp893IedexS
9JhsZx7+sSnpHids0+9Wxp1BqqvEdPH+Kt+vXD5rj+mj8xpPYY8gcz45oEs8RIxsOeIjOgO+OaGm
Drj+6MI2OKpYsWvApYuJHGNh99d/TjolF4XqZPG/ErLoYQcduZDZ1+ry2kYwx7UxHAe0J2muJhl3
3GITmx/w7LNWLgIesq7ZrDvzdzKqFQpcVZgC+9OqCaU8CHTv2r4zCIvnCk9d2C+icIRc0tUqHjrs
fJUXfX56NGz5l1txo2RipwjhwJ2Fj7Gj/TLk0Rh0Wqtbjek1KUj4Hlbun/lLGhnLyT24wgtz7jQI
zWBorZXJQj5O57pmMjJoW7FFiEje7Yb6SMBp82VZaSzyX8Tv7DrZWnVufyMm/ejT0h3osOKTftom
H+GjTCp/FqsHFf5/ekW+W/MxkeEro3C8MJMEriu5BbbTFqLWadUywsg3EnQgDyCCgIETkvnyXSKO
XuLN8SNxd+QEF9bhyHHJbws7LGTMs9tmcEdgk/t8b21GphxwphJZULSXohov+j+p1GoFIa6tKGW2
qXxDluKhBV6iLI027DuaRut6ekDrWpAwEWqKJNwZjRQ7jWiDcC5HxZ637TRqVEacHfsnZ9n/JA6u
edC61F7cklQneN/nJb3VoGHLeyUuL81cqitVi5HWWNf+4rH8lwx8O2VTzRb3o8Pt1vFXKHuqQiqh
TFSmk7I1JZ2siWwfcf50/pymeNp+dXqsLNCUb/qySiHCVSJk2WA/OKcIqMaIPXkhelJf/2eXxH8T
71WLaIeA08nBRK8sU+yMdeHdIS5DBs2NYxGIUp282e5tHgSRgTatV590xBLmgmbr8jo0mV/peQj+
T1Fi2gqXg8bUF6KgaJ+9IJTYl8aBMaUq9ZulIiJHO4GgrfkUK12o4TD3D+W3WOt4B0yCDGBXvV4k
/5JbiGdtDkwHYq4UpecjpBehaIMQEiNmBO1CnW8kUdbnST104bpGCjvb1Wo/5DGrdkGLDa6hx9xy
n+9EBWM5EMv6YuZGZHQjKJCX3LTEDTgHPs5zNA7CnwI3FvGerqWgAKX3tzQKPGiviuWlGdjBoW87
UmGv3eJ518EOAajk8b8eLzRO5XWCC7cEqA2rit1tLxlyrPmpj7ML364sGHPrnSQw1aN/r5ot9iaP
D9NPOB13NkMum77u9zRcnCMnU39kp+faestXUN6f7ulyBIyVX/Y7U5sVOlcCQtTn+Q7QiaWtlUuO
q19CF7Tqxw02+2pyRqpcVue4myhHUF8RHYz0zsfi9kHuJ8MsYR67F8Dd1bln9yq8j2M694PhWdsq
Oewcd/47eZE+iWQRM51fGAavlbrDwz5dqJjJgUVQq0MuZJtVb4JN7JachrnjrFER9khjI2SY/0lD
ZUtqiIqoJchHntHmJgl+PN/Yxl++QgPyVUWuLePG9sEl6pzP4EdzoWOXS/VjJ2vteJvuiXBUXBOi
piq3RD3IjJiwZmrHlG+N/y14Mm60+xiqrtBGs8lJgm52lLlVdogkvdvYjqfM4Cz42tc/et7sqe/X
RMavN1Ctn89I5ZdS5MC+Ls/wx4N680EhJ5j0Pyy2cH3YfR6tP+M9ILpvBs+GKVD+u0jmrabBfOc6
f6WmjPLqdSunro7TQj8QRQq+S28vmKbrEJDdTml8b2nw/GiTgJIeohSCwap/cAjMWn/rVu5PvldT
wC6+eQ5CADu0HcZeN7J+1b4zMEY8WJWC4QmDHgwq6Y2YkPCoZKWzgh4ENfrQOkv4FHMRoSWfJDuQ
AbvfTdrstjqOUujInAui/yrG4yz9Rppa/YJyem+w6S9i4tuJNpIHMP+r92IUlEIIeZ47pRQX/1+E
Od3gD9l3VTZ/8HnDeab06o90nXachrqnB7C4oAHMBkgMGx4ukEtxmngZeLgsYfSp6jk10J0AYGKg
lAT5KAASMqtn5Gqu+86i3CX3GGPwzm8Fs/6JaruCRejyzYJfyLWBd2wsLP7KSp6JSEygICxEsfMe
7b/J/UrxpD+DQDevBe1aq+Kf4mKIJKgmZ1t1+9A6fp6Vw7o7SWggrtgFNuWvcnTNwAKtgZJcT5jz
K9EQErj5JbvIFcB5LLJ1eiAlJnOCunSJse9Xj6so5eagUKv13YWl+XOwXfYgMZ4qnVx3KzlecE63
RaVNEmIPbVn3S6G5cN8v1jU4jP6upxC97Q5ITAY0nCR2Okx6QKJetcTAtyPxAPVRUj9Go+R8+eMT
vu4mEJtkHEY18h361a/91/Qo2kn8CXNDZlJNn3tMzLFsBJ2UM3axhdVaot18zen0rHA/HZzzvv1b
iT0EYwv4ExSEU0Tlr7V+vYvKI9Yihs98nEgi2PEJDw9NRNvejx1eM6LV+Ntx0AskyMIaJaPdV6zO
SIWLj36hNz5a7+WySdn/AExPmgDpfMXnMNqEVK14OGZd0oCFgmTe1HDyfhDSbjmNH5wmQBfSMfoy
jiuCwzE6EaVLfrzUnHazZGFGSTcGCPuOBLFJXujx4As6QHU94Y7DLaDxhTcNQfPA9RDNXIoi+/hw
phrYSqxl1OS9CJh+RpqG7l2Rj+OYlaMPll3V9UpvI7Rfeu4ool8ZElLcHHKaXL/LMty+soV0yImw
SfkAy2XX9EgrcoHX7A22dOJu2tXWkoQ8VMDzGQnSsBd3H5iy5AF38QJri4g8EQN0OnHESJPOQvLs
83phcqtv4IX81uXJa08T0YMn9qZ4lH9jD8Ux/TOhPJ5tG3cXMstQ6tepXYjj93ISuAVjGhN6doLb
vrJ9NgR+rnDDPI5g8ER3UgLkbOADPD3Ml5yavko5eUNolsNg882SxnaEzCQC+nM8kTjYstgUwXy7
jaWG0915rglkjQ2tpLmKhR3a+7HrEiinQDfccTDUqJ5IHmjL+bw/yknEzBnV46M+8DuZbBUJ7IEb
Tw+64Hj+/c6w+0VTaltOaO1t1x5OYVzbqKPraeSOZdq4GN9QIK1q0pp0jc1bEBT0zx8cFw6VNlDd
ObzPmVzBtZ7huxPC4N+GymU+C6pSfRNWH66EqbozIlM2qN8xVMATE/MKCBmLmYb9q5MwC8OZyM6c
jiQy9rMJKt8lyxNok6dGvj+xTgu7baCzZ9NT+thVh1LN566c7wSKDYp7lYv3Qu+K012sjHkq7WNQ
da32GFqq0bkrIPj2aFKot7z6SCFezrJTvg+JvU8StcZDymxE4vz51O2X0603OYD6R2BowwcZp5qS
l8mckDy+U+ZoOyz4mpWhfBw+GLdRYqVnCRKRmjl7nr7ci1NTp3ify2e3IUqnpj2eDEx8y+WhplVW
AHZzRolGa3SNE1zfxf3ENUrZtfiCkrRzgB20PoHtIdjeK7LAlH0wjisv5T0Tsh8786Hl5E1Q+lAV
cPTNyCxTDzk18ztLNoLDNKg61wE/KcIcC9AqmEA2AuNIprNcL5LxJ/llWr09ppPWOoF8O36ltJ8E
8Nct02VgyRmhzd08QfhqlPcFVyoXoi1g/40ouejgD/ucjQblac+I4PbrBUDGIGoAmmfjnGcZq+NG
HztNP5XjlZ909zGFzmioqgHHKgLGRt2bkQbUCwq2W6ctSyH5V4pbc2MXrm7XWhhLTz0960dbD5kK
q4vNQlW5qkADYm+4570umn80E8BxEwhy3/vBg0RtUrQBm+YCDRuzOVUFE3tD9B6trl6aV2OL+RSy
QYoFT4K3tu1LMTU4XnNBTAMgDOPunO5kk+d/GX1URvu9fnisbW46Q2vkEXGjZD7odUfjLcobAOKu
LP3ZsyZGR+1xdp2Uepy/C9xe72Y/e74sBQRAZMI8OnlAT5UZ0rfluQlRJKoZpLlKu6Afq5XwVSrc
jkIUleaqQ53FTjaMRALbC6He1zmJhLp3ZfEEeeA2QYKA1GiLqLUuYQ6iJBdqyz6PlIlOD17BDiSf
HucMqbWqt+SpoTvrAHuyLDcDbitpIh7MknDc7RHLwXYPKKvLEjOhTvvG8kABza4qGjvMSIZX6npA
eqV/bN4iBfBTKWBYV0AGxLLn1NCh1nnv1IebdxMdBPOk1ndp7UDYWmjB5GiM9LzIi/vXicsBwrEJ
fVPWmdCL80inIA9h/fwm3WhAikP4HLUrAB1jfkM9ydlUS0QB/nWXiGOX9YPSj5AH4e054cjuTANi
XaU1NT3qnoKWPC5GV8kpjAKgqklkzdQQNRGxDcnPFtsBiqfFTnTFD6CVSgWHlsxQj9PYd40XXneJ
YCnbpN69UYyzmKwqnrL3cUinyWL4WMO5DS10iQKnCAY3xnOMbg3gRhaSz8YIk0qLXAlRVse4LZqa
RkI7sfHBoQ0Gbk4kCAo1HQocplE6xkobqXLcIVNHAeNZEoCujSoiWQIQI0SIT+CPwvi2qK+YC3uO
6lzOlJk0ZAqjJG8p6Rvr6nblY6tuBvx6QkZIuS2Icgoi2wnzsSVZ8zBv5ah41Fmfnw6Zuik6OqX+
gtCbAz6cfUFlmhhnts0N6MeXHw6ZpP4U7Ix3XzxTKl5GEvRx8gQxLl+W0yJizio3ojkCTINd3PRt
NVMAyYAfmJL8chGcxJXKqFS4/VNJ5B51bRB1IZ9cgjzaFvIHaKzULJW/k/5X6vReXjLvPq8XKhfH
TxMV8W21EIt9eGVhLqqIKVyAXuMyJuVVvb+ZAp5EM0ukHdYPuWF1kJruGbTOuNMqYLGVS8A5s3CW
orYKfwioJtGuAcJJ2F2D9S32nrpA3ptFvLALTvOVUCiicERY5o8fMHjyY5cAFomxtvTRNPh0QG5M
6xrux8UyEr4wZFGFlYt9cSvi0EsHsu7gRbTjTU3EymZ12EtKOcyX/SBnT0/dO0vxnSKFAzu6qWUN
MmHZNvdIZp3eVogKGG0TLVA34LraeS8iZsBWh8RLpvtFKKiTU3z6duH6GyZW2G8RC9PATmbNBXUV
d2ITWJs6jU2PKX7AEOUusYmnBqxmM1+T627oabdboJ7pzU2wVOhk1eh63XWzb7xPI32ekA0MvYpF
HriLh+GDiTpnb6R6VsiQmy5HOvJJsSKkGo/Wl7M3qrXOmAfXrTz1fqPZwtVVHSt9vWPxYGcxmh6f
t/l62ZP1mSMzxpj0GvYvTBD96plZ6QzP5KeEBE/RAZ4FFOTgWJNzl8IOercNTUcaTLzEhEVWWbKZ
/mdnvM6+O54pTjIPabrq1UxgWB9l6KPzr06W7lheL8EDANWLkam7Ij2nBEgMUjT4EGgHDY2Muvvf
BNmwDkPCz8vvjKUgIr0ob7cI1D8N+Ze0BA3a7MQvOSOGs7EOVV5lHqU6KXjwe2RSPO5p89UccYVe
2t0aJG9uiUK1hWZqi1a3dVNsuUKp1Trc6fvVwnqfSdKuKKBM+ePVwm36jeyyUsw37EZfexyOJQC4
C+YW+F+GqoHJHbzWXK/fRACWZVQfMKW4XMHGQsHhz/t0Yr6YNy//HnZNYndxpq6uDlBttletElxK
m7Ubg5bXrWk1n3KxhPhQrXn7c1+ifNVbfKP8V4clHeJiQUiWbFchq7WHtJ9bqc/qLRmJjaA8A6Wn
Raf2xM/y7xE/GwN2MmfKgu0fr6TQtVunHKUfaPWyYQlDM8lCR6WqFB55uc8yApqEsPvstP8QW6Aq
KopdcPyxFDZVuPP0xG1DTse6DgaZsvRSEglOQv9/fFOjpAhcnm9ct7BCtXo6D/SMxAVLfWsEeUno
CvgPNs64X2fLkMqiBVNav6eEFBf+qEHYmXMK8EZXuiFDetVisiHS9nJG7anV8RAhM794PwtjX/zT
bccRHzGiJhzYFJFzMRmfmj3buvlLsDIHK9NOx+Gn56GsDhgMbTCBoG0jyPZn6++1yBH6q9bjOw+q
hu6kZx1SmYzRChM+FKS8+3TcxLwN2SUcNJmbv6AzlpDMCfUEBs40ds7tCmtdWUd9y/+wGRoioXCR
cPLkWr+/dcfa0AC0cCfRAdOlN5UX8oXITBdlAOvTNlaE7zB/Cj6ukJLEmhXb5AdFmn8nHkdPAZhY
UdzGoVJCSMLtv+EsM/OmGld1PLl/jUgOgqInsdKi4pjVuIJkMAStJ7b9yM6g36zNEVRvLwMophTa
KYZRObtkwd4ZWVltBvIjS46q1bwkTWU5eTtrv1+NpPWu8GN2m7ycefqqnOx5EdDJdbqgpVgnTZpu
37UBRnu3skPcVTPGVUMthyXzpp8VA7lmTBNrlpvNGMXdOE/NudC+ZG/idTJnB6iY8Fok4YTCjH1s
V5WzQuj6d59UYM3X6YnIloD0Q5LhEL6Qy9RNkPFXC5OcxXAQJMQTP9VRFoo7dMx/aByCINFIcY1N
I4LRaxXSDOSib4EDmxd12S0R8xiA7hj4E48J5nEoN+/F5+h8TAgFFwVKxQS8S1BeLAxHR+MvDB1D
KdwVXDmoFGAaljI6DwZtB4TiXkOWbgoJF/Nl0KYWjOIUJ4tHpzElxAt2249XuoMn7nLTBO5e8bJ6
8HJ+LZ4S7YZZbOdKaM7DFfSEtIjInaYQW6z7XP8OpM8hM3eLtqq2cWAQTC/PXh59Xi0Ic71fePiH
iVTK6eCUvCikk71EV6mKDBd21Ici+IVXti2ZX/b8Oo+OMrlmQbLhF6b4sfg4WGl5Z1LOKB9G5EYp
yWxzaS/nusw3mXdHJ/NpFsKjTKUeiAgludhSWs/3kMdpW3dewQZD8ykoVORuAuh8gE9T0itmaB7i
RHaja3yLMpSV+v+2M5qYu/CCQauSd6bOWEyiQe374s7F3M37HGRUGrVEVwbGZIpEyp7SNe7z24Ad
wTUk3KcLjPm3n/XdHrL2Y9E+s9Id4VBPitrYJFuwUS6dRImYO4/e1Uy63oU1dvjxXl8tmdaxm/GD
ZctUJupp6wSOWR3dDWxBBGN+1tJ63fDk/J33rUQLrcCQLcAG/GAVwAfPO5hgcnxNtJ7snz/V1JVI
3Mh8EnNx5f5ISpTgDWphX9U0Zk0GZYKK0d6vFWkW8x0qjUXc6eIqlM5BlvaSSMDlY+6BehSbiQ0e
PjGsVAcWj2X4AyGGc3XdPbgVgc8oN0507uh8vJSOR3LATKOmxrmyhkSJuJ3szHFfIcFbVnlEwngc
8auoIcdKLEvOjvYyE7ZsKO5FIpbVUTLZyg7pJuQntHv82TIkoJtovBKKwVSskBqtqgi8DsnT0aEM
qsGTQhWiEuUZH8Y+dS5nZLJDRHRwzZKSw9jlkZBa84Rn6hIdtWCgD/oPCnbKO+jXa1ERqL2u8bnQ
kkhpuGP2H/cQBzwioSJInCjw7oPzKVbfAcHdm2t9msTQRyln0UUxy/OnPxO71uD+8+gVTD2yWeWL
UJLnxh796ibK5DiXTHFg8qwnSHoRhFUM9zRtX+vvYBsSjqyr0YRfGPPZNeyQDDgItwua5qac4Tsc
JIcvZaVozoVn+I9sqaFTNorcdoUahbkfd3iLnGvDvShAsgwlB0Cc9zR1CKOKw0Hv554V3nB4BQuA
dBaW1azOAOM7Gxs2dnMRmf+oO2wzf4L9O/R9DGW0cSglm7uCl68VFj1U978CHdPAffhFYJVoML05
NlI2wtYevsK1U86FVSnult7TsZnG3nHJ0HT1BtZD1ZtLPEvyR+oHuDUpq3NHuxkpf5a7vfPRk435
wYvsB6nxOY6pQEURHciwXtMe341furoQaYMIJBhP1k4QN1Fdn5xGRUhhJ4LRnPBhhZmYd6eYvw99
120mcXlv7een1q0JNPJmzspQ/nBMqaU4qBWRmjtCLZfiembBjhj+rhxgWjP9urJ8CKaXPQLPxSxV
lbXAsk5RFSPNHrqzEM6nfuX+EOjf8F1xMeXsl52cOafPLEOaYKWwKRq5awc09wlOiRk7p4GBcvpe
UXcK2zt0I+l4dgQ877U9Q0+qWU6Ma46M3YqwxgTAcPtQ316gr/RclYwkmA9pFD1+13GJGKAfYXln
34cvzqUhIWBoFb3bjnYy8hdrLCsuisR4L+6fULOEOGQEQXuecuJkK9LiZq+yufxPNpqhVlLFhcc7
LpUmM3kBvHX318sXb64k84BPBsHgK5GqZ9t/ANjXOXwFY57BpW80QtOyiCgofQAvIlnLxszDyHOM
wQZtf3+jD2joSU44CwNunqMSL981wLbYFk7qTU84ntFpH+I8PFRu7vNZdyrj+QFQDJMSIOTevVNM
W8Og+KGsHVgXQpskDC1qnvvDkRCZUXfViqL1A5Qy2OnmiH/c8oiqc9EnbBVXF6hqPNBq1OtjvIEZ
cgeEp8kM1KD0ggWaohLFHIYTI11tMlc3OvXO7c94zIE75GYaglJ7s0JU07G0d+Oodhq8ny4Khgv+
08zUiGusw8eaX0WN5rZzO00Jv2yIrs6gWopxoI4abtARXTAzR/95bTKyBOU9gJU8XMmRs+WVhr88
n59cuB5mSmwnUaTfU8EhThO8LFuNaxu9hKCgvqhu0e7D05kpb8jHV4KXVUMUcPnqGB0GxKOCoofw
ThZQK/USHy3uT+Qk+HOGAsHcPaU3Z9ZEYs1z4DC6J8TSuknyn6saKrbTrr55ZdW5frYyunyjdDtp
mQekwLAIk1njlCDZDwyVucbSVpcIuMU0wS4uyOWQ0B5TVRMIjbqWPQ7Jk0MUbhHdyvhLHNKUHqyW
YiZSON3k8i16SlGB6lWQmyju99ISBAPQ09WdYzZ2gLDX7MspOzq09p2Pp23S+WW3DQG8LSDuk3Pq
jSeg2zpmOcY34ss6KPZsXvB0xmHeWIPeD3aoADeDNsGyC3EGvm4gZ9H5jK5wyeKso0t8l7SdNn8s
rEHtWzUfVJoi5XWZ2lzOO3IJHI4CrSUxtCSmwsWLF1aThWZb6eRXkRSttzqIMjhvZVy23jQWzzmF
y15S0UWB/mYZyT57iVjlFxFHkM6xzimDb+YnmrSjSZv7w19/lWW7+0H8kAHiP+NF2o4BoZHVNDeM
02pg03YV887eDiF7VziMVBee+dLgWSG9VAvBXW+19k8aZQlBusBL93Zv7fFIqLc+af/h5HydJJzZ
928FxwfJecDwgaicQsDKviz00NqxuKjauH9xIckzjNOE098UzhrHQUmSR9cy1ZgYdE9Sdhij5T9V
t+RGmQj/K2yy5ft5T4ykv6Ya50i58gKxm0MvPsZX5h8U1w6VEwIaP8+ni3eCnA9MFOVtnITByJQD
vuZyxL7ew29IIH2WV5L02yzfVan9Z+TpwBc582mB+pwDj6LmyuhZqvqYFwiByPx5wFvOXqPgztcd
iNM2rKY8oB3sSL9G17Of0I9j7ybLiqm86pGob4gxgjR+Mt+E4hLV6Fc8jU43ZhfkXtUbQ3YANnRd
wfk1qgw9+g+4bDpCf61FcZgJs/j5WKy3Arrg/GHWj+gDjtonkwUkHzvV5QbuMlXtNbdQaPllb2k1
cC9iWfBbsUHiHbLUOXk4TT7bYmfp/7ShMn0xuLSXDWhT4n2SB1P01yM4aPBf16x5RltMVB41rdg1
k3BcLDPFEHCwdZcZLBOGaAQU3oSHRv8hVtiFOztxQG4+NB8uQ20m0qy6JSQdQIm9id6kaC+P2cDf
1s2XipYgH1Jo6Z80CMCAkPp114jz8EzVfcY4O0jvQvEmPyEu83DzzSHcnmK0q6A0ReLl2F2Gs7AE
dDet8JfvoOjC1c3g9U/jCSRpADkjiCPqZ4X021UvnXG0278YfyhVTfD05uKZpU9sflJTW8xShVdt
Pq+KbI/DT2bpzKm/SslYnLuBFXZVrIoSpye2opdvP24KZQtk7avnB/ttk+m+xPW2G8zZjBQpWyy5
SPpZnk2uiUEjVba33BdaNJZ8Cz7xHpPiLHzmEiH8bkOqFDnWtWtDWNAMmWJqu1fi0afFD5h9AXkZ
mTZNLgtu1JcIWEOApCcJkaXCCBfQv20IkRkFF+G2OQVf81E2D3V/jJNgMZiCseJi6nw2QZ6/r/2Q
5XuMlxL2LFVnXtrmsGy792DpmrRroJLmG4yPD70Hp2JnpC0CzoUJiwI9DEGdbkl3boaPX1GAnxSb
f97zYQ4av9VMM2jTsI5Og7a0fMUiuprjXf9cwOWQ5UzcRzbOl0a3ehQYbvja29jSnxYEu/8I+Pas
Xx04sf8dEtzqe4RuoqwDfDNyJ6ytwqCFcN3apyyZ31AaG70SABbRuohmBNEK7NBg1UcAfHJDxZhD
h/VIW0LaLJQYbCnuRjA2jPW/zZZ01XCFWVufjpJDr67ph1DZGZQq/zw8VOBXnXGMe5xE1sm1NNqA
r8sJEg385fGW/X4SNYoAA84khwikcqip+n/Ve0tbaHPjMFFlF7VEZwZZbxdzaxGf/0290CywcXI1
e+xPtJO9Sk5ZDGy+uaFT4a8veesuNc3KRiGQ4YOtvynWhy/zNNn1oBht0xA/RMjTtP4TZdE1zpxG
NOrG5w7HIDmsNkxouFVaNA5jlO+XBRT81ds6hXFLnbFkr+WU28oAoDoIxXf0dlkIYXSTO+qfeyZD
78FKc+3iZbtEcb0vOwHgS5sV00K9kpNmRRC4Ro2UTknAcJ4xhNsiNIclR/uN+TZi2t7rucqHdFKU
UnV5kgvtJ2ztkozn4cVAooxOuxR+cDo5ekVpi8NTfkUxmWqjpUap92//hUt0MN6BHyUDvGuzBfQL
QgLMP0rE4rB0uWyy6OIEyTbriZ67B9SkJnyjDuebPJ5hEHLX1M4sJWFKOPj3fzeJu8d5twV7Cz2u
ankzRvYhQeH/CjoLIeKmiPUR8k4nHcZHAk3yK2x82QcTFqmQka1L0A3t2sD6Txg9dH7ZHAIFp6WV
CkrKUhZqmCJdwDi8SaOtckLli2SyH0eXTiga1o+HPVuCfqBNs8fnMJI2K571qH6Y4UZoidpqS0sh
BVzz2KQgW3DSqXONyygGKUDf+P/0rZTWBk/mvfjNuJLWsPRsQ10nR+PeCbTkrDZwBLQguW89e+wb
zeI8hGq/WT2Z3wRVUlkZaADnP02kumBmQxYElTOwQQNryE1h0+2+DXCZlkjNparsIzD7Le1YCBZE
TDZN0NErfTvT6YYc1huINwfLTjlpKm7RFZ/F16PhAKUsoqxLe9pYVCEga3vvy9HMEBarxuMj8JH7
XZcKnbVx4AEt1JieBMLkvs76ittTts3yhajCVhKzaZqlW/bG8qEvPKcAFqy72JmV9hDMcdNoMKu2
1xjizLhPRLFt8ZmCOrEtr0wsTn6hvSfKdT1rHL1L6CMdMGoqp1isPcOqItoFb3QhhVSHwotYfHQd
OTkgF8v1yAkJ90c7i3OXeURSWDpgKM50gmwcfiB5pshjG/wIgtsJsPuFRr9k6grWgN9HZvBRnzWF
thsulRkOL2SiwCwjUOGuDlS6ke9TCq6lGNS0ldWNKHS8/Riiti+qhIGFnWRHlcD0hpxRgESgBqTr
+mcYTYUpF171g4m9tfvBNCjKcLE6gNLc/F9DE5wlLPqQQyKP6rDPCiW1xwPaSfHvbjVJOeA9q/Tl
WvP1X1TE5wZ72EA1FAtO86d6uZo8bfrCspN3cNJBAMq5zPmSpQPrPlsgvBokOWWwln2QwvNUyP51
nbjeXysuOMGSV9pIBCQDKV5ONCO6aWs36GhiPfA7lL3RfUVe/VG9E7y250Mcmc8Kcg7cRI8EvpqU
sTY1dF5Q8DLvUo+EBgDBBJuZxYIHrj9NfzSh8IRCnndT3wtA/mekP/Gp0tlzveSPmeYUy/vZQ541
lbif/U1oyaJCbUeDCRm2UlMz70OpuiJVLxKGT85rtRJq7GWLBEaDB5GR7I0kS61d+dkjfW1PNfUx
aPNkPeFpk675aRgzO3Ld3xabmas1LTWbKKZZQT97NKXwb8dDWze1ceqsdlNgJCryTUCP4XPDf2iu
8SSPnxfcZxsyQzF4IXx0Km7KBWnfdWuih79qJPY5Wpwzw+gPw5fQr8pARapBBP74oNCvOcjprJoy
mCg39SwbXyx8hepcnKt/T9LYFK+20AVnk4xaRlRaTEWcq7ECIM7GQLzH3ciPElWsPXQVAeJYJdlq
zbBrtXwHyDiCefTMKL5SbYkVsg4RjeYU0U1BFALObff4mZCuonBmT1Nd5usDhU12WUufFiazLl/K
GOCCV2K/19cDVLjTPDs5BxLXl64vojpQxILBas/Ll1ajmHsYfEkH6DyCaIue144H+PwQWDWbbGWx
cncyi6sb5efLx4vWXY+OornUE+lnfM3gR9Yt5lewkbMO3D0uajds/RTvxdHPB4tYl4H6YIKy+6nh
9pMqu79Lvb/YQvKVcNUoftUA/lmrH4+1yi0J0ZHHH/Haa7GdT4ts7w08ncII/j0fPIvlWIGpQk1L
1NooJZgP/Uc0gZuinPDAxnN8sH++aq29q0HPsAxHp7TDYct0f2Msdiy1myycVeAwglXhvjBJuBrP
vaEyrbAups+6g5CgooC6fAaypKRlSZTKaUQqc4+OCKPPenrH0uVWE/u7lINJpzZYlCWJFQYffK74
GVonYUltT7+u0XAhY+7WyzptBQVQA5ZUnqqKydikm362+O1SYUA+jKRdzF5UAkeWLlH3+pGnSbj6
1XvdPm9h5ZfJPirYJOexKp5OVKJCtpQVsqLzdqoz0R4i40bISP9WsCMOYxXUYoHYGSE/C8nHuVjl
H3GwfXYz6UFekR6o3cWrA92tvOulNujHD7XBajmrCVdzgoCl/3IClgOKeVkMLUqktargf0vjo+xK
1kKmdiXsWbVNKVzjq+KQqdlRvIoRLoPCx4QsmJZl6P8cj7oRcmnNWH7zwxk2jB6BWfwLR/V/884p
sUKLP+pNMXK8zmoJ2KP1C41/dUMjds2hgk3izGfSfBt36TukqZkckftcADamcM2KvUgbWDCj+Km8
iV6Mh6MajSCkt71z8MI5qLH8tdELcpq/urk6Ml86KGg82cLnwiqQI5PzRZ80Tv9ghbpC1kZLZk5B
q8xrwNbR+gd/RPSqTiofs4v1jtohjOkrYGibABrn2vaqtBSocWAwOWytYQwhqfZ52FvWPpr23gba
OVCpJKszGaU/m7BI9IkcBSjEGPf11XS2dPhjLrU6K5vAraJa3vmtRoHX/T3Qz431g6LAvB8VtQEi
FnXkSop6pl/EoGxa5fqivVl9UK0KJ4CgafjwFixIWmCM6nrGcLL/RFBHNGO3np4KmMWoqsLzNKU1
HxxsfjJx6ZUfdng6+lhXLqHjt3k0j5u+0izP2E5XpS1w9oThUKysUPcYqhVxu/b8cU7AVQ0GXKyU
ATRU8FrSvoLMRm8f+s1Mf3xjMytMMArbBozt6KNNFTHrOsXj9eCe7utYvjj6tybBmym6g49rcCC9
ShQ4+ho2p4wSogQelnRIBGGhkaQWRxHf5TaQhziD59hjeL3t9bFPTJJl7pbj3FXP8FPLraAbcZRy
CrO7n9Q5bwcoj7og9Svq/KgUXy5GJZ0nL1lBBwxm6hqXfzOJqjiNMfwE5bcwwyBdADjwwmgepGZC
uY6tYoiTFQyhOBnJFXyFb7CDxl8WPihjzHkAgm6Y33ADEV3PYA3gEK8wzvrko8x+29s15242IkHd
JEz7WoxE90B9d5BaTm9ZXS8eE/PZZj3i3gD2QLuKmYI6DXHT/YRgMHL/Xxr8uwLl56h2VLcAdS/a
WGS34cDwKqNf3SIhbGxPanZU4X3A4JQRUTwpfksRRMsmgPfguG72StlgvrDerPfHngi/RtZn7Uwo
IXp7uvcN/inKCZRlvqSbFxdHQW04Adl/KFjsebkVri3zLWTEYY7RVoot0WJG/XHPTgzmQWUlchho
sXa1HH9TMR0tMapa5AC5jbXYp9M2LKdkPHlnCuy5tseSrG/PrXVvkj/HmIhO+ADPqDlCtfhoyd0i
maZhJ2dRCOmB4B+G0lILZJI+Ar+T9nLqw3gkhCoo3RX+wcw3pi5XQDF3G52esnCgpwvjlVsqJCWB
yuJ8emh9DLePQfUNh630889zezMsAIHpSB8ECdwfCuN9ET4/bE/mIS7uVupAMKqdAVreOYzKjxGY
RgGj8kt6+X4hL/DVlyFO13GAXbrq2oQ6f7lbwRXvFdff93o8yKICXv0l9Tw0qvi113Q6yA2HbIj7
MZa+FsHwyXTfpnSrmF37LtBUvuux72aMUZBF29Fx9dAKn1liDt+0gclaQokRJ5xAsayKqHEmgM8k
1chkVL4Qbi9RL4izzxPV5q7QuAcG+4yxMBn3A2ABS2M/HvOb3wDP1t3V6LpoR2WB0b/lRZUdw4ql
iIhbpUC06sMdEJnv92DFQfeiES9qXLfUN8ILnFSv5rFOwmIqpCwRq7a/dY0x+9FODL6aBhgoWqNb
SDafzbuswkR/gie+QTybvd48tZbyRPGji5XQw/gujt5eHFWEFdXEmFgRoSDhdEdAUanWpgwZ7mtS
A3NRvV8xri8qDLefI8qpZ8NHDL790xDR+vDOFGe+VTZqyWYE8P760skjT6bXsajEWbM0Ihif1vun
RiliDS2g3kGb/ZJkrielhS68OH75bAEq3TkXEqQmYCDc4vydQ7crcnzGDu06nFeEt5pvu1YaTgL4
v7HQbLqrhxXTYhnWPoq/TudSmM8G3EXIBzEKHrds4Fpo35D1psvNEV6NB+09NFNUGHkiweOk9Ow6
TZ8USsvCGHSI1WqDpDiw7xPZquOHdIOKUzKjfUH+96PinFqfDSj+LosYKW+MqYSAkiKodIknXG0W
G0AZ7NMlb5KRmG2gcwwp0+7N4lTvRDqQMLKs8VDvkMEHPkjVJL08oQNKJ0uaGq9H4zsKQ/PiEGsQ
AWVfMIyv60dCyJbjkKA0cmaeOONm6s89SSJw9cd1Xcx9JsE+J6k+Sw3BFik5+pXqibOXeI+lm8m0
57BVnaEBxDyaq4M24/OLlNhVW835YcnJ6f3RmsWZd7JVVF7TAWrslSDMRhrYsE78CRNvTAQOKaBM
2ksa+USF1cfzWoOu0sPM41DjzudlGLBGnN3yvk627unl8Qj+cnRx7faZjBE6TrQu89VMvXc7/udi
ZTWa6j6uzARxQcb8SR6+i3uZK/aZwJX3ZAdbc4sDpyHclzG3jIIjPJHV5ZzDyKxozsAGhRh9V6Tk
FTs4hsv9+YyjZZDRe8jNPk44kT083BvcD4DSFmmehRjytxJH69bfqCAVWCtv5OM7zm2UqVmUKoo0
O8TBmlic8XaARODEfHGx3YZrKKd+tgwR8Ip3/QsgEViyiZqLaV/m9zRntuhPzSs48gU/laDvgD4P
b9vJDt3ARslmMXfYzZO7lk0EC62YLv3rKnXVnPC8CfwU+9JjBOiNa4Xg4oGdnUZNFA8oz1pkPOnZ
ay0NzBFFebsilWcTH6hT5i5SBEbrvDPJsRZ4duncoCV7NCsT2UYFGwMI53Ye+KCE8C/3H2aknDib
cnoeg5agqK2C8a4/3APtFeKHSUNlVlPvjs9pQhf5F41V9AXmadACA/1pHPLDsUDoD51NjViTVqet
1w4U9PdXmxLA/IR3a2oz4f1/TChjwHwU43YoApxqN3/wU1knPqioAIzW0SjUNgnFN05W3JlzNPdf
DZwkxGTFO8G9Uzofw021c0LQgqQmXoHjnfTH3Duloxu+qKQECT2IcOp+4y1XbWZeUshKJpv4NkdR
u70syzMmKBtLm/Bj3TKihFKeviw63lTvshRN/L81iLM5on5XP33is9UQdOWKrfNnHWB8gK98MFY3
reONPmbWAIF7we0zqZcWMY6basaGURNTIMjK5UDAvmZG7EbHHO0BBKrOvDXcpxWNu8P5RfuH+vas
7QF6Y4wJS3zKma5G6P8qoQdz4b0j++bgQQzj7G8Sjqk2dCvn5gKN9i7Xl5HWR6LJoU/WwTEfWdjN
Uz6G2lh5Wjpe+OIB53ZK0WApEmhIe1HSh/CmeSzl8mNbvZtuUl8G+4uwX0JTibU0PuNuyUwnasBf
94AyAI0R6qyqNK2RR3OYTd0KqleQSs9f9T2gC+vXPXratkBKM7cXNeth2i/elml1NWgs7OImKOO3
JNBY6YHq9sZ/FHlQKCXNfbXxQYtR1sAD0UechrlM/2fOhijcOwNX5DwmnTSh75z8bdj5W9/WKObn
soin0T+BLLoph8D+MEB1ve2WMu6ey8BUKx5oarjBItNGpvHe2WWvXoSq7i8fNAw2Cm8R9dESSmdJ
Rziqp+emqI7mJteubVlZ/+vOW5NGKjfx8hDaiRmtxHTrd/cqJLNCsrkGHOuB4fkGSur60NiCakse
G81RkVqvP177SnqHqDacFa92bmWTUIzH1sJJTfpY/Q5fz1B+YAFrmuYN3XG80NtX/PPpUoFbnG3P
vx9EX9ktektyBVheTnG3G73ZpTKGmSgFqvvX4++/grL9id0SZ6+MQcOqaEaS67GgRo89rzJrEy6O
/2teUmcmhkz9MCa8c67+D6eGoPNQutuijyI8JJi+5rxF1wKfCAp4VqHdLpuBMgoyqgEOK+nozYVW
dz6TA48yFJjiEz0uG+2/k1Iqcjgpq6GpEqyozDmdXujTAU57INL8gxbXzGuvs3v36bimheeJYl4e
xaKLG8X0xvzph3VM0GDiRD3COXpuYEfhFm0EQtNEZFtB7hGycMjSNnGkbtlUzBtGwExyXm0O9sMa
Bxqt0SQwWiTe/6Vx6273zZqkcRG3E0iQzJ1jU7qFdM6DDxiSHPjaCytAJQqNn7Mp2vMmdwuPC6ku
V+TpMql6Fse08S6+Lq0OdoO/P0tEZysFyjBDcKVR65VGMNjykI3SuqltgWSlAf8Hx8yUAQUzg3On
XKzvp/ckt+Ym34/yYC0wXgJTvj1zoumCFh/mhlMUUyPtdzthvXq3TQQN0rhPvMbsT2rjwMFzhRVH
6MF1KLVKXEfpQieVuMcUa08DFfdHuwIoTlTGSvQSc4cEt2C6OUDcHV/kG3+ArgH83rqzi5KJx7Jp
d28M1I2RpCmQDhdNtEQgCyIUJ3LOXXl9gGHGlxs52li7NbAAj6KEFvZz6bd3hfTd3avgMJDQ4BUM
gYsraY6cdgu5sWJEqlAL2elH7P8+4n2ZmCpJO2FewWNpaSt70N8C41CigpVO7DPvBR0C1pkDBMUN
h7NIyAb6JQO/q5Y7+H12KrDIcg4emNeqmDJIxFAZZcREHBTZ4aW3WmOMQPPaPoV4ptSO2NHDzngI
AzOicDXVcDBqumR7TMi/ICqouWYtJO3F+XeXEMxe155XO6q+OYdu+hDygG9YASEnmlNke4Y7Fpf2
A35Aov42ZmhGqFMPXojF3g8pdpRCg6qBeGhc1axYNTxlyzFE0qONdgRMjGjL/pWABT6r3TYR47tB
rVdvCkMZ/6IEJEJz6fD9q6wQNN/9gjfvCHf/JWNY1TClAGaJRYRYsaz6OqJ3FmCB2cskc9LuoNQo
8pfvOscSNk6ggnyo+I1tmu/t5bcjcc6bfPpfwonRRcLKxJn+pGQcBSutnAlYEPW3ViG02p3PwaNB
HbIHET29x0qE+PZ8n/9PjlZoyJ5pL9z8CKWQLO/mCJoCALHSg2ZMBTzOQg70+X1ZNugSQO5cX3dO
33fuF4Xmwa1l3KmBcvoFiNBwTmkNIB7sqQmu/45aH+845pqsRZvvUN3IilA5m1GHQAvowXQFwT0y
vCDt4sHkqGGQD6dLGZ0lnXH6/H+p3+SPkKM+6h/t3K88/VbuhChnMSlIGKPZUixYmdQJbeOUuOv6
TaF/sr9H4/6Wz0Ey3fldraPH5MilpGlx7TC6Vj7YaPY0gZ3M9WqIqdGNlPIQrf3oMMGpj1j8+nc4
FEifdbyEVFdn6teGo2h0m852/xYYNVz+d3zHeMIVmaoiXBTF1loCc0gEe3zDYk7VrKhcctfVO5Ew
n2kCqkLxXz/vaB8ip6e2r9JQ5PDvuN/jHCwADp9ekQw5M9IdAJaONQfn3LPqmVBhaxCMIJULdDJQ
nEdCG8IohDvoZ+2Li8bbPiM+6cf8xxtUlx+E8SX9OOrYGH7tiK4ZU0pS0CXf2rOXjl4KvBW2eaXH
iGj0sqeNWjMYNyyo9PAnQsKdEOqhQubVBvhFEx2ujia/og70w0v6QpPWWLX8GnIm4j91Dfb24FXB
6OAfYyj0sHdMzoAm2NlMN0jZpVY2qrfsK4DoE1i9ROpm4u0PNUX7EeZBA2xp9nYpkd0yFEluJbUF
P/5gvLyT2tetigEhvi8sBWAIIjeQqFjISX6Ug9139/gNWyT/G7AZFP7L/KkaZoRD7LBDcAUqgUFE
3O71MYSLlGRz/Chf0jbuSfvsAiixBO1TUieGl2d8EJH69Wsag3XcY+3+TOSGnbRJ5W7xLPS2r5sP
YldXxG36ZSqQEruZGtmmgpaVIdzCZwBOfsJItqtwJU+j31HzZ7BSGQPIdODk8R/NrORCws44XkZw
4k4ghIuqcdwaJiURS0pOoX18UowwGUOgg0wNKa0FITs5wYv1aSZbYfWjhzZqtTbWhROeM2AcCU/M
LDAapLJHV8Xbt1bzWFroWEbLucqoyh5s/zuFtag1MZ3SuCjWuqKojQ0IpxYAVrURhnFc1ddbeNga
Z0PEDRHBAg7hhke35M3tTKcRg3/8T3jDSH8Mn/jsrA0ks1vhDIs8u7qHKDkXHbwxy/5S+ilbvBDB
G4xSpEN67d1xeTjXPqkiv5ztayR7C91N0sT6xpYYe6jLIUfDrhIse9SGmnIyhfK6+dwZ7PD5CQgt
ffZVdfWId048ZUX4IvIz955y/4yD7jesTlLTvECHkNzfSYHRcfuRREP9m4twHHU1GxISHgwa+mco
o1Xay6LLa8aqYuS4KWU6sQQxu1/gmBQrco1FeXc4OMG1yNwVGw65rDo98VVb5wAhBftlnSO1g1id
UfJmvbp3FZ0jwrU/2wZWTtFtMSEHWGXH98BG6qNHN4fWfDP5vvgCZkE5K2R4kHaPK5jH74dHWFMF
str2QFoeaPKVBCRVu92e91sEu7AJP9yN/fvxUH0umZJ11fd4Y9J5xUTYUgePXAHhfwEUAospQFwX
T+FnB2oaj57ntRvk4s7f3GrxoXTCwN+P7NvhbBxMXJ2LW/ZiO5hZ9Gm5gJsEK907YiX2GmjxknBE
2nafp+pfgoY11CSoA6uQWemU+TXsgr9hL90K8BTykTnTdTyQ4cpyMDfmJ/C2Ls11gzHrBK3tAdHX
yy1gTmI4g3BoYDlCZTVs4vzhJmb5/perOWJ20gR7RSmVkL+gTtQNWs5jsvUtQIr7KRt3OLzYPd3a
eEq1Tn7z0C2PqzXUj9q9xjeEq2gl7PtvYYtk/HihTCOmjojxcP+nToo1PypkH+Ln0H1u9DWzMSUF
3dRS2jv4lysFRv4yZOcEMB/0ELhA12eL7UP/J1ulZDnlfEb36SIe53gWM22q4L/O7slm+zE1pIpV
bDojTQC+9JY0SunM0vW64vAX4pFCPhUnGqbWWObA/SaNGS7XgyNyQ5tWJnLA4WDvTOqSxIHmmyth
H2CZw/ntBhX2Oo1bnL5aQXM4LAU6EtVLt6NFAPybaQ7bpr9lrA3HbLY/rGLbQPiI5o5rSC4Ji2tc
VyRbsJRSLXXV2Yaos+hflEK7TCoHnboHIvrCf9XSMC3FDscJk2Y6i5cRWPDtl/gVLbtukmfta8B5
0fSgnf7FwzB3sVvWSHcFehxu/u/xyHuVU9NS3VOr1xHr4knsUzPxJyUnbP7pISBwJayGTilzW+L8
bc+DEHC828o9cMcDMhHfz4OCH0oy+/swI9F97XMdHv10uBjWqEyDdhYeWneUijPcQBuPTDaC6T2E
q2sUJsV+x7XBdtMl5XdtDuYCWIyc3BxmqrIjW5c8zRGMMHMDkqcnCo1wiKbADtJw0n7xUWDmwN2+
YWLOj//PgxREhtFeHeDkRW7w1/xbsutHHRN/lA9i3+FETDX7pmVlkC6fUT5psqgSCFuekLHm/otI
X356dGD8wYUfzGArDbqBKpSsG2sC4EENfWv/NldcIzmr+ygHor7rU66V54ITl4z3qe3O6IRPBFCP
nNAcjuqzAzWBwyPZCBrzSN0pnLMvNQwHAWZi7hqGx0ggLCIEawHlTW3AMsKbRGHCWTs9iY8Dx1bs
QRBHYqBIvkDM68se8+Is6YC2r8dfCNnC8Q3qLoi0wyVZzXeFPjiKQFCJYsZ5HfQ1Zt+b7/nRQ/TD
CeJyIeWjPHbYo2bAOwtszNkm0coaCbV4zwq63G4JEXBrEFsadil7+KbgDo2jyelrLbTMZQMzzzQy
3dbPGokNTb8d3SnJUVyYGx3ndr51je05E+yL8igChYdmJStvQS7AH0ZySeevdx9irsZteEHaGbT4
m1V8l355f983MDyUCP2NBDZF4vCjHMFoZ6IG6tw5SJQyWyh/lWdOF2LZQJxdwk2JQf2nqD02+vCg
In96i2lr3LSHGO5K98+V+9bJUU80BnPWlnu6VaPOSI1gIo1RVMarn0E+wdRLEkL8jqshsgPp9V26
TT2bjXqTNXNlEazPwc2U6a14x7NCT4Ric47xoD404+vBBL3YD+9H8xgTWViqVgxzAUIz/D5v0TeP
VouDmwtxtpp+WrlmzqJaKl8NvFLBNhFR6zAH1L3w7VFwIipjV6N2QTCMuEQdx3ZYZn9XTo0l3YRi
wchM58pnPsF/QrbsM7ldjt7m3vz9ioLN2BWZSkTtVuKY/iHqHkTT+5ke6lzmPbabzjO7Z5iafTxI
DCKZCRIxp4YLLcdVaO6qfjM30TkEJwky8242qas60SiBoLu2G39CGmie2ZJITYvVNQI36Tglqo2f
n/NldHsEoV1AIOYRAvnemcrPM1U4ZahXYencYreP9Oh71yhWPQRAMr48jv+nPymDF1wQtqmeKFy2
EfGisXvJXMbixxKS/8MF4Sm+tMFEU+oVRL5G57sjSiaQUp6SAhXYdIRQbE7MOWbnqmZ0vBtDv2wu
asdF5fCdWgkSqLN+Z07U1Wx6k81xxQimzcn654C2XI3GYSzt8ARe+07YE46Gh1IItNJWkX3Ij1LH
ztFOKaKhCysgJO5wbKacu6DwEuAkJGjwZxwqARfiPi4y1BJ/3viYV64wm+zX5pPAi4BbJWwETrc1
sNICNU1xxVfSdQEbwXyABR1jsK38N/PQgxwbU+NoFg60v+wdQaiHBVLr/sZBZLmAxMGMPsVOkZpS
LL23Ox+M8c/H3fqLO7e5TrzuyU2+LBLCevAelCjjYNjy1RUc2daPEY02IwHN6z0Ba20lvXYEi3dn
nebln9gSayLAmyBWMUgRO8CMv+Mqh3MlAWMnmlHFWs06F0ut5J4nfQ5BDwP0IvOMNUrppq27GuhB
kL6DHGDqRJ+y7nbMGASgVbQ03aDPSzAzTkwNu1OkY2rq2FlcYzu6VPA3ONdZPHo3qPmn+6UMl3wg
Zev6cXkNATGbhMZ0dz+vGQrzDpwJp6EWh2+dP8eGlis2KQNm43FLqkkqe/XGSLK180WkgCE20iFp
dKSbH2H7eefdP+fDsQlg4PJwJDtIQM5N3IGNvfhPcbeMto/jUHarGJtaumTLzQeQtm6u0lGjAeCV
yv7Mb0GHdyS24zQCN+032xPqS321LFXtRArPqkOB7bdLMWAVuZx/yrteg+4Ep4XSaV7bvQZJjrm5
DePQoQ94BH6ZoOwA8Ch3cbZjp5tt5G63X56Uvi76Vw7bNTPfwjqHq/AX3ovJlIX0Wc8chycjwzD7
t4A5MRFgCzHhE+MjbbFyymL07jMomHjd4jgQ9iiNuj9cYn3Ppmy5ATuI1kj88v8KCODNTnXbftyT
2p1WMDIONX1TAUlOwC+X6vCuVdEIgIQtCa/buO2fHbVPnbox5sPrvgZxCdUxqMdsZkWs83gIrgg7
kjFabENoa+Yy2DwYH+qNjnunxgmx73AbbdrwZDbGWf+xoPnNm2y++O26ZKQa6lHikY1/3MWRix0E
PR9r5rcnYt/oZ6TbiovovnuQqzQuglHTLhgni597fWKkjoqbYShARO19kJJPT7eHlFAUrfX8PurV
TQMmXoGgA2pHfZCTHohM2TCy//dndNrX8zhqB9ZMyWBXbH1mZQUzz/sCCcaXkyVF+sJxUOKI8u7G
AiW+9y/oXHu5urKSCUrOmq3eYuaIhXPyZJo6RDWKNCgRkLovhjJ3S9BMGcJavqxub+xV1pvGPAoJ
09SzqYHyza7eLazJ6JXKDvWCjyX4f+pWrkD+TjvUYafLf79JkAhhTt4uKgRXcH1UbMSOM4m4wkma
FMhPNmFuU/idqkAkUT6ciMQEdrXZFTRqRFyNAgdH6SzieULDIwoYYgQe3esDRdIKsHO+uUEye1TN
3R9r1VWp/fdBnYLL2fiRPRJelh+ekVG+o78pBrt5J2F20U2tdlI4u2S1SFF6RNrqN0ZVJs5bniZE
2Iq7j7cwdT2ASVQkd0Q2wji6RclJXejfWZ3ZEYJkJ7TfTMSdkLs2vWMCoeTGCGnRlNa8rISuk5Ql
vuHXn1MFNEx+dbxXVoCjzTGBaMgVt9AyUZqn4wi1SBOiyy9ZqL2ad9qrpxOPGNIkaoAi+y+uKdj/
znHEsC0E0hV97oCej0IVNAu6Yqq7oDqUfeRnAyckJTfASmdBUZNWWh1F7SJN+59ad1h/rXRG+vjp
rBYjAo5d/zjAqD1t2xcjqMgt2VWHSrOpAfC4JKZZQJOpHnRmvgSsfurLOTLlytQBhzzlJ/18c6/S
kFcxmtzbtEGyeSlT7yAuIAggDeXTWP5g5UrOihaz6b3zUQ7aeUiVM5LQtHB3buhFRkRVcm6jD0D2
eKX7EzkWjptzLN7qjqye06hRFdfwBC2uLQIxS21lJpYjVv+8mrz+3yFNItlN2gl7JTLoChEfpvPN
dEGxuGrOAUkw0izKVs+6wgX0REdxwUMQHM/f8G+MiQboGjeWyC5SyYJYFBRpY4qqneedd53HW2ag
BL7uGNNU1e2kzwBGOU5V9r0DLKOC3NchxoccHzuHxTcuJvJ70v2mGgaWMW3KFmzC6IzZ7b4l8jHC
OiRBmsJIToOK1eljmjVySWtE4bj9w1WaWPgaLBgfDzpx34btNg2G6Gz5z861Knahj00gbtFqr46z
hMPQnB6AxmPwmifIP4UTRx/m2EMKAeVfkHal7QjnMTdYqR/N1aySUcVkwus6TnfOl30WpI94vR8h
PvdaHnBIivC6cDiJF0If5xCV7R4ydAAUjtAP8EsrXS3T00URGQ3lvv/ptfN9LYbgi8J+WllPLvIy
9L1wzbtvGfdaG6AOGw7vPU1egJoJ+4ouCAvHtwPGetjgMWz16ka+9mfdmcWVYUI6EN/sh5zqBSA3
9goyDSg9fNhiTCMj4PUP1VCn5LsvfucKinubK67FkmvwbRP7z5ll/e+znPVoWDOyrH33VCPQl/tG
pFFYHaV0MXgSyZvxjERLVJG1m7XBI+WoagDtT90A4gV3dv3JcqS4lUd+dUVQDtoZ3ReccZK5n7kO
OGAiQ/AK59l3n7dgG+99bL94nMp7Q7cW1v7Y/36eudr03zAZThKZ/mCoN31C9VHCqMQnPE26BFMm
cbljmkpkmH+LQombu4yoEF2ia6bnCNIAqaLGdZcUetfZ/EC13/1yAubG3RSnS4IUk+H4cK8f7Xhb
fkzMMAFR9vc8KnHEG/OyFy7wnuaTu1ahoLCihUZHweskDMgPtNoH+z+atfmm6LE+FXASd50sZsb8
dQ++mmN4XQK/5eOvH+yVWMAgAzXeVDAWLPrBU9G2mCp49atszDW+SnnBdvAekab1L9J8ncX/t6bF
q1OiMsYmKuSjjJt6ViR8E9o3haPJky3bhggM+Fpr5pM0ItRrNRp0aRmcy+XUnBpT/Sq9Z3iPgO+f
n6uzs7G8KuFGCvoVmPI9Bw8AAfFSTmfWDbkaNV6cMjJmXEYKmFPgg0GOge7HtDHuZdsDiiEFGFpB
u4PDrKr36TBEsHWWvOi4NQJgmM5idxYEV9c5SpMH83ctYzeb55jGpIIX+P9s+w4kcC88VBydSxO/
ODyyXI0ZxYDf1qLZHH8CqaACA1VF+0dYKWg6JFBsrkKJYtK99/Cs4a/gvWoDfJiDQsXZdfFgk37d
qSylXzjMjcSejYfSSL2xaREu+kN5k1RI+PbBGygcNJ45V+J5DhZYNP3b6vxlWoxm41YWJk02frEm
ay0vuw7bAcZiDEoCC5QdNlIXJOPxsCDh8wiLWRu/mm1luTC+PksOIAxWLZV1tH4QxlqyJr/mVrN/
Ob7I0hle95pI+JHY8b9Vo1RHtmT7VugvLBvbJ9OwQ9t75GqoyqmEqqFRxPIzvW+bCpWeACMHpDiS
CDa48WwhcwhfMloZ+IFXaZb8PHwBcTSLwA+ZPhqahIZ1Ec5jWKWB06xL/65QTlrCp3JjMFCJynWQ
C57ZLG0v3pDIpmf2KMS6HaXK1OAy+emAUKM7ew+qqWNB3rOQ4Du3Kuy5Tc2S+QhREvZpJB6bbNZQ
+Qw68HrNab/TNBj+PFIy/D8aSY6YFKDfhQ5IBMS0ELFC480xIgbT/6k9ZgldbbKiZBAF84MV/iZ3
EeWvpQQ8n6S32sK7CLhajIH3oo6fy0UFc5/3lLupVdg2Q0SSIe2U0oi69V6xMw6uQ5hlQDTkb7sk
2Zr16rKZWSBTAS/NlPz0/eUgjRVNyoPDfvEtjtiNkgyrJIvBhuf1WUdNczqKdTiWOgE5KXwTvD6I
azrGYxsJgjOTqkLJUvPBsAf3GEwzqEniPR4yifXTXnRI8V0ggY9j6KrCFKJlDWY8jWT23IViXXgO
BBtJy8KfHT6N0LU/w1Sxrxrvh1uhFsuWU62zMnCFDfIWIystNi1NzhxGAPNgFj5JyXsFOGcWWEfW
hCt//gAhanY9Or17yvfifQwU1IS+X4VSVBC8VQiYkc8bxrWKx37UArJ3VlYFgau7CgawPDKZZiwK
lsEscYE52FPX6sd9fF3+ESOZFLNxBQNkZ44KMfbnFMWpUquHorth1oJsXmthHSPbKcNPQMYETefp
rWOI5d+et33xy8y00HEkSfpn+1NeqiC7DZyiYc8CX0/1qTfHW4nydt4EutykYWkzgB8jQFvYIFSU
USJ22O5+KkcClIgQmA8QPFSzvHT7NlUDgoTYi8c8+SDANWm5l2AghHTOhTcLlHTwIGm9vwSxnvzP
hCrE0ZE6KXoGCbJvDA/vHVdhvZM3azkRNE+JxMRZvZu1GcZZRfiLX/iamg/OEkvB27kecvDCxj2x
bBY8ykCNuovwBPsvNg0e4/7Szh9RffRhNtJ+jetnMoUk0edtsK+t+WSCqoWRJFBHLWDhu2AXhrSv
AVkMJuSnqdLHLJVUOzkfIwsdi6zwN4tOd5dwcNTt4Vsf3o/5b5MM4y+huReLRnoQN8WehRv+oB91
0zGe+oVlSGevjxgN0pjGHlqHgQTvPehcUOK3l5C+ksfUL+bQuZK61dnamVip09JprwO8rPuTJqgV
Di8K5xNbn7bbsfkPAYggpH4nVWQMeC0DLwutI/QWKQ7j3C84QbHrA2muVKcswj0id0h0wPmNgiUb
VJhkl3aMFhqlHAQX+cP3b1AxwaTl0cc5r1KoEdJTwB7R7blfG5b+laJ/wZbIQTcQYrHEECY4DOPx
trsEaDwYAcH18C4wJUYCqUytFCT7KC2fSt2W3lEUXlk/2oDPZTckaFUg5jcKI/OHxx5rvxue02BH
1Ggx647y0uRsIZEHmWV3TLAmNUyk3mjoHmuy+6aYqfnYH4OjZCNLBXmKa5Y9KbColnZRsDeU/92u
K7ZRaBXRhekCFrNAW3wWheHAckKxLqw0P0o/+TCBtGi6Y780R+7o8NXpCJAHZ/jHDK9Z5NbJj5Fd
1u0DJOjn5RpIWBCqx/kAcsmKXza0v9FWub4bgoombvuMHTq2TT9GXX87gI4I2Hw8IE+lxbaYWEAR
oM6K1dEo3MFIwvYg5brXysVYSiyLMq6Vahv63xq/IfXq7aD0PhSu0D2G/bilW0XPx3b7jVuZ8fSl
E8KhjV9FB1+1uYakdG9IW6v/TFk4+9lYHBopE0FQueLArkBB0OTgNv76oJ09ZavLC/gRCa55/Tjw
6tyg1uqyN1Z8+5AT5XQPTEgBV2tVyeQDt4vvpXzKzUWtjbqBErBhzQkjtjM2EuFCpG7VsYGTfcJZ
4BwKHubcqATMDcTYLPMVocpEMiTYmp/6RvI0YvrYCNGmOd8sj4x5fsH8h/e9a+1FZFw8yc7fCk85
3OGY3R9KkfZSkjf42ix9KG13ExcEO7ae15V4p/9/MN/bIINKcxqpHTVchLrLey2rbh2/5kRVIaDp
nERqo5dQKZaT1G2xy1/o1D5pF/nx+vz+qutD8K5CqqNV+GzdZHAbUyWaiA3LKu+o8xj4XcwFyWzE
SR5bxmq8hVPDHR7M7Oych3c6+E2jOouBnP75E2vdsZH/NzeI6M94PqT1pF2lKu1x9j8FOQ9gg7Mo
vbYuFv5Bx2P0Ng2nQegwqWjUpVz53Jvs8OfHgpjTQe+F6/2j7m0aAogRStncBut0QLf0CUo7uFhb
5MxRo5SXaP3Ecz1KVGTRLpkAHMNBNopDk2dfOEN8ij536XNCDAcWN+Fbsqt8cEhWkiR36ONYbpZu
QkTEA8dWkopHLDSM2m53J1N+D/aZcwKW+YKJR7pnkyDBDDJDbT+BvQI8YXtcCPsCPEm48SvuqPo+
mllFcJqfN5G9Czar01ViH8TMm+9GDFLB+mLg8YLdhz+Jl1GPA3MeyiBVP7B1RnSLoOnvjUVNOL1P
d27cSlYRhB5vsfZmriHllBN37LlSBfSXsDoAX+w2otP9Mo/EtWiWPozZa6ayohsZXuZXwjBkozoj
V/JuigSarlP7bkTt4nB7WeK9TQzKwy0mB7Z29dphqGgVvB87mRAHQki4tTD2i/QE0NxMsBgM33wj
UcOSvSZuCT7F6mA+m8TfFG7N57T2urOakbo2IgEW4KxAth2fRbWnUU7aWiEUZrKId4lAdFms/AsG
tpLQab+NleaJowZ56NhXDXO6X8pOBSAXG2XU3d9CbhiEkGnwVYLA8qIqt58lPjWqtJkuyI2D7rB7
AWPk6oIyR37Y4iH1E5QPZWgw5SpgLsGV9zZc3cpQoOKVVjlnnJUcOPgHRGIHXbrWsGLRtknAHt5r
jSF00FC+XlcwELFCkVPvD2no3+ZKF9yMSPS36ZNrFyTgzwWXmbXGIeSB5RaZbcU25P+AHYWVj0Ol
8iayCgdWO6GfBwQ4qeWYrbTbFyptQGEaA3DrKS57Hp2qCGYjp/gEiSbOvQFwQSWfCjt7PABLB0Nj
qu83pOnQz/aSK2v0Nnim77L1hERtdn3q+jVEIKDjLPMPS6NxajsHaYNQQLX0mNYMChf6xVTkm/FS
W49qlTWdCOS6XqGVuAZQ5qCBvaPHz4/Td0KQiUdOH8CfPs94S1Xm12xzg4XeTsvxWkJQp1J0kwVu
BWs1CcfzkFF1LKPN5amFOOS3/lrCmkFkk2I/C+c1i+VnmiZ/uepu6ldh18RqBImnDAgWirzDo5QR
WzPw8+0lbdhhpNB0FRAM8F29cRFiXhKTeStz3r4Yg7y77P2wSFGwWiRMngbo8S1hPGLAYpbYe2uc
9AapV1jZ4PNWo7+Ddy7Ou54JsdmtIgMa4GmMYDReq/t1osbGokQWe9XfpYy27nwPOuEMlsJHUW/D
QNUeY77nLjN4UcUdo1Jvuj4CLZXaYKOsalOZvBl+4nFLjT8JIEBID8wLIOlhiT1mn5E7Q1hKVKrI
2ZF0pLAF5+Zzq3Xlwcswx2nljuVnLuCmrOP0NJXo73qmdIH1oMygiOxteenE0tFvZza2rLph31Y/
zGYaToysSvw6bvcHw4krFPEft2cXcI0av+anfblf8qS0CT72jcVD4Dog73jFqM2X+9ku3dnaLdMu
CVjcFsY9QLu0Z6g/yotNd7nk88lIU9A/8nKOlpJZIjOS8dpcipZ7gjrvpDNj4qHT1mmTTUwwuFpM
XjNrwUzQBwO4v3HaXRY7BXiDNuxODQlfREYxN0orypARAAfEalKOUlblv5PTvQvhhCH8+HgQT9Ye
PRc/PySoA6XlVjcxQEyq0d5AW9jJCmocuAUgb0HF5TGwMJ+05Af13EBz/oosKxJqfG/SLuEA1cfZ
bgW7dNCBQy9jdegdxSuYGe2qEIb2UiGAvjozYTKNqNTBgc87CXotVAHjzxAnY0UgYTdUT9UR8aRq
9HAHnE4vhX7Kl3xw+zwcvwYTrqUxnpgXziN67wnk48U0Apky+CB0U//WnE/UnqDlWVlyNskVVcrM
flCjg/USTlrFT942W/ymGT2HPYjb/n0el6HTeUY5tpYqKk3/5JGNHg7M9SdzbsuEI0aLalq+hbVz
rxkYrXx+FcaMqCEz5C/fqB6f5bl4zD0qBBwrn8wj7MLl7zJnOrUyFRYq9PTGgY1Yy3xHumbRnQ3l
b4ZEoV6ySXnpWo24v/iTHJBu2QhTllp6PCw8czeo2BKl/rJtZVAItZLT5eTnJagXA5ks1D/WSh5Z
pR4lCcKs8YvzUL2TSb2kntrAYuZWcg1fGJP9nVwUeymOXwePcT1BLFbpL82GmSwspqLzpqlyv9qs
cKfdF2P7ox/GX/nEt2sH5A1eSrpLXHCB0AVesV+aVXzeYfHjsWPnDdKprmBw/xFxxdr/zEnNmLXO
n0ib0eRr6r6GEoNrAAVCvh5isOLgjSYN+HpLXUN5lEv9ykqIVGMg0iWHuu1rfHWr7xB37GLSPZ9/
cQgNEsK2xCjZWzrSKJRpyjAATJDsmogduKa+j/UCmz8GBP3uBknIRdIm4m3z/zvwtsNT1HNjGRMZ
fO9a0VQ17zO3zC3P2W0OG/lKFWof3e/YCe5YOUQ/dJPLcuzqKUzWqJIXiKLSqR6Dqe0QHZ4pg53r
ZRfo6Pq/SgBG+2dqQEt/q/05xWowt/DZl9YUvgHn/5nOCjP4+dTgQJv2Qh2ADqm2jKaEmKyB50kR
5FuGEicAIyhYZtspzjhyc9GHqod5taYoc+1q1kA6378/wN3mdFB8nBcFpQ9fXdFZWoizjgRT5Fan
BDuvknZHgyywgPdby1XuorTpYIjs5mGpEaAZs1rBJDsVoAM17tsUhHBhcrCLv/ScrQKCd0IqW2nj
3KNRTUXmHwafjaRTKnEthkRCTxiCyjji4vucQeAe2wWhev0D/CLFEe8Ge+K1pIlzl+TTVM9pAwtZ
tkC2u9wa/3KbCsoB6k/9lRBLiLYSqXnLqS6sMp2TSvt7/GJwv1UGnhmFXDGNmy5LZR8q+Z4XgdWB
TKlPi+ZvJYaq73ozI9ewf4FLFOE3z+Q+tOJ3cWMuT+C4lNcqoV6WXhARazxgkzQCRl8J5wYVVHu/
j0LqznMXbBdWIR68ujRcUuzmVaHDdwXbMVMyOSmcGRq36H/hpWZIn0HwIkhi7bvWZ04q2fgcZl1o
Fn0GC93wT8q/uaSjvlQB4Z36kqWt/zHjApBneFvjyTThC4s+dambatSR8AoDj6zxyKxpXXQm6nJJ
nZRr8NfnmfIgpTT/hxaq34nUkOOFVs5mxZP1OsHjUi2sPXS5jSvAUZ5lyU7UCJ6Yrf1ck0WlOQ0Y
sCzndRUVYXYTcPtsvKAqP9RdcbTc0hpYwM1DTLlZk4aeixAJw8Io0OIm1BG1KaRqIFUvK2HYt1u9
Li6pWNoCXHuybuOEnQXBW8K3zr3PnmGuSOWL7lcr49vJVywLytayDA+5HrHjhBFku724teJkeCN9
wPTm2eRmVd/DN0BiHaUF7UwGlk+7SJo9YpHxAFSKZI9M6vkL1AjF/KiQkyBT1OCkc5CV7c+LVKtm
rQpAQ7DTnirI+D31viik5kyLVK+4+eT3krTTyXiyJ17AGmHNUFb8kZB4fWtFFk/mkAoxtMy3l8qJ
6v8g4xK9KSuLY2SDydUtUZGzJ9LkHMaJbRDVynpTPvGSirFRReo8O8N+Nai548a2tNhFbjFK0+/0
coz7a+he36D1eJx5I8m4WBDGtV2kjI9dJNXlaJN4mlyMqzpSnMDqQypX8glk4jx4UyHi1H17NTa5
GDHNsD0bBXoJn1vt2H8hRfRPTkczXvyu+bfeoEBVIRpfirrvoYhRa9Qv+1puk8hygqA9FfwJuM9h
w9YT99R5cnW9ekcFRoCfO4te4mZISVsSyRqyvRZF+sr6fH/4rX7WFlFc0MHxY8IUV6qlift3OqME
YJQtwtqmkADI8x61SD3FQ/8OChECI+J5+P9qyV1CapkMCKLE5alwlLryULd11eIUDelUPuwPjLhf
baPjAhMGAynQC4CFsYuKCdqFy+JYduLtAHsbIS1/xgXNm7mdCEW99yMTlVN7whTseVdR4fD/RjF7
u1f68z5K+s/syZAI0EJLlHEO5OZxmbzqArBreTbZocR2A305V3r6X38sC+lzxPGV5pKgi6PRI1Lm
1vzrBkH16xfMtvhwGLCbkfO7/iSrjajFEEA6EtJ1rCoPCP+IiurByBJNdG83Yj+bX58byIIhZW46
FeMs+RsWi/xNHhfM3YGMF1yBB6JZihWQiUMiJdY7W6jev00uQenmRwbbMRbeT+1pP6+x7K64Cr3R
sICMK40jMui8QxdRuPpPCvOmPUTofaAaK1WeZY+MPUrqe7Ue8UVyYDQgQqCkEYFBPWHBk7v91qJg
ZLTGl1wztjFo4nOnKZ+smzwJzMuxBM8MlYSmcX0dvIqDMJItgiPE++fYASUlN9AtZiyiQK3pe6rY
wcOqapYFCeaD8nbIBhGGj+vN5IUyt64Q87FJFHTlTNeTtasVcdVMoRXqxFE+YT041B2O7SiRLoQj
Qkm7QOuJjVi9iOXqnBMsMm7GjQE+6IZoDrb2KabmVj3LJ25QeGLklIjiI5N2o/qIUizg/HRxVOix
wQ7A+Rcpnn9VU/lwJ+U/i9VU8ijHZo8keuFvNOdrfTBa2UggcFT+9qvEBH53IT8GCL389uCq4YQR
jJ+1JLYvIX8maEJUzVJbykBUi16xDWxOqJypnhLnNHC9Xc4+apSGQ51pKboGMBHERDFAiSKVf4/s
zc4yJ5osQHsOOGtknrrCoBZYR8Lqavpwrtf+20q/vy1uuJ8f0gkAn0TY9LXKO6dVouBV3yGP8FU5
gshBQD5cgEpBS8HNhw83dt/s11U9mj7MHF+nLSBmTqvMNAmLJIbqiTRgjlisq2+PYocDoZ5xBd8B
YuSc8flhgJelsTAta6ln3CiO7CGKonQ4vem3sTgumkPTaXSwUzzt6uRoM9YP7n4S05xl3vtREM++
ElMAD4szZTXK0EmkHEcrvFT92Kf766lOlf0gwk1Hj/M5SKjlaOzPbClTCjkuBgkqO/hKS1VZFhOE
Te57SM/sUAi4JQS4Y1dz1QBdrAIn+FnnQ6Ex4IS+lxpkhKUysFMHVsuIwCSkjc+t0CAV0zxJGWYw
UfX41PbKh/7E0XVVNa4IemDEhLErmzR1kLl4pXIZoObJW2p0986PcRCegaIG6e5SbguYkCkgljDC
6PvruthLvkOrVAG9NWuvdOS4txq+3D4s1KHMIW3NSu0RZeK/1uNED1bjbSFOH8xdOC5HWJgnbnHy
Fr7iOtfd5tr8gdhMm7CFXk956PAERIYG7VX4esBMESTQzjnCVuMWgf3xRgHjoIKTYB0hpQM6zh0R
A3Ru8FPYzKl+/EiXzbiJ6Yz4BVCAP94U7AyThExTwNIvH4jwyhmNBtCwtxWyAcV6i5TPp3INxf4x
VZXkQE8eGeB85Dnb6lt7qKYhpaQipzaBNJo+UD9N1Vwzpk5TmWba5ny7r7sdQLgTYegIJ3y5r+I0
cZG2sJ4PCnP+LvaIASZ10Fcz65VTGkA2LUcRmKuQfKJw4Hw0AYlYtgg6oIA7JRNqqB7ChUyOgPeb
0msb3J59TkDruuUtQt5aWKtr6yrwoObA6hq9fYUbn4PKd+rawok6wny0v0KDnGyYlNU1A8FH/iqb
ONvB5Uy9lc6Bd7O0LSrBH02lqH0UuBlCe1ETnVk4KZrw79thMp9kSezFhov6OkKPDvzak7qH8/2q
0sR56pUD9zvYGbRW+GVrKK/YSLuewRJ0PgEhgVCyx0tuIQ4vezdV1ugNRkyGCApeY23ud0loyFSk
7BP/VmZnzJGZztmFfPeY7tNBwANTsL47yjQHZTJJ1SqTxkgQ4qhD6aQc/lFd3VYXa94SgFPYFE60
zlxQL2tO4jqfqcxuQoY+gK4uxVGj63UD1hsxY/Ho6CdiWIYk5ECHkOLbdhxQvR61nua53uFjgumy
/DhOPUF8VCCaB10VyB/OMvJt++Pc9778OP8I8RHh8Tf0DyEGsE0lkYFciWV40TXHhNclpXbMWPuD
8ZhLjzVZTKdHYaXW7My9DbFXUHAIwoOzpJEIEKFysKMzn1NLnGnUDamy34QPM8cG35xAn1i5/kdS
1wLcV+yuI1y23vgsvLW4SWDA5p2DeCymhPkI2b+b2BYafNkf3S55xI59E83ISt52McQDuy7xXdVo
FUEnfBUOugqDq+Rx6otiyPyVlUYg+BDK4SmV/TylpvVPRfmQCaX6MsHSF9OJndprihAHNFfx6Ywr
enKvRSQcN5WtEAnao7BzlCNfhpWFdZfdRu4tTellacc98B8f6M2EGD43cgbSj6Pkx20hBv/HIVOW
2jPB0llA9hIBpEUirzMond472DSAVodwFt58RFvaj+gtTPKqhTKi5fQwRbPGwbdJxAQi+SCpN6hC
2tGidqvifZOArx+ETrz4fPlEYzL7ceEGI9ovy+PM3VMP4ZcFV5RvIngVO4AL1u+iVzX5ZNvIq0qt
R/KSo3/SFveNa76rPEDE2e/2OD8Ua4mlGgKHb01uxgp+bGTP0h2GrGUmyPayzE7FB0OQ/HgTTica
9lC3DU0HiTwhdl/0NnGREb/fk/ssu0DaWGI6GajwJ65qXYwEivUpLO/Tvi8lCXKjscy/fkebwBow
gxNUoTFF4YsAQ5fqP5Bn97hl+TVO8AO9uPGHHYd79hQak9JNUiVYVFnKcmjpyeksxCkN3NdJ7II3
J7NfXbpQdo7EpDwYoJjV7UVvd6qia46CHU9sC1fYV+LMTF2+9wURQ6JBsST3ARVbAHRNGRg4jJzc
bePZTgjYT4aCV/X3EkYCn0ctKa7/TWpyia+1EGYy90No6+5FZNuNS/VUDLns4m/jpJzSGXhpJKsx
KYSzK0BCpSr8ljEVLMVD1r2o18cBX6k1Gw+azitVeYTr7IYgoHXkRuG+oYEEA0I4RdrbjNKQEXP3
nN6z4oNEXnwCGvSl3NT7NKGF2n+hqOCeeS6tThxViT9LAtZaZZS408/ou+/a9ipvBlvov4ihzsP7
bhosdSnI0Vsfs9tUZfHLj4rvURlYxi0lZBaC6HFexewsysx4ZWxplaPErJAta/UPJH4KuW7zqHnc
E5SQMl0jQIAIrDSwl3w1ftThTjBixY131m4G+ipa/KjQp8wnquDsLGgly6XoeWvj1roTGVSjl97o
mdxtkIJjX0uYSxzYLbzqjC1B83x2Uho5n8SGZg9DJiBMSxi8KmT46FkXsdOk0uIjUPVoWNPMwdIC
JdqO50a/B69qG2wAtCa2AyP78BKbx1BLX28sZayK0YK0ZOvke8l8CbnP5fugAx6LdUjue44BbZlT
xheKB4/cb8WFQgZEiAM5Tj0Oscfjt22KdCaQF52410ZYq27Ro9sN0lC1HJPUBkL48XNs8JNpgGlt
I6npDWlzkdoJnIoShImQyeh+deGJADK2f1G2vPGsTpxxF4l3TYvBszj0uMAu9eSwpejN5uOFG050
FDLGuTQjmq5jAHn2R4JVZ6bfI4rqBTKK1/HI4JXRvFzVFfL0h+TMPGlCB6PWNDWa2vP0pZKlM9QP
6lZy+oNy7gbMzabwlGjId+MKivNCjdfi/nc39sAp+dRan0UTmfmRaLnB8/Z0oTzj5q84ZkylEFaY
R2yWzgQu0/FNZ6jlIxv0OzhjaUCqoC9mBZCWgfTHoOJ7exSDzVa/mq95m6DaeDc5fO0Qe9gkW9mg
yZWGex7gPHdXLuzxZ1znSsQTtLKjEWe/aA1QLmpnDTNo+8QD/C/9OZZK0GCITLkX4xFlKtSJPxMe
DQyHAvBA5TziqoAqL4xwDO097FoVqRgGAWfhC0XlMH8M4y3yW+7m4pog986bJD5N21rG/2Q85uPU
uMJQY/JoZM7gcjurSVWsCv0ZhasH2uDPsPt2gN/4bVek2gpwBsUAzjKV1RWJ1viZdJSPKuhJHOb5
8Hkbux/nEmA1Kj6wQ0HUpUUSxv+sSjYwBm8bp/iqGEUIrii+ZbQI1xTVqzkFxcbjK+iVfNyrYphw
RYEcDTBdjT1KkYC9qf3H1gNy2mZktOo80CfZuZAjWCAwLSv8yKbi1L2eklJLj2Ni2RuzRA517ic4
d/L3Wzo4uGrd3eWLhgypFCVRpXItFQSv3qlasVFkDLO/kZ6iaGnbjDCpL5vD9JpS1Baiqjc18E8H
lnwMsLzBlp8IGB/UB6q54hmIeF0c4NZDpWyiaYpXgMKyJc25kssN4T3+EkOLKVU+1qdzd0GZwmWi
3sdipmf4lq6GB9rpJyB9TQ5OX0a4WV98JxoLgoLMHMN0ZLlL26u8nxlDxZzFI/PuWH66//F0iZRu
h3vIYctZqlD7MNsPpWAt6aJ4Gr0VeOkoXXAEuViJZjKwcnsH7eJMGjVScmfEIn89Tfg36xUt0pOl
pb8ovKs1KFbfauVpxpqTD6U0MBYb4EmcuCO81dcIeAWqMhYxYPHEeZ3pH+Tz6ebDLjPFyDnIh5qN
htkqyPTgDu4uhzcllL58goHuMsXiBAfDn5xV1E+tT84ex8w9d9oqceOyktH+E45xupppIhZS4nzq
YgYfXFFsu27wo4OaqULRJNM3Uje/2rNQivF4FSeFPY81qs5PtOSQfXTJLBDYh+eghMWIOyi32IRm
JEbw8bxBqZtaxpAS5iXQo/y0QUKpsdHybjadUIZ/SJKX0C6x3JJf9a5OQHs2PheeZsyOOIOkmCIH
2HxBpK99h3xk+wI+D4Zz2J9aDHHE0ZjrXDoKIIqb/OvFRYN2QALktmHn3RCuOwJNCmgp8URNa2Zm
DXNHKiOqClWghdks2Ebd/sddzqHv0be7RN/HDxkWTjmMW+hsXrgaRF/6htqVSVgJ3JRMuivPT4Jc
a6Gt9U8G0ZwqDYmMmPS4HX26o1c9wUrk8aznSx+gC+GHkOPQHEO8paZ0iErT3b3nZcJ97sJfoj+J
W9WZ8SJ6KITqVB2ITjDTD4UuW/nn4B8us2WjW/LOho2At6/cl0oKVGNPela51WQPUEk1jcPT/q+g
hxTuCpF9ovIYDRxf1Ws1x63l1XL9cKp74D2EX78nUm11AiC7f5dDSXt3YwW+b2VFTgNMLmywGNJi
tmb3szeWIdZ0OWzcO9rH3krcfUwLyfd33xMNQsord+UHWhDzS686UUb1bGAgX7FSNbtxaby/4vd7
CI85htymqBTbxEPPshg3HbK06D1VSJPAbGKZ20oLOsOylRIgpGRRseQzrDldgrwiA4/zd4dErpt8
dgM0p6kOk2suher7Ph9/DGBXv31CxaiKIBSPsexMLZchbrMUlzSLvzSnnd35JUg51FeLhua8tMRl
lKBV8v+1wNYCgw9b6U3p4HEzjipwH3wLnwOxMfDwHLhHHMNm1WX+fqwSMcoQnvLl0yd4ldAesYdw
oaFROVDKz1PPpdVchVbjenHyl1mZA9HlxkvwtdWW6NCzNeS/+/ofW7OWifSlF06nJ4VLRJCRw26h
NWE3hobmFm3IcKnUJN7E9K9bPEH9Jra9yxJ9rtUhtcBoocr3kohJlfmjpm74tHXrXy9B/EWgrD8v
Hl6Y44KU9CtZNpr1JrFSDzQrbld8XGfHvxVpSUC5zl4b4gz+fquB/g2N+pMQBBU/uGRnttQbTw9S
n7IGZjGnSSV3XArSpnyMC43SiLpeMa+o0A8zujPl7GjgnQDTIakg2zUB7BFdSyQGDFpwkXiYCDGo
DKvO8MlOKe6G4u7cwMa8XmmKZ5pN3CP5TIpGjZ2+DQXM4ARXs1p3zi77xLd35uJwdN8twe7lenhR
33jD0Ozb0Wk25PIXGZlLE5y8ht71QPxP9ElnPiE7BVUC3QUPHT7z9ADF7R8K1yy5u/yJiXcO002E
9+KPINba56DUZAp9Dbgwp7ArUXs4ELAMRCyoZxGTkko/gdkJGyGcyfx5+Ya5369rj3TkRXhZV3G3
LQi30N0iUkU2z0tp0Va5lPPpR7jJOy0SdBfAIjeiEJ5z1nweUh9AAV4VJM8adazL4KuV7+AKfe8e
r9GeyAXtq4xy/dT0IpbGCBu7zp/2pDy7430i61tdOCYAnxmF3eg+LcEiw6EpYX0+hOWb5Yts1XFc
xEdj7AhTCq04VHhqujJi1w5d6w7n1KsvjJuSGL/KqfoMFgept2TDBF894k60OlYKifOE/jE7hpAl
ZQgLyXra7Bd5MicRtRR9ucHod90LLl16YUKDD1KR0dLAb59hy/VPI7jziInk/WBDIFFxDvPxA+ST
zDRi1/nZaWVJLSEv5F0L9GLmhvBtJqguLpKGijoUhX81qE+zbBzDgwljEImjF9cneYpcu2PrNAzJ
DmBHX+oFIs9iK7chJIDhj9pZE6BulACDowzpyzdaSUPv6WwhLchMG8X+92Uc4wH6oBJ/V1mmkd9k
SaWGRPFxeI1mqHYuIA+PizpQnRfm1HggA+fBhWxSGLDk3ISTyBlua5Voi8QOYjyN/s9EcTna5Md6
x7JZkNyYoZIgRy9hYbBmesmXrgtqBXn8EoEAGY6YGFFi2/oAWXS08/4N46Ei+abrshfmAchVzPOG
8MH9I+KTnO1bkx29LanS4WOpOMVUwkJ0ZhYDemkfDcW9MOoDBvNwNSNHQjYYOl6AupJzqr9LDYmn
8IPa7IFStP6IYL3Eztlv1PU9Sr3AVk+8sK/mxJcud26t/5TOClOj6ECYCK14M8q/z1XI1Syi9IW9
6uExD9pGZd5CR/MwCmakTa2Z5wDNWFWQpU6sL6P9njA5zP0tctVXq5s+3vQyQMc/FAMUZQZwWufF
xUoXWNaRkmzPCptvHgszy/TvJQf0chcVywK+PxfiAEZG0cOnDfzv9D53ADWSAHJyA45/qlsnpK+k
DjwfkRyH/G10fsLDGs69okpj25idS4li3QFRqmQkxnBp+oAYtqlGAczj6JHdwSRVsaiOf3S5Lc9n
bv263jcC90Bju8ENcy5ThLv+uhTZB+C0khWcvjx6yQbcfQHA1Hg10q5VcPImIwqX9H4ymTzg42PL
XcRgMqwBfxgP7Af5TZtdWI74OV5enEkUUxMUZmiFVgq8mMdbJtvIL1nb0/XnJsOEByhSuEkX8DTz
gNGI3g1gKyFxqWxmYcc6iTJzNT61f7CpZNuZLjaybEbquoZJuarA+NTO9mrFMXm+ybDa6NZ92LEx
1NIsC9KwpNVDipaCald9VzASKu5JHpOqBd4PRGIDYqSxD5pQcHYmz8ACXBOJXmQir6pI5Z+mQ8Rt
hnS6XzmryIY7lZYmx/Hlh6XdDW593gMEaAg497jGM7p068rsYipGtryrUzzQkNsTaLWK45I4QiRz
kp64V4ZF5Wa5Gx7GM8x//aOqjNwQIga9rWGWZH9zw4eyLEOJlqJSjY++7O0MXOQuRd1EJVpi427f
I1SKg97gSPUXLX4FHWIwMy0FV3aT7SidPGJOCjiHRUkP85OjMhVIe5NBEAQ/nkptz5dQ9vPvUEdE
gAP545YsGaf6Sc80fPyS8yJMZtFRQZ0b486IT1VQGDiHa4tdWSPPZQ7XI1MNQaUE2SV7y5TAJfuj
r1JX8zlA7HaZRoYczauyWODN4Wd+ltKsHz3KZYgCboSUzhz8CbHaIGna9C5/qMCY2A1746VY8WPo
Pqj0Xikbmmx/ekY75E8dOD7//6xusjLKyuWDnOQwAWm1LSnStFpSzmf5iZu+/VnANruS4Dg+WRJR
c+XcRVHdQvtJtE5NqZXVXFmAhAUPu4HPcET2cl1UHAl4NvffAeqqkAKZ2wVQphuQ+eOBpJJiSw2r
CcwUQA6xUhp8Hk2Uk3HAhCarUMRNLQS7mCO5/IlmZlKuOlfTMAXM6qnpO46O5ZvhT63EtnZsyQWJ
69q+Qv0artoXwdGXPW+WA0wr1hOmgVXjY9h3vAMiP/c0aifJS3icfLoHZs+YMkXmn+s9n7Gc3CoN
SEbJXXE7GzpUW+YfWcdg3E+NKwNwqfi146BPX7DxiQSz7ml7rBFcRzc7ELrZFsdvBA/VCHY0147E
aTNj0shR6pmcLidC8zuFDbWYHb13tKa3uQemEbghLLDHN+8uDZNZPYBx+Yjd/036BwaIp7KfkiKd
FWNu0CQhKDykJ0yIPljzb/72AI2Pa/3uOE6xnvJ89Rg7M77LcCTVqGlLaN4uh62VWHytVM9ZaUZQ
yL2YMK/9UUXyH4LLwu+0hqpc+W8Oc0Vk/gJ0KC7273b+THc7Ns4sfFKlmyRc8+Xd3c6jOyyXRCOC
IzIxvEsIPF63945ZrRvUOQUc/PtAlL0qPUeo9yu3CkrEVrRDwKN2lwWfbtl/7Nf+4+T/vA73Eq1B
SNsdq//QxN0WS+QhzC3ykbzkudJllQu+HnNiPup/1vcF22LD9qud+afsLIjNuC38wWlzjE2Hsfuw
QNE0a+uPsz/qQsYI6Bms7G8g5GjHojJYHUpcO05Sjyj0uh2sw7MSXLB3Hf8GuODG0LGMa9HuURMU
Qtwx9L30B2dm57Q6x1vnGkW374qw9KKW5nXeQDBypmtRfhLB2+k46HrpeLlBPuSr9KgsV7/f/o8d
GE8mgSno+qfnvVHe7dk8dnOXfvG9xKgK3NFtjeB0XtDER37S2mrM5Og+nnF/8pIw6RpzlBkxTR6Q
irTmiXfoTV4XGl+oEHrPTGdj6pOoBPDGOhDms6nXTFxbycGIf75jqSP1HZdewWhF0qIdBFjvPo9h
utOW8n4xpnuGAAiRFmmTiZyjnG0Si/Jj8L9wbsCIHvt00CF72JxghtXfPZG/yFLFhOgVbrWeKArg
z4keKDd2cH1lMSR3EQV74iMfJSIepJTxaDJ+jselxYX4/GkLgQLGsuaAMfQTdtN6BFxilS43xI/S
FM9QD141fJ8QeBuwaZ/UrqtV3tYhbQd3vSNIFGboxKsOrfrDDGm5dFYlj+cM0q83fQpSYT3VMXcl
Ze686mHl6PIsl4ccScjR+JYljvPtQXg++1qC2Reb3mzxo3dz2IkdQm3vhEyYKJ2vPPF7j4MQkbq6
KeHJ7nhY5j4HRTKkxhR7NHITSHwMlnnyzyNZouoieAcn6woRMy5EYcmJoKNqVZTNtqEB0FIkb99z
69QwLpE97xdgSC262hKoxCcCRPYOurK/eGSCZ3iucS6lY5KL4MW77qW75S68ULXvsmMEhzRMHc4n
zDIcFNTzvKdNhgJtevtYY62xiT89boyhhj5lnqjHkcPoSc10LEb5Vp/+VAXMCosAC7XMsgkF1oBi
L4+cfVJfheR+zN4VhzWYKjX3zpy9buawZun2RJAjwHJn28DKmoMS3DH7B4vAKzV9SB7CGJpJxqCy
J6RcR4HVt4sIynXSJXLds15ED0cl2oQwuF2jxwWm0JXrkksWYIhWCExu2fIlu/2TDR5T7nCJNSuK
Qb9Tj4W3oCQZQbRpRfc02RBsbH7uhFIktYyGk2add5sLNP6Xnf9oUaZY4O7dy2+qMro3w3vyi8UJ
y/curoDYomDGoyKysywWN/KoOIkkwLIAXR4BKBuSmaCUy8+mmjrZeWZo+/nyMV9jz+PxgUNCjiLX
iBQl+m5bcScrp574tQf+rjzeHjEM/b+JpfMOOqu5q9dYkcI7sPFUDse6KelHlsR51h1umDoBuNTd
dwj9z21rlQV8jmfQ6KuH6IgVX3qlQXTI0+x+xmXws1BEc/FV4isDhI4PywONp4CBNaK+p8qBQhS6
qrcC3uzrzGpKbAdgAHr7sjR+5+6JQEfFT5Qb+K+WgXyCn0ESdxih0ugPfe0w3pyFAnYfDVj0wBg+
4O9B6PSqOWVQ3PFzBUFVx+tIoxDL3jkxmzxkF8W3UOG2RW8woVz3c2ImvoHFrlfbcQvGN9prLKn7
mN6O8UBxlA31uoTX6Qxeaf80jC0ZfZaxbv06ZHjM1hPrUNhx7cc6gft2zxDUy0k8DbGDzwEGBjQd
97ivYwRHYUmnGXHIVg7bIAOWe7eBO7QfWdIWInNDkHNYQcJ8JIPEl9aCPEexiaeK1JBlJLKutj1O
usbOw6szfrv6Yvh9MeIvmjP6vQesFbNfH/M61YINWoOSrmGQWU8s5Je3RtX4DE7w8QSQ2Ei6KiHj
QIIZfYVHkhPv/oGWdLUYM8X6gFCTMLROKDQmQlXUdRrwxFeu9RGbB0N7o3MlTeFjkfpgvKc1Ckzz
zKRvC48FZuQKqH7S6yExGxyhDW5xrQUJUEX806tqVohKNHXQKL6M2rcm89oU0WpcN8E/piTa0qfn
HsttAHQ15UxesLJr5KB6g9MDSJH7MP61e4eOod2JS6HlviFom8QYWPVj1tv1mx8Yz1No3P7O7jgn
ymkbZV/NGSB9KTeG+8fjTnof/r9idAZo7wuaNs2ARZpat5zoQBKfh4fzhk4RERbfTNxm7M5bM0bS
wINIkbdEIftVsAcGvtDtCHsibCOhDJFkOUmrJNH+AXjqaev6usmUVlsA5vyRvQ1MPIgk+V14ViyW
pXn4RNuihCH7+e/C4qH4p1GxSItZ5d+l+vqxeEjGHMUQXtstKycE5Kr4RtkF2vaBLDlhTgmavTdI
b3Vb8HUaBqWr+ezkhngR+yhNrXu5FAcaqeRQ4DX7Q8SK2lFWiiVPjpiwvvAWPvV7+HH3gj/dkW4x
UrBTFXHsR0IpPy/wD4r6yPw8B+2V8k9czm0JkG+yQ9+Mp2gnzzjBV2IKDe49B/41FvCvngD+D4ng
947uLVHXYNh3X958vOdAcWubPBfcrFnKgJxk31LUgkFZN7ykmfmrTrej8FHrZtScnWNYRBzYihKu
2CZZXoS+vORFfXzi/imJ9Sr5j4BDYVuy84+Sf4TEGLQGOb3hS7DuGOEp7pcWc/FSnzY9apgsQLMJ
6ExxH0O5IOsSIP+HGFTpNhxVLT9M1zX7GvTzguOeNGSpTsr+Bx8ZeMKHQTZ5/Sje4Pn9SOkJFbyP
fku6yOGxUjqGWooSut5css/6ODwjbRDSj/nZRwIGVVQr87YMvpLyxTKEu/0+h2pNb6Zzh8IPG8SY
VudPDfcVhGTSlmCVwpsCz2RQhLssrqK6zvIIrk+lGcPvOUjQU9fZMK8PlkW9RUruGALy0dgW3606
Hv69yE3ud5V7IZPLOttQs0qWifreEras+I/7B8JBdPrAP/SIKMFarn8Bo0UnctQIAHs6LJcrboy7
/f6nThsS2b24ACxILyoC+tXeTD/dWSUyDF3+iLEqkynDk+9ZAPr4DcUUTlN0XE2EOQkXtn8aQJhf
Bv4i9Nmg3wYXqzvwNTtBV2hyN/WVpLu+gnxMufEM1YAf4uHKMZ/R9VO6gXumubHW8K5r+MI2kR5T
nKMIsp78a9CLz/jSSZNwD1UkoKzXy+Te13DPKbeJVycxHDXdsj0D29fWk4OTjRe7V972hckViy1a
H6J7zWzxWvNSEsa3oLYMt6LyrPhaf5eo+l9j7AmyOz4ieHfwbbVYB/3yD20b8lZoabLZrSDh61IU
f6pJ45xNU/eFlXO79zwz9A5H/UrgN/RYGtdATnClPiuUP045tT3Hp86/fLLjGNvEPIifFOjiCBnF
+bDSQCIfRYYXErbgYPPnseQYV2OUbNn9HvCEKdVP1wANnPSUMXB7Guj2Ft8amNoAWm2SrDJxsftX
ujp2G52EGd9VeEqErGtBKIH/hTVH/d3wGWJlkSp5HGQFslN0glEhbQ/Q6BhvXqe+vUlC4nJNtJ0E
JN1Q2oBQ+c0eFEzyS+pdnERQ2PrHl7ugP5U+SSr3FXW5ywekGqy++Uxq4+PVZ43bXc3mZL7CYapm
RYYkm7/YvrxpK2zwrlZNAZTDE10V+P3Fpd2pVKDU3sSDRPTZJ0EsNtUMOZ9LZuexiDKvXIRlV53V
HU+eIb/lll19j1J7g8mWVjO5CECZWQThhSvvcGpRXEWM+T8vEj+344+9hFPJhfvnTSskbJaT8SXC
NKod185EIQSXitZ+aRC5hD+T6S9lR0tIwPFjxyat18mWUHEW553IWOW0HFImrB3GQdbkR0yBJTXK
F6Hq/UN23gQx3gQU9yhFojCvwpWDaNcY3mnhZTP4lFF0m1rr/pPdCpAciiX50OlGFnK3y5QKMNs1
LD/Q8YvZwrWb1dYTNpj3KM7gmD9jyKpsdukUb6VPqWaDSePyxZPVinrQwCpgq8OsjAambLoVOKj1
xIJpbvY3gHGsMQp8es1kBlmKbD3dDSuOfMpVnNS+mCGIgMVFdXCubdqZhJIZn0LAhqW4Ka/SwPJA
XN6PDs4j5WEWs1aPCEElq8dM8pQZ7wZUVP5bX5uZfqb0tQfRGvA0+GMDu830/frAuvyNkI29jQUN
flCtzMNEtIhRWXMedozeKMTcOfluD7rdBB0DCPO3Pd2SCcxKN5qdTAHioCzpizhC47tRBxVmMLcW
e7y1qMPcnXOTYK9Ps9WskJtAjuty3OKe0Vo5o/NbFCtFEioMg7Y+gqEcUQUxave1ZUpNXffkpdih
GLQwCxQRByISh/1d0/CIPR/65KiOj3L0ggjAZEjaqDplxL1POkE24T/XOApGvXGE0Eo6NWgkXF25
D8nfuiaO+cdv37+T4g3z++yekGr2FgpdMa1OUdIBEeyxBDteFA0M2W176kNwe07Eqv13CLFL6Ft+
atsobU6pz2SVjRNTHr9wxYROIT0lbYVhlVX6Ul99UqFin1b8vTgpN9HeKM9lgNcTYiVWMOZQSopF
eokc7bRESiEnBLqJqUAYBHXQddzl7gsJg5DDYggL9f5zKq8fJ6iKZScAGYV9Wah33Qv9KnBPV8nM
natV5I8/s3UQvFtORWmNEka6tR/R9yGcJ8F3VvgF8CsErxo0iUC2/Paxlzq0PK82LiPOAYomtNGr
dnBXmxESLlTTnb9gUGZOp+rHioJa3IPC86FmlzoO/4eCUSamdyOzPbNA4gE6nHoBp+59eROyOskR
kJm+c77AtPX/cSigQOEh4DyNgx+MbhJMqL7Ex2bPwCqZYgq1JoLk/ofWxtsf1S3E+4aWXI9zmkNb
gULzfjiu1nNzSkqH4bybW6snR1vQWr/RWuS85nFZM8SZmmSqaP/o93lO5QDjgppI5au5KwMIOX/r
Mg5kMI14vRYvr7oqniMek1b6GmOhVMMjKTyzJcB2tT7F6HLp51RD0Xd1Ue1l8TlZ3PtVjbRBV69h
oQ5MbyqRBh3p/5KHkE4sAFxsNGVVPdpZr/elOG3opX6pbHSat3B3v5HpZa9wiTJT1Dm1SmtodmIf
R8Ee8R4Zd71+G17zs62pMQoC1oSR6TMNLyE56HqI0m0t+Zx2a0Cv/SEXBrgE9U/ooHZ4OzmLqO3/
/vDbYqtigX24s5wfpg2xEXrIWX3er5j0L2PcomgUX6U2VL0h0ds7RzKvKKCvjGUcaH5jMa8zeo7f
j+ess0k4pODFHzudiXN5mJ2d0RyYNcFPwFESNxM8PO2rMEmBZd158NW9kCsFW91g6u1VkiojIiZ7
W0eRWZDWPyd5QxCdkZm6bJbuXlCZluf0XqC9haobohV8CpPWiT4HJbnB6qja9Swxl8KvFUABC96t
QWcTxVH5ZsBFe/jSWQOxS89pOCK2SmITRQCtZDUIo6QaKX8XE/Kt/h/ZsmJLs1/gemOXTd5jkbua
+nzWO1TL02l2vKCgtlar+QuWTEVh/6ZkS2Frt48MKrQWA/01Tah7hOwdv8gUL3mjb83m74gffCy3
pA8ioBBmhPdGmgdO40NfTzNOugldnXMpecci2K/h2c94VKMO7nFq3cIBzxZgorlfxYEjc94EKDb5
tJGE5SKf9apCqL3OAILM+bEDtF+ZurwBzdVnPzyVpL6VPGQl76CYsiXgeQDlpOGElnphYTLbDCLP
pURGUeSLsiv+MPgzLyoflSrsTL8Eoa8oNTNxSJmFVxwKKgRyk4NYAI9w6Wf0gc6fTMMePmOVxras
1+LuJeH6q8VwqMRZUbM9hDGADuRmaA5bXn+EwdLhFznnadJvJ3Hnw/kWX2Urz2+siRq5E9f3NKDD
izpU7He7o8ueZnPIqwqxZ5Uxd8Icvcktfo3FdzBE1YHR6jsPGlQk1P7VKwa7izOldFzqg++KV3sp
0r3tmLlR4vjXPP7Kz5+v2XD9DGVc5CxI3AGT8SI/LeI+EO/7aXVR1m9BWPgLXUzmIFXXMd8t39Qb
9MRRO/f6qsX0GRXqr1j3gpB5Ksujl3haNH9/0gkinVDpXz9kVp9q/yJZM40sJ2X1h/ZFiFUI+Nbd
3E23n9Q04i+dNShKGg+m5nWR0D6W0DhC/CoUsGcFxdpK1vp5OpvTcAozFHIVpcSi4Pxt+fvh63uC
DVsKbuHm+x7rMfUEenKax1xh668nEgqIctR1M6U4x9Cj9YrJ9C9L8wZ6he6f9mV79UlxspsmEtr2
hRxugVwSuilsYsdYfuSAK9FLFa5a5JQqIfP+M4wRy46QU9ojadHTKMFVWcW0z+3bluUZ0qevehdU
7oZLmfMhPkCmOZqVGldzg9bVBrWTXHzp9n8vt6437Pe2mR0cFXBfq4nop6cKrMx4QHaRimHJKR4+
D4Uax1OWV4HC+28VQAEgRVDT6lSxrZCc6Q1wqWOP/hhXxTgzGSFrRpfO1imKpufElylLokqqZ1xk
nKlIk4mAp1OWLbxY8zdUY+cUa8CrnxJN692A+DXVI0yU3j2BjyBIXzM216UtTmUYm91p3pSIhlzM
dX0XnWWlWD35HmlXFNiNSD2KEKwfuA/yFNTA4cDlT6CzvEa6MKWSDy1INPRe10OGntCvy1OCSK0y
Xyn3nwbAJc3XzapkRGUphj89DgztnMZADLQzBbpqK1SOGcDg3KPCXUubZXmkd6Vizt5jQgctb9SD
UZxb3E14gH+5+lXtDUihlufFzzvFyIgeFdRqyijwCqFM/LO+sBmSwbpw0605sF+iFG6wGNSzP8ur
49zo8Eg9q0TnZxTsliz2lDMzd9etCPIverY/qqK2gcBU/yrM9NYuGr5SKa59kfm/WvW56o52yrHf
yPpbGZhc6dRXjktLW0ffOUzwCysQbDLJU/4qUivQ1o1EIpRZH50Q8v8xaIH9pPgm6T8fNXjBzqGI
LdWJ2x5CsMkLZHu0YoWkaGKfzpF57yHWYMRWNdbKsTRrPDhMvDRlvKOatykiqpMEV7rQZHWCIhcd
gPQZA0Pl6jnWpdBS8wljfN5YWRCt36caKJK3Gt/pd1npg1BMXayp/3JLOuM7XlCAReYRNUO8amM0
vH21Azzvf+azUwnouRz+/xgzGy3il6LjHbsyDiaLk0RFlMZ4/gHm7mUD6rAn6nxM/8ZH2ILP4ON+
q/I27Nmxyrwv2TBSGXQS7wkNuCtYulqcypt9PdbYd7VlpP/ugrlhqIBBHm9EWWsrI55umLRALj/4
/kEHqEkdCyICxzL55d24cqnotTehOd1H6gWnxxGUx9AYbPb1b0UCCc9DpCXArMl8KZShUrMeVPJj
Q9bQRDME3roMIYPk7ttWKkcoXeelw/YqEND9+Y93KGTdrTKy9TsJmdwYjIJLaCH+BCodhZMwhpqf
kRp4Rq8vzE2aZq0EzOSB0h/4VsVXELEe/2gUPVnbDP1tOL88ZNZNrUz/3gnQJtv13VLK5hHANOck
IcPhx5IZeTZZUBqnRQGXrG0no8CUOurnV6fXx1G2PKKVyyz1MARicMgyoc2vpM/KEMvfsmfvh1xD
irQlwL0fSGvoYGfEEXygl6Hl2D7n3PHRFyev/ZWr/KK9RJ2CXHqTIz57AtLpQeNA474uvzMRyn1X
xmF5/o/FlMYwqFjSowopb6dV2IVmV7c9r0hTdRd3QTIxR0Q06sB8TBIcvTs1c4XL/INhFs75dE7e
Tc6Rr8E0y+B87BvnbPl27pLklWo+WzYEI+0Qnzge+zrSpy1Dv+W8A9BETlj9fyqsUYrD5WjPzUEr
Hn3IyXMUfU6hDnAOw3dRWBOPgWZVJY3OwiZuCFvZbD94fPjAwdsgjCi6ifLUF52CzH5I8//XGtH/
fccbWUBuTxCXQDvE2ScQ0Du8GTK1bnP0oGWeiYAJMRs6gfaLcPOuhPFNt9gUkRklP/XanqSAsvXv
zojj2o+7+7eNmSCd8E1pyHxQc4eyY5gZn9Yi8aMoJlMiDGBjFKBFzqRx1M13b7GMwtPTZns9Qg3E
AUlqLLAmZgLo13lbZ4K5S7oLqYgV4nINIr6mEmtmSk6lgLXhQardPGChAd1sGS4JjYYAKED6L23p
zmrl4dTvrveEjiBYc3BA+rpowkgzAW1z7evsFSc3c0inZDIC0gv5RTcayET+AtnpY5/WHOwp0N4I
isvIemG3tO6pgbFkfyk/UiQ1MXCYrMo1QGvyP58jOEv1/QxOy8niRTSvtxEh/9JGTqh5Kwbxub/B
ziK1rQrqu1VZkKxjBmZo/NZfKDG+BE4KyzBgUIwCd8zByarQGuwcX3zGm+QlJU5Oc2g6RdLoo5X0
Rn2BvAnVuPgnSdjb+jE9f+qoQVaylIeJxFuQW5U5JOdWm5L6Ng4H1xM3TCPdyI70pzIfLG7HEzhJ
paZEGMq3O8Yb6GAY5V2ncva0qNAuhvTi5Yfc435rJqFf3J5PgtbyzODRkzorc8LijwYLPmYaB4v7
9ZTKN3Dd+AUG/Qlpgt9vAMY+pEBHeGvUDYXR6AGqjKpkAMn+VjNzVKjbQTFerroqkoXrgoaCkOgf
CQzgzXdHVCbjin/9l0HJi/ed8XgJK8xHaW/LzZS6dgBnbbtViWF+Ny/tAZ3bZ1Ecd08vJkSruwTy
t9nsnbu//arTYrU9xAWM86OfGEKb4i7ori5B93FwSE+K3t2w33f2p6cMW5XayTvr8hk5uR7+QW4x
eqRtDDpDBjgtUiOdjjGWfI81ri9Z5r61IxKSRj79scaAJuO+YqmMdRWcUHfME3OofZY1W8r/wfda
gIi6BqLMbM8bYtVhUM0iJjSU5xrmvuw/aQQueL+EIvz0sTuERcgnwmdsnhrrvtya0ciKNSefxzIl
cnFJskBN+2jXk8PQXsLLZvW5/iLwrRDoS6VX+h67Wn8FIRvqC4xZ5E+9MFLN/HHl9vz/AcXOcHQ4
cTw5xqT2Hhvlndf8UPv3mHJyOhYqPdk3XWAoUlN5osmMSJm507SSqezsEV9JNv1tQTBWrsYbNeQC
ALQ+sTtewjgGSB08VDby3VOJMhUfg8mgRViQvPLmofmiNEiklBihx0wQ28dfzBknpkpKBMKxeSAr
fwSdnKQ6Yd+HYDJup/JDpOgCPlY6tGUqt5HpGWe3wC6d0i49x3ewTOkvmdum/9Z6zrB9yNnuEEpv
Oup1DS0fwIOzaG9RHMzvx5uhzYuPd2kxrHEkHwWEaw7n+YvwKsCuMmAVXosjofbuEjvetZxPr5KR
h/xdZ7JBu31elQzh4lzpNKg7psKQ541s6v/Cwt5WUzDx1HpFE8bccYT3Iyj6MLfedW93Pi189+Ij
ZUnVNtL6MVE6LdeI/e7McyYX5JL1EHLGg0miWQDoibkaablMtOLS8rZAkbXBpShVqMfRhV7ieoLr
OCy1wipApBZUd3Wjlp9e88fnh5FKDXCsR8jazHM0/PtgQFrxQUOw9RbsIT5ZTbkUljYFGnJUJfVB
FWbWQevgqY7DJhW7EtmbXH3vdiIuaQG08Gq0H5lJqr8+sOh0Qlm8aXQLhjBHOVYvaVVzlg5vJC5S
fmNyDdmT3lcUVOWNLTKxUEb8BaVoab2Bpe1QjegaMLIBsTtE5GygwZubiIHk/VwMAyzWaPFt6rj7
v20H4V4unxB5p25fjTfZQRTp407ZfQzBTr3w8EpIUVFK52/hU1y8/4TRJEh5uqrW29WxYA0bs9KZ
OrJ8qETwtj+RHBy8piS/KtLOwCVxGYCV+yyX3/9qAV5Wj1STdxTGpPI09Fj5OIOMuXf8shwa0djf
MtyLXCA0ypQGfdJQSvJTfsquZS2K4hp8XjL0I9ToGPR2vod+dLPUFv36JaxHgZl6mQWJIkXSijZl
9TXVBFXwG8ZQvk8ZWE7YO4ut0HNCRLJcWLBKuQ4a3t0kSFrFvzHcuhW1CPZZLmIUR4PAD7l6N3f0
FXDUPAvC4r1QOAkkdz452t4xTkFm7alwnqb0asQkjMCcEhZl2P/oFlvxEPxaCATuIGt1/TomBq2b
I9YdB49G+FZZ9LTD3J3fbP/0+Z95EGPvcxjzX5CblnnkFSDY5njSiO6yIHzghbHm46cWqzKXsYW2
9AyiwaeTnCy5iPZHcIRZsz1EWr67dtG/Ujzdi/uYmwlW6DGsHo4m6mwEdQ3WvnUqBPQTRYJ6aukA
kuBIwZawZjSJRQfDaMMAfqRa+FWu3jGrjdz7asztyydFLX3bka96pnxOPxwz7FtlZUox+2/LyCq3
229AX5hfKmMjkSeMID8SwuD1HftpwUbGiv/5ib31Wu9XioGX+xkpOOvUD0c0Jtqy+3kNVJNjYDgI
uL45AHhsNDcuUVOK6vXR1nHPDzdImyR572ZhPG8uLL97ybVk+ZGa1nkKk8BCRbFh50zo6ALwH2yg
6v5oBH1WfxzL83NhT9lZlTz+a+OKfNak9pa+c/7jFNHwbTNTryw+Y4DQT347KyaBDmUmf5fDKaf2
4D0p8Wzo8uTpEpRUyEepYCLSN5nijFKOXB27MYp+vyEumw6plDdSRD6jtuf5CII/+9il9dRc9Lc9
wDbut2LH2UrRdRWdxhL10xnGj0ZcOlL8kmjOkjsVuKkfWs95cxbhPVFK5ltreTHfyhYDtHD6jZyA
AY+3p+/T3aLPf3hS97YPVUzjAmdr14hXwj8O9XZmV/VwY0Fmx9ZK0Bo7vX+bPJjaSKaYC+/mdoWm
8E+XEy7a7JWCwJjAauwx8xeFLB1Jwrn4LBySRG18x37C68y1jWzTwPiSPSiXfedO8TzMB7CkbuPx
6jgldfeP/seAi1A8GhyHyFAthin0TDHtB2ZS2wfbxNdG6oKU8KzbdHvEzg8Y73DMB6FsF0Ksr+7m
0Kw/ar3iOdns96JuCmTI/7JfwBSwW4f6UqDtDzhO6MPx4TkN+FyprDSGqSwWXKBMrdnz9vFxDIQG
YoP/wOAM61Olz4sohOGfe7G3/kqJ1CWB7T/qdXUtwrRei0KZMzC3CTJ2pQevhgEIHuhh9uOV5Us7
nZy0diQHiyfQiomaVbenWsz/9YicveBbgwIRUbZ36gqO7OL2J1MbYrsDbCTIzCQbsXSbJBI9SDTd
v6+LKBhwzH7+fCF/aCEKZgYxkDvOZ6vG0XtqcfpooVesvtaG14XUktBFs+L90y6vDq7nyI0xAML6
jy43wk3xfn0tpe38rv5Z1UGR5cvIw/7G2CmtBWFh+Cx1HWeffwXH60jG5o7kbhKt1pnlLFyraWVF
40tN+3sRNgDg+3vMjdEQgdCICxappt0liBGtjWuwPThP6eqqzmsWcTLBJ3YznYb3NgSWsF9RHcaK
Z+XUENX8ufQM+3xV0loFbzC3w6gB8j8thges76nLIxUGNTsuzP4NhI/7k4JzbHgI1dX8ZZuPLYPR
Rfn+vPYxXYP4sSIeTAnaoiHv4LkcOF1ObQXb8vzWj/tP3+wwF/iSwavCXNLJQ4b8RXFCOnK/6/Dv
mzlKtnjDjMADwHsPdlkgKWu1N89Ac5/602oKgBVHqE0/8ye4hlyTmneb+/69MUonQk08wkSnyFji
e/49GSp3HOdH9r742zJFcD7w0KLtj/G2BlTpAAZBYV3I+OzHhBATHU6lIjtUbeHmvzSffM80Mzzl
PamTpNrxHXjxqOoxUpkWGKGrPk08XsJEbqo7db/f0BbM/H3+nuP4qo+4ato3WMeVBc+GlIegQFhL
3wZPDdUgYbMbD9XgLmOzcvQd6j3YN5uCifIRyjaQKEZLwb9cMTghdEKS1fL5CIJ6NCp+1UsXXQb9
C4zN/WnW+tFfysUcsco1IpaMi0LbxMEqUCOmwoDp2eytLDTQbR40c3jmU2PRnheCLfz0QKaVTgBe
MyD/safwfiTqWEvljqaoVnPPmtrdtBPrTWiTB7tNCVl8ZIDihTthQC4KgPSP7NuKEslze1khRQDr
Wc7WawKNxo7rCyjhmAJ4bCsv6jtw7a5NXVuT6cTrT6xonsO7/J4JixMe5QqeKmM1b4spZndpfPfn
5rSKVQptCgGnedCqzQuEc8RMQFJfntyLIgQ/YUDfa+uxvaM3eOHIst7aOoOhv9WzkwAdrwH8W8Ls
Fa27Tsy0cpt+7Q0bmMxrKcxw62/YLcnWNhoVEF9iAYxrhGRnHnOdq2UN5AtwKNlL29E3A2TKUbYj
RhsrQ+QGAJS9DZa76I2GjLCRUGgOSXR11hMraILXM57sBONKZfiOFhGAujaUz3N3TMcYc5YE7rKw
HvgDo2kbj4Kcqz8XXM4KSRfhTF4NBeV9hzaKnSmadm2TqHXURXWrG0saFxDq4f+JY5d2SaC9CXcA
MU/MjX/eitQEt7ilRIa/NQkOHE5DVyrvKzgq/UzQ2BezSS0mdnSb10A1XvGlW1UeG52ixSm6juDw
yUQSNtCpdXXBZlhMoObTTL1NO74mmoctt8ki5WmxSmbeRER/iaG3LmJSpHNbmV0+P7pth1oo2dX8
afw5d+j8s2s0c+vbnL/TZ6f7q8p8aIo2YPgD+bQ4V9FKQlWfylsxkVOFfP6CzTrJT+quPVVSUMj9
4iShUB+qpK1zOcXjb59S/syfawhz2e0vO7AKUuxzYjV+RHwVfHAlm8Dou+7nYKJ/8e55pmVzP+ME
/bfljOaRQ2JC2UC5BFQJsxuPGRtc5fjIVaXsq9lUGMR3XQrts2MFg6rSHv33saasfqChp0N6ctoV
6hzuFWHWDm7WiMa62tPQ1f7JNaf9h19a+Z4+3POPeXwMsmEkGQ3JL9fN/QuWqUqQFBFRk6SYNFHr
LK5DDvqqZGklfpvJI0vvt5fhNBPrskPNsXyX6ZozDCFpj2Zd988PZUJ0fu3PQ21YBdkR7caQc4Pb
dysywwKu7QvO3ifZLhPQ34s0Ixx7A9SqyUHc8jORQhht+N6UhvpLXz57vwp0mFwa32aFHbbfS87e
PI57UMbVQkVy31GB6O6vPxjNxpWBNh721GhDwpq/e5XT/kFYgwS9dWBHVDMpdRhILXEzxerF8A37
77MH2ADabY7cEwLSXgKoIQcRGv0+rikR3iLyAULZ7Wf6Ej0YO7irJUdLxFFsbqhUrmLCQNU64hql
EbL6cdWTlYsWPZrFMlKnx7Clb5CpyZjL/0dbyRLVxgB+VGok8T7f1DkQvQ8vJguKTQHY6g2lxx6K
R3CWibMyZ3XMZwzOX9QwRDM+apks36xfmuGoZ/WdTza0k86Zl88V1VGzyrY2ENZjrwFkLz08wLUJ
3/KBeLU/X/4JJC+5tTB+KnJPGQ88uRiGcPsnG1bZnYQZ32DXzN3X4g++dXEgFBrttB2TfYL01KSi
mIoDHQ5vVfbCTFcUnyK4ItpFCKMBXPXN5RI0HhlBbRyXnQ/uIWBzlUe0FQvC8IbZUUFBTKOSMZYO
GbZXH1dzrQStH1uqfw9hjwaOfuD2xzU++AQTYlDix1pMPjg+Ns9S2lnCYFIwyAES/5Q0oC2HcuMz
6ABBhks+wQGCEYi1dKb3R/dW6pBHY2TqMTO/C/KUMcFMwg9c2Wq7FNSxn/JL7cjlOrvO/g7A/++g
INJhK3gLweliciXELFFGAuRbBWiSov5nVRBu5chxlLF+yzU5al0P2ERp0QgabLZYedtMUKsttfV7
xkUp8/wV+IXvN+qK+wNnTVIIEmKkGgCjxmGi0E4O/9QjVODMBC7F9QUm71MX1G4T4MjiXJA1yrL2
riZhCDmDMpKhk0OHADAuAnYkovTjDYRCX1bZ59+qXxHpx9qKNa+diglXssOpVA2HAcv8b7wqt1HK
+1m50UFBxLaxrWoNmPhBXhwTIndPEXVRP8kZetsr2UJ6ROgFdREzTfuFywuzvDOqjpoBehCIyaXK
/rKuth3bpytdENFEBAFGRnaY73k03+uAuZb+pkwZtZrNTaOn1+3JTXMYYLlh0qMZg3bRaAOh2rTk
a9GMBTkzm2vvNeT6MzcQNjgH2xvfCSBXjnhP57RKLD3QhKdRWhnVSP17xjx5pfN2dQzBx6mhOqzb
kFv6hzZhbmDse5n/9W4UkGuVXO0a/Hl5Vik3eg3t/B+LFiq+jnbQH2Gfe4rVOIotO+CDQy34Ja66
rIKFGFSv+aahAw3a2fh8Id8eDUhPcADPjswYcTUvjMzNt8hmJYRf/5Rz4vuFhGAvOVSH4NzldO36
mdybs+Rk50O7CaPVa0JUrp1lPQZtOemoxbdJRPdhSa2HEjuo1RxyKHLOkrpk58IHLLeMVjftdbfe
9MYXujdUDaIFGK3I2NJzU53DhOJt78qLxyU5uyguTa4EW5oMK71aPzBoSz6JKkTbCNJaGhjg8951
iQXdh9hrFzGGOPFeMfuX1rnzu9xuNzRmJRLOppYAUWHb/vxBRz4psyTRJ/jIPCBt4+VHYdxyr6g6
Vb3cDfMiyJuBfnY+u7xJCoPpMGrak3/ViR/hvoOFJn3vQpSAZ1CdLDYvk/g/WA3H16djBhcFvn1O
Q3cYZOJ5TLLjyYwfJCzqHX72PY7CvKwkOiztO3/ZudO20kV8fmzZd4jdfR0ilbZylMRWZtHVbsOK
h3wUz5wWrPS8JipFO3mg8nGW5ktH9Cr2qu7ws9klxggv8P2YjAEDl7SIZmwl0/GHEnf8BxFSC978
TQGvMDiiCF+W4Abztj5yl4tssWpXDziGj34qz9VqRianBNgbu5FC5xAbXeoxP05+hXltEW5/jLu1
68sUovkcKj2FUW+LCKXY94lPYuTm1746cAjoh/A2gIPwSGNOkyDAat49mHS2UI2yL8F2Ow/ezHWK
A3XGOMNAtqJmLdeorb4Yy+1aK/Tj4WavoBWBzJVS4B+0UruwuZlnYe+4hPaagd1DAloAPWGr4DUs
18pIxy75SWZSGxW28gpMIabAyoKwUr3JAsZ96L3IN4206ZaW1DhWYXMQvzzBiFiPnrQIsIfAd5uA
bMB+EaiM77d4JR30i1RoDUiISkcJqHLQJbOF9lkZoh5jDYmeM+zAJzr3649vWLbt/ZhD4NUPKlG9
Cb4VzHRUc57tCICNWEXU9B0qBXafpXaqJpVIsAaJvJd20lcQjhn0SVS3UqIvIvnvnytf5lD2JPwi
bFcBSlFwIc6Y9wDaAjSW93vfml1+CJV7ft02pl0Z6jVvulFlPelefZDD3gdZ0LlElMQWj2l4wKaO
QJ63C9N5BGboAb6ytQL7ujtH6pt4/kWmyStUBhtjyUnHpNZW7nVYk/YcOnmuHBqo31vzE98D0Uqv
o3PCy0pJA6cErObe0P5AHsH5k+PgUiHz5/jzyA1h7mo0h7iPQzumjMq1R/mUdjgH2fiMALbTo894
A6M4PmAsFkBrtVLJnu0If9RuFqTvYPS6rW75rgy3iXavdyRTyDHLL6qigUPw9kusEYD3f6bOu/oq
tWnm2HcQ3bWBTBzC7vR39Seyvrw3CbuTdCN6A8bkd0YDDPZkEkTZUJKlbT21gbLI5aQRF4gglqDp
pIzV7JKpygFL4R8pIvs36jObaPdIzQT+Wom9ihMAyftZo1wkrnf+snTL7Sv3qzuWTTdyzwih6C9k
RSQVDWXwMR7yHBlTbzaYeuuRMTAXRDgYi8YktSImK6wgnXJmJW9MsToKug7K5xgNyic/Z7V9iDg5
48dVJfu246wtSgpuOw1hkSfN25ety2XOPDtM2gAWbBRq0/ax+OrsOwhZxhzckbaInj/BmIGQU24x
FgTmU3TbBff2pXQKL9mzS51NJDn9xdnTCp7PxHty72l6LhdapRkpvFpIN587g1jnALMwHBMjOSaM
OYq1SCvxOnwdjF06SuG4+Dp3bebDtEpPMu0D36+J4StgQseeWl15BPOvfRgr7zjVeVP9Bq5k7AYc
Kt3Xikt0fIvsfPNhl0VBsL5WpWXCTpoFTGPQ+RWD63C2K8Z12w4GxbCArsb9sg1rabMge0FWthEe
TRISvmggz0SuGpy31Mo2Fe8ipVipE6HNZLf7UKgF73d7ojr7nugaVAtBBIwbGXRO80PYCI6rrO30
x9vNvYmBtKVeBc5HOrtCgVDO7++oI+xfGIgAdYG0uSuRs6PtxiwODyPmvTso+MxG1DQIye3/zqit
OdTpLocjNLXdS0pih1iDrJIlwP34TJlQ7HNwiKkvxIdZ16oOpPfj/Uuz4ZuR1uxtwL2xrWr7GHhk
YSxVdqaQkiBdoZ+7GOGOJejotk8oulIQi3UONxjK6CT8vjdg4ueLiMVRmFyM4jEXiL+SdlVBtjRk
/8jlafKvqIJN0UYgSUy4Wp3CXxPJABxYcYcaPrui4a2NVrv2kWNP+ao0OlPWMvAz3se2q2IyblYD
Yw4mcazTtTEmzoynWpkH9oYMHP6Na2hGntN3tUI5sgbIObdZ4DfEQKM342KzLWmjn7o/96PLuHQJ
B1DT1URIl3/Dki3pYfDifzp0WmRFMYZPo5Qwa/ETUvJ3BXlaXPXdcQkz0ANNQE/yANOa584GvCT8
KOBOlnSfOq5RUG6GJ7Kk0AQUmNWoE0CObfSmVjO3kN0ke3AsFrUrtSKoJtXTBIIAyTc4uvRgMZND
iJssm5uJBGZLHHYRZf7/zUuBuUIwDLfNibpwGvPbP7MFwYeqgzMzhyaq0zk0aa58Nfp4qBDbMX08
/25O/GviE5UAi4gwooIWFNJKtseaiu2oR2QYnN8xjwDzCrExK7CFvYET2KSATln6ylbgjDshN0Dn
AlwrB9QbWny1r71TAQbEJiqjcfNuS4Sk9HM93h9qruU+rtJ5eZGDDh8jrxmh+ZnegSzCfz03g+zt
gqnGRy79jHyBs8LE64LnZ4TZ9livQ7BdLAtljdIdjHpK8mzcN4PlUsqf/UyBYdjjvOUhej45owTE
qJYoTKMgR+hf7NTZZAwP7noxIEJpRmQLpKTYC7ZN4ZrSJPTd5o+/lMA60Ovc5TlVtGqsfHa0fQ28
u+xbQmJNGr0saaJ1GfZBZq7DMHl1gTqoaVFbS0wCbF7eUfTXH/17Uxk+alKEwS96oOAi++oX7lCb
qVIcNBJyGifBEYziHjplk5vz8mAsL9nMwHRvkr3ka0xTZ+enneJ9kREw7ZCl8K7WpP0r3QdaLKdL
3OlTOCr1EDTFHzS3absa/saJfV5VW3RlepBx9X5ECQUbAYuvsZeGzc9EUMFjdcgb90T/IYvXohud
BG06oBDH6dEKQs+++A4iyh/FeotpBwPfdlfahid4B8zz3lZN5QogE6FHxP63sWI5Z/DjUHo9bJU3
co2zIGPGRTcz9/SRvfsSZII/I9duEBwyT3NPcyyGyhZQ/4YtpVTk12+L7ixYgEfVgUK0Zyj63LMh
dSviVJIMLc/ZcAZTnUGc8UavWoGuS8SAW1+Cl9TvXZuhNS45Uev7mSCSjH7R4ZFwn1Xg4AqCUSiQ
SUz8v0TW/WUl1ld0qQYLOkvNN+0FswjyVkNRHjestbJqOM/zqAPqve5w7lMF1k10lTLeXc1CXeIj
ObVcJdH5hJFvT2f8nJFZKzd6JoggblJRmFerntBFpbMErUNB1igzv8dAX5YdxO1ehEWdY8pUf5lS
IpPt7qcylmLjbA73nF8wU3SZBfS6Y5rIpoiyTQjl/Xr+NhMuqSoCcbcs8xCgjoqw1gjM1VEsJOnu
Ii9G1mNMnvhCrJdaBHKn3bUnkPNMI+v0uXKn3oC9BpjfGrcTpJPm35L7fTqwfkB87egeLTeBIuTE
KF2qQnC3H0tXpylYzHz4vtdwsjMYZ0TVjdHCj+wciE0ap+JgnROEh8AqsiM/vMV+J+FcEzGg6BAx
Ped+SfuR4fHISJhVIOXSXbrfoC0qZBFi3rWbuWU4udFMNRPYXiPeNHn/2hce2UO0DeJ1doVzHubO
psRdBIiO/MXo2u3aJ8W16v9rYIFiXz4RQBzLlmWQTGmy6TqYGv4Y0UynX5dFYBYdf+XC9mL3sIrv
YnRtV+xmVQmNSxR339Dn9n5kR5HzqfoJ3i1HylbtVjuZFQhQp+oJ0B1/FD81VrjGCulv+huKafwo
lJbEXE0SB/MXoyZjc7ZRgTka8+00+Hqj8scRzO9CHKQfWVTjzpLxr91S1CbKULe6UX1o4gchnpYL
H7k1g9qgv0yXzpYOtrMNfutdf6qY0i3XObLKkw1JofdoH+yLic6hgV5jivffQd/X+OwH+AilkIp/
GFyxyiSNhm2x5Yy6hWJprATycvAFEXZhMnyFPrLrOXlSC61S0jGUaJJaMWa/YqH/fAKwqPrXSQrY
MSUHEE1hGV6gOYpMleiPo/Jxz3tCZBpx5jvchsXJX6CtVFsFz4SQuzosytzKFTQoqtFk6XS0NAOg
UXW7syvVaPz66/sT5BEsFjT65rzcsWNbgpnd/vbpYuu5d+pjCiIa/SI9aArSpUQHFCeTmNdIq7Nt
iNbQJb/OrGyOTbc+pd7sRo7HyU+q9ICb9vSoex4anLo67MCzuh9PnQlxvUQOk99MEMFI4iwGEvdM
MBbXYQ0evD1jd24xYaKQOeQAWpOn0CEq1TYgZ5f7cBoyImziOULCVSTYXWlHbmRje2Ub4iEAF3ux
p6rFTfV3RhyBV+KSIzdXAUuUXCQ2UPIMA51ZxJQuEUFPvjnA+cmTp8/oFUeUfbmevbs4W60SNWU/
BCpBuHERXJowHnwLI6l71sxuH2oxaXDp70ERwu8Q1fH49kVK54kOBb1bAprouVxrbgTdpXKy6Hv3
YLuchGxDr8jqHHb0mVUwOFAChLuS8FL9aWDtIF34+I62pchHT9/pn2PgOwfXvihmSJEGKLzdKoHw
qGLvo6iyL1kOEOkcBO2f9QJDlcjQD2JTr1cO+rarIUoZPzFeDq+DGHix6KmxET0r+v6FKqEvhEz7
fDUxTdfwo3YqRX50GNPQT/FkXdDMFST+0Rlp8s54SEwKEs25/erYe11D3vsAu0kKp3mwKz/J3yFB
VDHoCwdps514vMst+14GDiJ5TFPM+Fd6ASZBTvZG85aYxl2cPuG8OLHtC3GyiArhMATuXIRsKOaa
qAW6tgq5r8Csz9p/Nlz98w421S3Wn0sfjwHll+SJfZmS5R+W431+ymj1FRytacfyfenKAW9Qfpvy
bCQ63E7cFDo3uaqOweD0e+uz8S8hgdDxUt8ET18d16uX8FzXjW4/Ug+e8ZaNe8ce3UcHd5wcGhlO
A7tMfm0QusqxU7GAgav2Yu2YPmsc8py34BO8X6bQjzcXZAsw+TxBnXmdfYUDE5yRiaCrTeQF6nI2
duISnxnCMPtHPQxSvIWapTATsmq14Xg89gUkCZVbQ4ADe29RNN4dxEHaTC6U59EPIGnquAGgZwCK
0OFxjSLhQG6+5fm2beAUPGvMOzUClU7YDDV84Iv0cUzCwLmrTJQ4LmbtUuHHTeGWBCvqDotcCJzr
HktuQCv4pmvf9igpmjaf+zs9b7lpZNmXhjhLWMiKL8RL1SwaHwy3TwJj9sDi+0oT1q2hcTL9DBxv
I6jtO2CnrQuAyPvv1AmXrn2x4gJnf96mtdGDLvbGKF/lMXzBR2PSTyWfHokdgDzAfSywMeX3/RDR
uWHIppdR1AEBe0JR/8CNzvzVtb5Fj+f8Vrz4bnXPEOnnqmdWLq2y0MXnNJ0yF94XcAP1VfnokaPa
t5NwxccBbc4Q3Q2Ohgkrde69YtBHbW3Z9oq5KTcIRO1ZJke1W+f6GiVXUOGEmICIhHN5bkrA2Tty
8bxVi48DPy20L/VahkXcFoS0NGcZefbCvFgeUPYJQAr9EvgYdRvzsnPLnCpFvff6NBXWSJ+dhmi5
MGIlyDpX33Z0F5uf/OIqC1qgo1Lx9o4GCQC6K8lazQZWTwWx+GQlwwOTVRvl4MFgk/YsQjqHZ8aO
2c1nNizS/4vTGRQ3uk/9kACY0KEd3m7+rIbri0hzMJqMrxqyfNmwCqYIrpW5LfL7gWvUhz+ixXUn
QaFVNudbnuSDlrHoS8681q0TqK7LkKthIa/LOOCUi/wf5w9Cyhz1d5D2m3Lsd+HgC7fvKpGtCvRw
ZGQk8qlWuHucSqEC2RU+GXZ1DQlBoi/yjNl8dmblLH79pgoXmSsIZnyHPZlj5K7cANUQ+UloDdlt
BxpBIlhMQ1MzCsk28OiZCgUWRqkPEWf2092IhDhgwptXFBMiUq2KdJ6eTI7m1VPx4LfMqTVYyPpZ
/VV04eDa8kA3uZVxAHHf6Z1WNrHpxYfpWf9ZjYxGHLWiqYN6+ECdBXKBUbeZeSkJG59Ds5AL149y
/zsP9XrtlTzIGdELDnYFPj2lmIgP/qVCD/UtUuX7KQfeEg+PGKQwTb+REx6NGi6M6ARuC/SDyNaF
uoa0CaC+ojleCdLUccsp/cT2g2bwnoPkxCz3sT4oCWSuZIlmNZ1bGwN1G+ypu4zUMUbdId0nyX5Q
uAhdXiihWVAQA7SM1FNEIGUWw/TsjZDRyq3NgWrOB2utESeQ4KLHsC0LDtSFk1eippv/KER8dPt7
O6PLy8qflf6b4XSYAw+t+jzu0zm2VeKjePA1ItamhRvpeNvtE4GDk1jyCdFlqJXP46A2CeozwApx
WCFiWEBOOLET8YyRxWfxp9hSB35VW9RI8sMi8ZG6M3vYOQMuLVtoC9hbu9mW3r7doni/Xqt+ROH/
Ox9Yv+xgfZuuxLA33KqkEYB58WKs1oTibKMtFysG7hDz+45cnlSQ6CjFBHXv77hi9EkTEx0QpoSv
Xi/LGfYQ+sPMExi+qZqURCldhHFdaoDQCZ/S0M1MD8DrQShe3oprFDX6ZUvIDuIcL/RswIVH0p/6
bXaHcKtHzpCdxsoXXgHqUXUOlI4sTf/FNIQwxNIUlLWNnZ0akSlhVLVBH+wTGu9KYQeG+AmHMmSr
4NeVw2LbNiWXcic+pIL3Ruyu7G+5leXvlorXkVbXqnMg/ekRzIc44n2kE2YmnvyfSYVQGeq8S70p
Wpqk7REpkys1c7AbpBeDV1t4YnE4q6hrtKpVkyW8je9ggdlu3PpCv0B57IjkB9CU2poTtfR6wlCx
CgR9ttHTrHhEZefTXah9CPPkEfN3YCQ1rxVHTm9g1lvZ3J188wMMcYTu5fQUphndxBv43B2HMCMH
ieWb3ciBb9k5N3AzPfjVNlqfqkGJ1yUTuUP6Fqb9ElL6K45en0MFwFT8sVtFlqDD5diEvZFSLFFp
rhjtCe/Jo7Q1iX/3Ch7eQvq9eCHXXUw6xykx1jE2jOlb0w3u2964MZMHCAQdSPoXNvOr+qMABAz6
A7y/qIx05VZOwWqbJJm6FwxauD6sG7jfAw/wbLu0Mf+bTneL7XwRpBpw6COZSf3dAl7sdacaZVAO
fUIGg7djTNu04+hBWD/WiBT//Jygp4e26c88w64BHHKISyLkI3f1dxl+KjuwvNEOtCh7zDV9iziV
/FgPZLF2qoXtr05qafWf8OQ9qtHZrX0CBFHWZJhB4ICR70nhcNNNslQjG09k7CUqvjD0vUp8Dgqm
id28u1OGJQl76Knr7kzTP4/huYYkKTpQNICkzIP3nqxokkLPS2yPIqyE4vnmUVykS95+HhzNvhtk
atKQiIxIWmGi7TaM8GKCG4v6+4yjzkLMJziBzok+WJtWkogks0WSzV2YImClE5ylY+2fFUb1lPeF
IrdpJ/UjfdV8NjxXNRmeiH9bRIqvSK7XJ/c60jnHw6TfOlO8A5yigGth1dT2VQZ8jnE/I05BXGWL
fWoIjTQ7tQxwnVxNWnrSERiycix0sakoBl2mYGT17Qq2XulWJtVg9WLh+ynnrgxDHpTyjQmaqjAw
i6AwSTafnhPqNbBCwlzWl4lHTCdRDwo40ni8+wzST6ezqLKQsxQpFqr2slWGnwupergShOeXOwKC
mFGdv9Y2wHWAt1JEvDeex0HgLQNomK/QZfzWh/7Wj9QP6tEuOax3bFSAeCmnxr3ZSWsvfW7xmwMd
0nbjaM9qEDxSnLsWrSCOv3kru08ScoFeqUFscoVV2TxBGC2GE/gS5oJ2PYhYgOLFbs/V26rxnMDh
bAG3NI7eH1FF0Y2D2z23QyvouzsftUUjVdkgSuDtS2Y37+PXFJYAdxYCAy6kAx6Fb7j6oYU/TEMP
FP+QtLVegJhS9ExwvccaCdS2R+0ZEnVWbJDRgh1dYyetkLO6zNQ0iNF1tqE1+5iQ7klcf1pE8gdE
U4YOZVVpniy4olqwUw9m3fKLnKqIkcK29JSlPeUHOg2o5N+EbwLdclvDekV/y7EZFbCm6WnztRyR
B94lSr9AI3fY1AVaMd8JBgGv2gQ+gekhcNzVODAGhDPGkqb5dj5qQwKnO4/VNnCOPX2LA849y0lf
MAU9dKHedGTPbiVAizWfTZSC/Owo8yLGAQq0FlgZYZTutaqDERtQRFggt1NqsvFzgd8BCQysB1EU
VqWARCzZ3msd8xC46XD9GDC/wf12mmKFQaGoxIvzvmHjlQMKjlxAYdmYOkjjbRUKeFQ7pc5vB5fN
U957/f8qhEVWF3p3KJdXTa6823KBirtZglt0FnKfEQNDvpQoOmw8MsrYu5b3PAwMIjcR0VpCwFkQ
Nbld88+MSThQF4uwShbA+cNOWTCvrGOSjmIiXIu5PkdxRoCbiQ9qA6Eq62y9uWr9Odk74Al1uWOl
rQnqf+w9qkGKmrVleoELJIA7FmQMeqPzDeXKhytCBLxi8eXimdUT1tZqK4v+uivIvDorwCvHcFNK
pHDVFGuRfkeX4nwBGg/jJyU7EBpHJtUSj3Gzlq37KDnwYOar2cInmD5znZ7NU57AUBD5Xhz1y1ui
UGbrtuAUlYzo3ZnZPEOc6E3s6tsZPJHOmG7I9SwkFOUx7rLgd7x41AP/YwA+2/7ch2FSgdG2Mqzz
388wW31u2lUldL7eUHVUDoyh9dR4MDRX8IKXh/nZiZmmWncNwYg2xQ9E6XwR/r4stfvMNhXlSQYU
+Zmc442la6ZhwTY3+Bd8Ce0r5szUs1RIve4gqVzJRpXl/6W2FofHAHiX55f7ONh3yq9dDBWp95+o
OR+1GvoihIuNGAw5X2fq6m0VZqYJH7vH9lNxX2COl8bO1cspkl4FhAEKJH7F2qdAQzgJqLDfksvL
bPankCPpFua3uGcAIyCm6//kOynAjU2oeGpHutaSHDIQIRriEJiPmfZL2tO5W9lroWjFC0q6eymv
y+AMCZZVMrlqOX+ROC9iUr7yPArQl0aAVf9PegayBLhEJFa4ZUmaqkm1DjIe+B8Q+twxSD9kQ7L7
TH1uhcWn1KwhlsjoPxm2D8kJOYZROPgJpDZoZlourxicD3qqzHOgBhL/LbJnUgbUBQGNyAfwd0Zv
rqf0CHQIr1JxJqBORXpz3ghKQeG3XtSOI+hcET+VTN7+lz8i3ULWyzNJy0G/LvkgrkEYTRBdxVrb
9wefM5Lv3CxrRzRr9r9+mfU/T9ZjriZTSXOUaNj0JG8KjzY/4zMIBhrKrFr7r1u+YfnT+wDuQj6/
9s26L0HkutkjYKthPwC8xBUINgyQVw1rxYLT5aXKxCKEr6XCt76AmZQUl4ZX/s0P86BJl9Xn7Fmh
3GTPehmmedEnGVwsajX3Z7lcFVJDI84Dq9n+8lNAFdyuCIIXTWNdbIYj8pLwzbewQLk3foTlKnEK
VTZnvo5jjjuYpsXCoCMIJ7BFed7cDT4iBE8rSw/W2wt1OA60FpcqW86GlWlwZaAwG2DJtattfsM9
JBi6PTRd6i96ZWMqya3NlOrBye3F7Uq7xrtk7PKDrDEUchj6Ho9n04NFGBUWyc8u0tH7QLH22Z5n
A/tq4g7G/nF2mU8QUeOqcJE1lAPDTeitY9rKtF5Qa+5sOpdxjmf3SGkSBDl1015swSLLbRZsgLVy
5eQaeMI8bf2HuJbJLYBeUpIQHzjrwlcYi0fzi4ancuiyoO5AIKiQ9+9czwJ5Pj7tYRs6GsweHhd1
KqdpbPr9ETOBY9yPnTCmQRP+Yo899lx3uRqRbuXnRObTYj2Pg1C741oCHJt7YQDcWvtwdNHwhVMz
FU8TbxbX3EUD/9j/6ebMsF3LxrJ8m4KejI0DOof4b/NvbE2uwSRer6itObuOrpO9vuanAdYcQ9sj
IoEbEFgwODsvuarDR+00ZhJTqAeAhUmxLvbYAKqvjYwiZIdTlHqGqyfGWP68poI4Zf8rlmgS7vRb
Q1sfni4WwnqyYhxxtfWbxhLhgkIi8n01UZf82v9LJS8x+qoBfICJiQKqQrWGeQi+xpS3mbdRx8RP
ZaczDYrFPLdo958AUbJc+r8SM2bEr7BxzekGMdx/gNlsL33P3voCMzqYUIdp+eH9vxLRaxszNxOK
vA+mUXVbEHwuZUgg1K0Dd5pPQU+GwENbgmYjNb7snxeYdZtYcYNcYyFSxxEFMoGyURfTYN2GP0oA
a6suLj+tFpQsdt9fMl3dnyxxJ0M5IM1knzYH9b0UV8HT4MwbZV4/mSpHdVB7hK4zHfn4j+PiqEmS
zrYV49rcVY+NBE0DWTvmOpQMJh1/jZaq0HiWB06Lg2zA/O8pkyPPOkSj/nTt1t1G/YarD0AGJ5FP
6eVPrW9OdM0Z2S3+s43VZOFBYLLCAUuOMJuqREYEP/E2ajoFNhC564SP+Nfr95vDJeYShE84pIv3
vRy4ARFcVli1WYwUOBcnE2dFkbzFJEWScs3l4R6gQirQJqA6fjLk3amMCXoLtgQpVmd+2CDGt+zr
/fE+Ru6ldMWKUsINkvu9gwRNMEOtEyfcnAO2srKMzo1STDWhLe9tUBFL0GWBG4RjUdbn7TnTHp9G
J854ZIBClOQ8cgX0ErVFB1CUXNjvjmHmf/BstFCUHbSN+k2zlAlcTnCpGk8s0+MnTAwZcLwmpMq4
DoCXSaETem5rNMonnYp3HeD4OVLT8l13HOPdGjILs4C6UvGNeySszd3ZbslBQTvkQOiV95V0lFra
EICBl/eaqcEWphOERHDJxDyGSV10663YzfKIJ2iaBdLUoCxRL0HwQ23KcR+9iD+7Bi3UtaHamG5h
ilTW2uGmCJ/kmH0WoTaK/gqfxT29i1DEt3CwQlMAtM8U7Bw39TjnvKp6l9t3uNqbWu04Be7ChEVX
lkLJNZgyE0EONPfsYxSoHLhASuFVVlVcf+H3Kj9veGxsvO60RfQlLxyDIEbtbExStw8sMYQIczyv
pWukdQiHefyBWOEPv+SljUKfOE94oNYQfiORILYx2oW4xRvhBbhKytVqsHz4vBVzkpk8ELAIzSTj
wBAzSzEdWayG17LW2A2GNd1BwXtf4kiWqVeQ6jygJQtPa8J+cBnH4Omz+tnCjBXYlS3LnAwarjLW
Vdpo0wouSBky+xxAXcs3rF++Sia+WYs/VzyQmJJw2vlDttsmW1nNEzMaUm2kht/1Zi4XrZcUHkSK
aJXNPPTLvnjGJ9Is4CQYxBhwHSPk1kmV7dNUs6axaKlr+KXkx1YOnHRrkOV3ryR5nAh6KtO1Sfab
g6f164Wq0YewunJLtJolYP7KWCNVjHbXaKexXCMAMYlt+sxFkoTFaPfSLR6hC+QQa5D+8C1svWVH
JbhB4LE/rPKfkRjlE2XbKAMHEFIvsoQcKV1PXsGXDGuZqiigvMAefGP+0wruy7WYGA57ueskRT8I
1RpSVUT76YM3Y2ku32MjCxw4XTtHD36Xz/Rn35q4MaOgpcXx4SGDdtktEt3EGZU0ym8yd6u5SGZn
67lEKd8D6pdhTcnjpk6moC9dA6GF3Mrhu+vW5P3JCfJyiGbl9lxMXuaQMT/K3pNBKkMW22EZ0IL1
0FIg0bd2nkJy6WPs/1O2Cinv32bMmCzWDfA6yzly94PNjpR+zxYLT4ffjP8UlfDPheeetaNKJ1vQ
vAyGHvmcz1ti6Kqd7m8iys7LZBV+V00WO9TYBKCS+zq+npSoxes69DmVsccLEFHBuQAlWx10gZqH
xHfNgp7wMaVBJQ30+j6gGagxMV9Fgm/DMO93L9luPWpfA5ioTc9uvayfuey9jff40pOeYjvubYUG
VJO/lyC8kn6KmZxzTkyO2sRhVU/4JvzUfioJbt2kP/AmaiN6F8vFNlXJADl80+yvLLcqZ5LqFe6N
GDBycG+Eh1TQkcuPER6hUQyckLJ+Y9Ax2D/0kG4y7Vl8f1ZOkoDixhgnasfu73Q4BvRH+5Sr9o7r
5rNKcYuGQRbGfvuM2znARP8SlgfLbV+3PZoV+sBWzR0HD415ZfXN173Dk0TjiWNJJ1myP+GnFnov
kiFSCsYCduUVIjUmsffluFIImVao910HosdiIX+Wv926DE1ZDKsnRS1P2RDwXjDQEbpVDg0Xx9XA
qsIb4Z1RZVeXxVsYKZEyCBaK6nC/nTOZ/7XlVGR/gouA8abYl9AqZ+3Lu1Vjxf3Uyfa2gAhQh9MZ
kw1/CzkyKGL6jnXS2uQczHh3MReUJsvODg2mKB5jUKFwr4l8UFX/+XpwX9fiSNN/DzrUfiUVmays
Z2+N94w4hChdqzmeJAjgCTnefHQ2dQ7qP/MQR5LGgb9AZ4oqJHxrJNtZQIewyziZIiL1INHII88i
PUlyyd/bA09hINKntFI5iSVGuJmXSVS01456yzKIDeto0qEc0mmcZhD2DQoAZm0qZ5eIa8loVyXn
AYgIFi1TfJg8CqAlAVnB+Z7WoQ0HdShwLWpRW+S0PFGReecVyFSRtzzUiCuUOvlhFYz5kqvspE9W
1dSR3K0QlhNunzpNiJ/5XKyoavXJXiRE7ahxAm77Zr6uCitFweG9pj8oV10BOs6MsmvLgCG01s4L
fEWuk+iWX3M3XuKwIZajdWpuilSfSiOSfcWHyzrrrkiZt15s2EE6ZJY+a6EJduvqtFZrY/awr/Gn
MUMjy3vx5xix+Od9/SDk83I3zbJObeNqRZK6T4aF74kDrZKgMNy+3oVWb6IUG3hH2MA6jVAyiCYK
L23HFp/jjyIahs5tIs+kShGlprCqPbSzequwOXJ5o9HaZLUSifWrsftpfwjOZU8fnMu+m16OkalA
5C55ALQgGK7R+OPw01lLOLWPMhYHB1oSn+1Ps8xYQBP+6DYsC7mp+L/TF6DqVucdWE1d9INUxVb6
qS6MHCpsEmCLRXbZUmZ0zyOta7O/xKBHYv2rqzmXoZFiI2m90f7ywyGc0Qv9DHRwRR/MdtRP2/Xa
JpPPS3wMDnsQQOknDPOM9yr3TfAaO3emROsy8qi5vghs62v2MlzZVRDKCkxnFRzKqQTWk6xDexrP
gA4hb8+mEJwXkPDvU95toy7x6xkJwcantmG4JmW84MzLonOv3I6EKbklbz/iI+UJKuLvFr7hkkNL
rLWRKdPht5afuCctDy7kUYTNgH7vVclAoZzibOkUqwZJ4UKLBern/5Af30by0ghqiB5MFQzoI+v0
CHOIXbQMqRQ6ol5Fxksvzbpa2JuAR1WRawh7AJntgKuffuj2qYV38RrCdfIrIgJc/X9hhnFgQI+7
gHkpz7Ndru67NagM47MwqxVpcbp9OW/gJoImo8QJLqz3TcA8AEm89ijkK8c+zIqgRRgNOSHJNpZ4
A3x9I4eIjjH3I6DmHR1D8uiD5E0+zpiPIGl1lzfkrd5vG6u9Yqm8PqmlrUjx360kEOfKgQKifodW
U+ggPHsGaExt6K1u24KcRtFRtF0BaRQBFL/VlfNGYAn8+yM1GGcOj+x72BL078UMgpre6cWSgaAW
jt11jWmG9y9XUSMnb1m/3B0+VpQ1W/58vdroqebkmG9SYS/2c9r0Si5C2m3MOjZerFD6TqxgGx2I
2fODIJ0bS+FpPt6UZmyMiOEd9SL6slNwmhqo3CUvcWx/xgWXu9c3H7inAcv2Da754FR+BDF7wVJq
N3JVoTfpT5+CzQgBDOWo75Uc3PnaZNeD5o+hAZJ+Y3ng84Yaw7GM52I8zHVYgtxTfwGifWpG1lgo
T8yh9g+7I/gFSz9HBKjNTuxjq+3lFRFDb1iuvNFPg4a3HkFPF6T18ypMEMQ7jBJGy2bmhFS1wzhQ
J0CuGQBiGE14NCXiecg31rP21OO+e6bdEDKg2d+lW1u/k0vtPKewLJxoU03IBh9hfa118QSp4fWl
TJUNw4NMIHv0qu0g3HW/9toBuxNKwS6Hh0EyW4M4o1zJvPHoqBicsMa+d9TYmDdbbcCPyvaiXdiv
+wueUUlOItkVrtBSTLwLMZPcGtyMqHd6UuDvOpJM4fLHPef8ygAcJQn8yHDcM31d7v2k/EDtIrvy
2N5CjnDp+wsJpnC3r8IBLafkXSybkmG2MBgn/KOfQ+AGfKjQFM8nyL8zXVKKd1zry5l2rN7AGD+D
ezx659ZtJmB2E5q7lzWQJS/+q8zQUmGV03OE7muNAcyb1ep6mz5ZmBIUZjmFRqvg++mXQKI+Red3
rq4yFfE2YWky8ksAKGZzREdmg3ASFRvZy2xocJv7oF9xHtkHfnZo8X1kO/rd1cPKJ3fg70VAWE3R
qzveSog9hMAysKCkz0Yu57zYbF+MMqpwfxYJT5dYq1DcUdERBKRkCYDHzabNptLYxwbCd4BP62fU
gm2bonWq3w8SVwwYTl7NKMmujMiTTlj0A7zoWt0cyOBp/iKZOQEbDUz9dAKwYFuh1AWOzUVVUPO/
6re3rDaS7zsqa6O92q8sMPeemnmK12JHy1oQVvhb0GwdB378rX8uHmjeLiJFoLeJBDrqeLA0PAYg
shhTK4NDcoTk5fhdMDENclmdICABUR5cTlNMF9MXomFvQ06VFy3oo9PbQdBLohH51AiAU/OVfUAG
r+Pgm882baEf+rlJ8Ez63/D0vNcScYcfrgY1XTEPa41VbIh/VYjOtNnp3eNIvFES0T3QNjTT/HEO
+eMrvdvo20pAHK22k3j09ue1dfb8dGSlkfe85GBVSNAfBaZz//qgRoDhZiJOm6TuomNp1Ulrd1oD
eRPEi2+ARJP5irgQC7rsHdzjLtrHC0wKZqOTaSsgEH6TPKcyOXk97UZBbnN6PzzdbunHAMPPI384
3ixd+exwm9endH3ri+JaptEb6ygKK/Ih5pInykO3wSmDx7xStybahExmgOilrSikcaTR0Y0Y5Au+
J1LVqjc4ihBmxf8spbPSkl2/RDbeqJrbFPPIGVJtWPEXUm6w9A6C611wwyhZwDpwfgjTnONEUAnO
m5pQoEtCWKR9wSudPTX3IgE3op40vqfmIe5TlspVllYMtsp6ac0X5EC8PmOSa8aZ7n9xx9E6gLnn
n1a1M87WALzPYoDBHsts/0w/sUbpWY4bzPND7MZrzlpRZrO3ISYjOkd1RPKvKhpGB0uq/xFrjs1o
7vt6ipaRKh4J8GwRp/eYBqbF7iCw4+Y9P7MXEe00pixTAkEE6CrXe3LPy1h9E9V7IgYEjxwZyNXO
3A8H95khNaGklSLYM/v77MTh16NG0tPL+l47cqB+QgsBNkEbGWxIOtnpb2Nt+93k8sO9uQxg31Vo
wA9TJ0EFC1Pnxh0P3+hCx2u3F6CwuTdznhljt4b67raEr1D0b68wy/KC0afsqN/31ot3cpNghk/z
h6Cd0daX4bnMEBcKsHdVKG/C9wWWBl7J+vUxRDKJhNLx+3AL1se1tS/76On4w5X0MSoPshc5lbfs
UN726u8q6ii48iaKHYjRiBKuZuQIlODWxd4bZsXL3kKyJDk8v6iunPy3dRlimrqkxTzDOn0fiHXd
b8GjAPf/PrdLnu5yV7+TxIfXXykKq78+/w7PKce13QdL9TGjYkGJxpQn1tDlVW25I+H2ygdog1TB
UwlrWVIQsViivBctZa2dGwMttlPAPubTaWGzpB4CR1tP7f4uOY22C7ig4pgRD4mMuK3OyWFQS0Dr
I4RcCBL7P6a+k/S3I18maJVdbMEbiklRNlF0FJH+NsPq52TxHdyW/3YeK4rHGEqdScLNc83hc1aN
AQzOfj8ruEeHco62sTGqYo+reBZ8lZHtbe9i1X0NYoIsnXgLJ7XPGL/UQVTt74MoSL3nNXdwmeIP
92Yanqd+lJMTfVa67j/polJ1AqZ+ArX8JT+riQkzgyObEKGcnfdj/S+v4Yzt9FLw4wJDjEvvW2C2
fUmiv6yi10nTvGBuXxlI2H5wxt4oo3pgJ5OD3mHCP0SpB1EZtK5onPedzCTGA+nYEJU29snwJDj9
pikfvyfL6+7BQSg4Ei3bcB+T3h1ew+IDEuHVDThh3nhyn9JWLHI8KutLitLKdrucok2GClavlus0
qTa00aPu0ZdmwWHVSwQUiGk1rqWUGhwoIwvvf2sSJa0leJQseczdFA8dQhEGXm9p6MQIhChwqA7H
llbZ+50GWP3UBJhiwud4v7VIoyzGIRon7tuNLUH9j+on5MUlZlqfPkPWCGMa5vdYFnie7IkmsKKi
lXPug5vmxouD5I/LdJT6JwMBJUf/BqBVL20OdNYQl9WPzIsJjXYQRKyGqIaYsSZod9ihkWNSGTvn
+kIS2M4i9Iydg6tVXY7bbX8nPL6dTfRgtFxaV4HnutqHBkUp37E3oopVd2PswB5DN16le/yWol9n
OhYTEyXxn5pOXM8BTSaIQOL6FpGJLSYdQErt734x3lYxGPQy6s8ex8D0L00lJo5BSUA9pnnbQ2tB
6OSCz37MHR44sFcM2z2NajZOF0Ix8uhkVbRO/FhjgsJcIuNrI1Z+hH6VAvAzF4zOmbAqkrd2FD9R
Me1YB5g+nmpI+izAzWuxPqeJgqCCK1xw0iBG0DC474DGKIGwi/wY5YsX0dSEosZPfij//6/ZmOHa
Bl7A4XNCJalUOyg4yTOnz4UH0PqvZjTPXpHrkFCOlI8U28NYAJa6frFu1WDAhGMfZ0N+JMchc3ft
vXeWz4b+bZPrCVLb9H/ViN26pq5tVRE9DyaDSJo9o0bxe/IlIOlU3Ww6Zcxm3h9+KRwRaC15+pkj
pGbfj9YhLBVGkU4M/3xrdlwnZ4yBhPXajv66uklq7IWa5rNXDgUiq5tVs/XGjZbdtDZAyI7MH3Yv
IJnHPm08OjagywskAbImW77fZBqN0MrBzQE2h+hlFNP63OXbP2bKQL7Hg5QVqPuk0Uuskp7Y9rMz
cAVH+iqyu0cTit8+GH0kQaX58pa/nuGLxd5TFi6/g5IApHd6H8GLjdZTrY+sgcqqxS83dTdIJAcf
414S9BhOFNsRMkTyI9HU7ZFQkP+LsE63NGhd/vhwsg4Fia+NncWywi/AO0GXrEEMvWiuv3PL6/Wo
wRUCSlGiZxPeH5nsdKiW3nuzFJCCm4bbgC+uwwTZucjCLW6zX1UmhFcEl6oxinsnAU2+f3CsEKuc
RbTGFKjGdgkrpm6fJ+c1DHoQ/mW4NuEvK3ekYVfu62id2YPLS2zmt3gBl2zAwvKoT5XG864Dh2jE
xzc1EP6prI1u1McdO7Own+b1m79ZBWKJzpApRTjxAEn38pcUNZxcgZzMnUf0YZKg9HZX85MyeC2t
Z2UNoJAwFKG8XLuUavqu9U/eUwEwVPwtFApgXhbB8+yC17MUxiJix9dRv7k0Ekq4gY/itW5uJq74
9rSLPyqrx65yJUIaHIX9su0FjBS/oqEZ8rTVJ+Q+FyP80IYIH7f233uT6quoquTj+5YbJ08MANS3
RywhoAaIu3hstPiqm4MSRzR883owKxfJo/mTa4MwuUVjgQKHcosfbKyUOcvUqknYefND7qvh5eo6
jPJ4Rgumg9F3b9z3sZgkL6O9A4CzqOYTtDzlbj6EMrZmUyEKFUNrdaTgPdEAkWNZ0NLn5iFGzo4E
DeQnGs5f6Tsr/ZZ+E5Sk60AE+1uTRUBrzMEssW6TYsoXbDrKQjtFPIYZkJdkscN4V2OeJTjANV7o
5y6zFwdZMixKV9OjQiHV91gpQWDZHFher+cu1YmmXpDtk0KBzKRra9KPCPKgRhRc3p0ABvXQUSvh
AzmgJKJIEZSMwKFK2t6LyLmo3NilD74uBAOGcl+K3d3Lg4m+RXqLHJJSd5MevuAV60Y7Td/PFejP
zQPc8x+iQ6EQYUNHHN6Bld52j4tldWqhjE0UhPwh24Lnt2tCQtJsPVxSBSF4A4ok2Ag0SI5OpPoz
59krVX5lSM6khwGj4tjKcGnGzEQqS4B0u7qXdNyKq8HhFOEQD/q0hOLKqz8MBaJCl/K+9x3/ijOH
ybJxpz8RNfD+j6RvHucvmjwzIV9UtqrCIzRln+/7u0jinXd+XHFSUi/LK84tsrw6Q6ni1bjQrAQg
V8LX3FgCZuKJXe3PjKHHvjMJdjAj+gUM2rBIj6Hm/xN8vXDTnjiS0DracF5b8XVUdhxWbVqfMsnl
RWDUTXZKgGvxEUkMoECdCr9Zei9I1Z9zyTNLew7g27eqjvjqtD9xqOl3KOd9ooQih/nYo8cTWPVs
0b0iUAIxFDiJ9pKaDMQYq0a130L5au5pUsfBmtnHQVZg45fVLIYs8Jd05TuBTe3pF/YrgwSrtE4C
rM9GD49uIcay2NCYMoakUqqk55sbCe4mJsJi7jmfEk2YktMaKkaciyNWR272ctatJKG/vzgbDIl9
ZWccgDFy0qWoigIzvvpxVgfXqUYI0uJ1VVHHXHLUCiQpEa9bdCaEO7enmbDhzGRiTKF19bdPuxyj
3FPt8EBdnO5CRSu/gy13WExt2rBhjjBOAoFqt88G+1wBgO6xaNDTS3AYB13CoHC3v+IzPvkzG7H3
YUmv9vzNZQ2MYvsjMXwEA20iph4EXUDpgC1w/2twxTEW8QbYdd4A+4oUtfE7AENGTi7SVHv7o/w1
UQ1qW4edQIKOoZ9NOSWza5krWimXDCw51KP3gmcJVv2lPyiukecsM7co5TCsrlRJDw+UhPXazTNx
lrMQRSL0HfLlQFokFVJMH4zCAMsiSW4GPuyZxYA0oDdm9D8qXwa8q1yDgEEw6ATXt6i2Mx9X5Wrh
8F2vX3fYvbxpEj46GrFkNJLRSRwd0fcaHJ9nG70fxsOIVwJE3N9+plcbyNlQ5tfb61An/IV96Y3u
/j8ax04Vn9FBXXOBDhd+Z9yX200cO+J2dNuEjdieNr4Swoxo152z436GOGsth6tqq37Y4HZGaC8B
ywP4032uwje1nAh78Fcgn2Vv0Ml0GiptE/sIVWDWZgKcG+XMMOmwjDtzakia9q9y67c7JuEHjUaJ
fRpa9kVL5wRR0oLzFUe7hgNAa2uV3XN4PCx/zTzRqr2Td4ryDP6TqnF4B6N9bFTLP7n4U8YsXaVT
eGYb4dGIAX2BkGzp9YhiitezbgEGkyD5MSUKKfQEwnUoXs8sNbjZY6Zud1L8pWLVBJRgA2lpdtlZ
40+BGT0gbeX9BEuP0i5v3POFkeQdgeGBe8pTFEG47Fwu/LSyogF/U1N7a9eEXrwyLH6WY7yPxQub
ooGJtufLVJaEQaeL81KSp7TMZUZMqgKnQ6/P8p2c0BHfTqhptoZKU+HtfvY1llGistT5pJetCtxU
ponIALKJcCpHK3bSRdBsMZcMNZQ7Bi4DEL2eTckD0MPedmoNQK2qqjeiilHzJNu2QX1cl6b2G89K
WkQic1AoSzi86igDw414ol7KQrN3yGo8eRy3MXzGQGo6eXhSscQjviAJWmKFOuI8rqOXvc+1/y8+
myumw8xG6u4aJXEcJcq/sAHQttdAvBxIPhixcrrJqJjvJc2HMAMe06+KaulSEyMCCTsaGK9zFlP/
5Onw/dYnV+ryxyXQBb4HBP77WFH5U/HycXvD/L4K/hsSpdCcAS9n9CTtLmyIN/mYu3eonkuhHu3l
XfE0PmSp0EVR61+Pl6po7ZYPotSKq7UAERKyL8/GQhufHfbXog65mnTwmvJMLho2JuZXqXaZb6wQ
xTK6X5Yizn7ZL83dlzYTuOTNZIIPS/AcDfr2L701CXFZP03Tdn0gmUcnPywmdRIvGiPH/4DBOrKj
limpctkN4fCAfuIJPqe3nfYZ/k8S8d/nXAktLIKCOShIOnxaT1+AxCUy3os+v1LD6AtLVZH0Xay1
Rn0eXgoNsWhWJRk6Zl5bg5ki9z/2S6yd+/rtla+Ptpk+lAR2mg0zeaODovja61Rozgmbe3cwnaY8
BfnYbjyQe47nnvX1zaWRezbkgrbrrSvkbjOiF70vWDn/tXjQcAOhuxBrErmE1DSYlulBzXThimId
/cgrXnypOVW+H+zK7jIKVsFeZJoQgAQXBo0rk0qP5Erub/+bXErOayFno7dGYhkUA1qPeVj7pzLl
KdTHKCckWmBmxEmxtF+WF0Z4l7LqQJMb1055H9swU2NThy9zZks8tYpxpwDvl0D8O3Y3Y6x01W8L
qB/VBP5Nhx0JOw7mQcd1cPbiSHcQr7g6vP8D3hayRQe1hTAEA0d0u5qUm3oB878VqPLFDCpiyxm3
bKbRUsRNOk4eizMvvUCDhQdO/plRpOm4Nw//cf6dfIuDfqhsdqtV0gXzhYyW2+4or3OQWpiVWrcD
dVZCS/nXOWwrBaVDZFdHesM6leAil0qi+ISBu/q6cLaqtgMvHabFjRU8fVv9izHKoipc+z2MhOBE
JX6DKSXIPqpyVVG/ZMQ2Bxv2L0Zy71Jsjfl1BqxuO6kJx75QUT0nh9zH/lgbhtyeRghdLhaNmJLc
ZbglUgiIvH1Qq0CKVd+HEfXfWCbqR/t+7TANwE8Mt9XQHD9kN9+AqVlLmXy77iO6W062tBjapIw0
TssklC9MD+BzdFRDBmZyF27MWMaZGB1Dk2B2XkMmnRGxRFL2K8hR21d1aynn4S4YD/jKPeINCpok
tfUd9JH4ssefzsaPkS94z9D2cmZ1c7fQkj037vox6VUdW/9N496znpZ/jcj08M2cWSZHx1H5clNQ
tfXw5fL6+/ce6vS4EE5sT4V9ezLyviFA179rGJITJ4bM1O3AHE4Iqa14kR0WYwG0LmisAfD5SZh8
9Wi20M1lEkIt6N+/jDT4gv4ujGQ9SU+hGLznTVpHVx8iAm73AGD87yNRbX7yJCouwn9iJB0a/6VI
rghE8dtin7eAzB4PxpIFbF1Cn6fyKJ8Ng+jxrAIKHIoQEPBHpsU07/BjR7PL8v9jtGprJxjH5kck
Nd4r2WES+OmZhF55nm+26hjFrGOBq3uq2TVpUZ+GV5qpaz+KJ2f40ansaDo5vZ2j03Dzi8vDGZVS
p2kDiHEnteJm1MicnVy4gbarQQQzIkHtqN7WGxG6tBrQlvZ4PbldCVB9Gbxb+nK2MjBBZcKxwHlp
+v3ds0PsP2VmlwgD9FlcRUY2mLvNEpSEWv3o3otiZst+puqoCSZXZr8Fp09xy4tNFrq54dqK/vhz
K5Y5yl45T7MI07Pxu2tB1mQniiy3C4Vn7T+JJ39NaoLgmUb7hC+5t+MtauOW2x13tAdc0cpJvQ5R
Ks+KlgGcokzp6VmR7rEEBRJm4ay90tQhw6OuMHqWtyzBQ92ydJcbfeE0dd8TeRHHKDBW8KmKlvLL
pnETVjU3V/BV7+FqbA3Bh7bhdJONe3Z8PCPO4fr4AYFbj38GpfAGaX+DPoXQKDG8vMK7AX7KcGkO
oAzAU28rNZTu8uTd71bfp7m8O69FvphoYahS/nxeMFmlTG2cak4iTEp+/3Mm8m+PGO/4JCL+hWoT
upwDnmYgXj5o+ekT8B4I/V51EBVHHk9FGhf2LOwm6vSxL+EAg8FFgMRu3uvc82oxSoQ2kUHDHVFy
AR1GAvpSQO0dHtn2n/9ihdN4nvDHZtePyeOTQaWn2WJT69GsdPkqLHkmp/mKleV4Qrf+IIHibMaK
ZXqy/HjN8wcUTtz1BrhcCCVCD95z6dIAZHK9zwnkXx8cwuVGwiJUdMVGfazNesF7iQldqkK5HwYL
iOkMB8bhUbt0HgbOOd6l8ucu+7zxEeeOpusqPh7CRVmkksdgTbCjcxQC7Kadbfg7rJD8r4ihDTll
nYMqnYhv+dFhsghSPAGVZOu2XwTzgmWSh8gCrYv2GVtV8ji9kqIaUkjTLkzju9JmlF1MQqyixwZv
PBceF3FIo+A//VKfGg7wor6L3D+S2F54B9wCkCoaS/HlyKrU8TqCLNCeb4Q1eYtcW9suZtw711SX
P/3Ixx3EK1dIvwY+I34oMkKE6wF/LYwV5obnvhPCyeGoRLngU7DQacRIO3g18ebcD2NmUF7tLCKR
9T2IsiSf3ctOsp7fC2YNs3kFPzur+uSY0lrPB/C23wEr9u0MbV7YuD6PKhuT6vNaEqVRnfR+72cl
hvgv8BKiOFc34XHLuJIWLJMH2zUM271w4jmfqZZ3x6qYCukez5gsD+Z/PgPI6sjCbTleqBsWJAIn
G7k3M0Rze3T35T8XdI89aoWbrBm1+Ajr7Wk4J6K/SA505VUWcRmAe2/NHunMkBz0cz+Hjwr66EF7
1nKiuETN+KV3vlLISi3NBvCV3AGdyl3TSW+9DrAYrEZwKD+fvYvu4GMinb9A6Mc3mMWn2yeYag0D
6IRxvc0zPm1fgGso78U3qEfZKY0t4zNJkQHk5L8CnrvDL0SCVLMBSbZeXrZ/msJ8+Rk93nyhIArW
FBd/DsmYbPp9lD6d8g0/aqMrDHJkz2PUQq2u4ua8/k0hlf+t4mH41v23xQ30hsH3Y9YwziBcFixU
NVMScN5AL+X78v6RiryeQyHCihTbPsYMN2i4a8B3zEZ+/FSZJyr9UGNffUYPhUExf7rWTt74XL4+
loJTOvCNq3ckjfXtvR1vv6C8J06KDQzCJAIJ0NGFqJeCSCppddKxBC+WSsg1LrGcqoWUoEfrrxLT
cYEpgnIw8/y75ceRM8z3a2nHsPWZCSWsHktchAge++DwzVZ9hwlqVmp8WP1aGy6/kwuExdiq0Ua0
BL1ohsNKv3PttrHOxxJ85RpZEKijcoA6lCPpE2p3Aj8xCXlYpCm2UBde8CRofr4xid/05efIx6cn
4BBSXQnpQqJLEDRjSr7eCAtFVve0gctckY2hO36hz4h3o8yxGcNSVb/kyODSnAalXXIhaInR891o
Q1APN8sNuGwe8Pur9uflYrhn98VCVXvNmocmNLfNpZfN19hKPAGCCNYXcuoX+dwrRePc2CVRLfev
ZsJNUrOlNr9JRE+yzSnUaAw9ALNo2pJp9zrfVC+HCbDwVqBP8qsPUE3sJq69sfjUNPI0pojS2Av3
Gdw36pgEcJbXmWKBMOZvypMvzTZ8YbRlft0iDWe5EZEmluFA4xjD5iDO9qHZYjTB81olpuB67yVQ
FgUqYRhuy++HdS/5nMncn6+y6+OVrZrtv9vYNqAGbYvl2lbNkwYS4an+VWneIvFhHgM3lrXbnYo/
/hJXYtp3EvNhJVa6ggom0sqADIoHNm2D2fsdYXy438UlrxqSYuXy7WWQUnrLFSS/JTQqmJO3+Zi5
88rBpPeDjJDJDL0222ALskbYorPnT6j4k2ScOZlqDRl6XYp70reNlTBGINpbSSjz5V7oxIhHnOae
b1L4kU/PyLC8KUdg8TkQl68CMP8VlC6QKNmtwYcRY+ZL+QWExP70h1u6ZUxYYEbbc17p5ZmiBYnb
XTc6SQbUL13aBzTgwiVgVVniKtv3HuDK7F0Nzn+iAyPUTesciDCyl/kWYZPUXyYPSoloeAfAFQ8A
mydYAGnZKaw9jF1NAYZiIAWwmbXAsrsUPuWJvd6++lmDdMX/ThEfzWhOH2FVRMvGrVqqqM5GNpen
Qj0iSUpGIyqbMBJEHiBUz26bCvbpcPy9JeHq067+JkDgtQbzI0cLp5G8BwHoM3I0hvUWuzBOqjIp
9d51mSTUoDN0Rf9AIqLr0ZtpsWuI+gwwAMwI3Byi5cCVWvNy4QskIEIDLPh6T76DdLP+rS6SwQMV
moNVUkqgnPtcfLs9aerlCzNrTaLJynZEkDJQZVbTI4s1fnsei/v3U2T+2dJ/Bc2cKy9j2T/hK6wf
rXJupFM6j/2bD4jILH6lgMsko3YjMO/aFWdt53Gtj3kJR+MZuGpTJOkTuJoN3n8PSVbYDviyv0ij
CHVvtyIEnKEMcvX41wQfU10L+gcOLGpYd9NUNh/Jft4zv8xcKyGWhuwOSSIUbm48NlAqCWzxl1nT
IPNIzYhuz5K4vq5SoSew9WsbXd2zCu77kue6UER/57AkYu6eK7OmJlZg4caZJdrZADeDFjyHy/Fy
nJal8rp1QPpQHW8uEahNWu9cHBpSyg+SWlHPU5FFvedbTtqFsH/LQwL6fihXYtOj9KBfBFOJSlAU
3qLeLENJzN9pjghjCn8RrPw5Ig3T+7wcKIY/gxEK7+rkFP/RycBSxs05hQnGPz1I9kzV0yIvot7f
UEofsy6xijom9yr3NB+zlY8Rd3b7/XUdlHAjIsJcPX1p/LFpvcLufPe4VIWNu4s2y+wDR3iFE3ep
WEysEeMgdio3xjwJN0YSBoyaxuetU6gJAKUFMO+EGQ46itqVZLoI7X5K1fjlDd1r3RAiTtTXaxpi
4tGUn1wefld/CLmJxSL2SMWFXSho/JNpQNITJVrXLuJZ1lU2f6qG6snrI6op/sgu2FsAwMTzUwfd
ns/MGHnU46GX3IILoT8lz67jrCmnQfewzaYIaV8Lo/cd79QGRmTUVKcaqLZ8GBBJKv7lVRI5vrjr
83UCsELTGSD0ncN5Pw0yNhUkpm7GlRKgv+dghU6oCWkuHdq2Ku1NhBDYdJO3OE4BLpbuDktQqpPf
YguO+dFzrEqkZ/wBfpFhOqb9JsyKTwbGI0xDo1t3FYfXJeCo561oKXbL7ZRAgV+aLiCylec/ArxW
txI2doRI1sfn64fvpOHe+oB+autrK0t5NA/KRP4XCrjC6YsAz2kUN3MBsTGnrxOXxa7YcbMxqqq2
U1cJC6rRBqmgG6d9LKeKWOrRJBOBXD+kW2zaHFqnfDcYKxPRzl3+FDMiON3f6srY9ntOyXJGDwE2
elYA8xEv8dAJc6eLY6Yjfch2Dn2LMBBX3nQ8eiNQt7ier/9s8dpTwzQu/w9DC/yYy42cDzJbVHo6
PKjDjAEqI99DOE9eA2ZofKrGiI0gw4s4iZEzwZeC5gifwosAk8aPvuJYnS9xuAUo/8AR5X+kPnF7
S27yszl6AA/sVeLdIoYLzJPp9llMuZLwG6Na/ZmRYie9zTepMC9Bs4tZxIN5KaTqf4ndZNAkhJEz
JvSnuHGhuM/qynapQVx4Yu3D5NsZMJl1oPFwkmBz1l2dAlFXupnd0RkRJu69IOm1wqoKF5feUjPJ
oh1Ojrlj7RWjHTeELGdKdjcf4YGWEdScN+W3l/23SLgA17sUP/2aA8X4igk/AWRQGgZ8xHG5zH3V
nXqZkZDK2n0iwHWzxd8FhMg5q1kFYl3jgH5S8Gsuf4E17NlvoJi/2nXWQHGE+/mMm6Q6cANSinTe
6UTiyYeZGR6IDxJbZ3D9BY2pTiiIVmAFUZpuz4PR49jSNQwVGSpg8C2aCjeA0Vw+aI7RzdJg/TDr
mSbSljZOe/qi2jWiozC964RSbTb46da57U2ex5LD5kHIvX2N3quutC0EvnU8LikPlA62JyIyTfwm
gK3HSFXTbWKmyHVtWpcLzHzMg5mHBDJbKo4oeTMGLehl9PUjWLa8hsWX2+wBlyRZz4GwUt4dlOgn
0y+tIcXfN/q/RbSh5dhZaD5Kfx+D5GEpf0vc1BI8EBCrx4bClZDDOjsLyDEY5cQCGtKQGal2K5A/
yv387LC91pwlY3QqoRJ4ADaGNQyg+QYAKVFc89KprQFpMKpQU+eO0cQ1siv82r+le4g+WRu0e+Sm
ahg0QBta6NpP49TpPiHHF15OsDeriU+ON1b+7/lO+yj3DeXEHvY6x/pQ+lHzn9cflvMFQ008jXLn
N4FQCSOtKCgLLeLFCakYwflzUppVmADO+vha4i4FUtpSkNHumoSSCXqmSyGVYfpCr/XRX0FpDlFS
B+yHsZf1o9qZNoBw+4lU+Het2pftjHpWoHu0mXWe/a5TzBvdE+fZ4gQfAnc6aT6zcdKl7TIzMqQ2
mS6+N8Hjw+KaTqiWvsYn5uZk61Fi3Ka4VQtaybYfqXO7emT0Ew5ZHyQub8CHJ9VE942cdw6NfJd9
4XrnXSBf0l/yC7I7yc9PIPrWhb11t8tqAlL1OG4tUNjo4b0j2GVkg7Zp3730AyxpWYMT83UqwQDg
xxL/2R67zDPUOgNxZ3qNi+E0F1oXgd9uZxwoXobsxrCKE3YY/tT9uOg1ijrLigZDT8gP4cQmYK90
Un1yj4tq5r099TJcR5jJhvEJKT+vU8t/qcbTDFpeVf/CTO31RzjEE0KY5U/gUOtuPJf5Uhr6CDj/
mvtMl5v0j0MBWgRHTehdB/zKs/aPGP7YvPWmx46LBt5QRrBGhfYHK2tap2kHtUO9BR1UxBlIkxch
BpV2DP107CyWm3j8P4prMwMwybMtF84bvJ11IU5o0pkmQoui4Qa6bfpgApZvzWbopVPJzSwG1ZDL
J20ehU2O8r/FbTdzNs2Z4ou/4h5cMd+1X+OA2z+MNF4h+x8f23Kg8PtiWHhHeHazQO7wPY1YzBEi
xV06lPe1enrs/SmsLSk204xqelxYRWeledZtAMv9eTxCVoVFj3KYdUFCPCcaXuQK44sJxzusST3M
N3LbzIUcDrWv7SZ/t7yJtdMrD+xfQ1TDb3zZPmU04o0wJBvmd+IbN7YeBi1iu9IAVOVf+Ym52XQB
kBUfC8yw1vq6GgZsRXS1ev4Rwj8u+7gIXdfNdby+nlPsiZPMVCUm2+pcKpjmEDjO5DA+Ba6T87uC
dkLJIPAGGqclqHcxo11OMylNdG00sJSN2Tb1peqdQQWgHaXN+e0b47b0NWyOZE7DlqI0KxO1Bq5x
niYpGbJXchaEaQV17M3XgvxpEy5Wzk38pKWNwij0Al1j0869x7rBsyQB6kKHEtrE+1wIsGDeomCM
SHRugar5CzJ/aRV4YQq1mfKg2M+OA/9PMyvl2pD2hxjQxtDoKUC1pNuZbORW76124IQ5WtbS6mQ4
WKYrUuu1uOgeeOvEOdlqmiEZUFFyZROgkXwKvqgCuevNAClOI5Dmygf1JTxZRIOYkBLqSOhy4wNa
8+3CvHqCAZ5H/qGgl5Jh4nWXohrtakndIWrjH2q3Qur7b/Cz0LIn8jc2YVKWDw94zgCKyXKasbtf
NMRYxk27FLkloPjJYe84cZDN6QFK0DNhJlAvdN7K15FEWSQ25IbRkH1cWH+grZUT0Kt5bdva62c5
0QNeNIU49n68N/5LHBz541Xt6mtG0VPuin3OVdxknsfiqs6OjImhsv4bPelgaSr5mDNvkM5qEUog
HBRRFCt4PTJDtLL86kG9Vms5uBiS0t9dscoAB0RJ9nwoAIpV1iM4PEJBm5B/0N/6eLal/KWsiHYu
GVGh98Yz1KPLuhD2MIGz9GL0gsCmDN+IidwPY9SKHbVpDJR1Aie6O8MPF5lZwaPA7eOXK7R/hlHY
DLRksG1dZ2DJagGsrSQjuyWhOzsLiw9xpamgrZc4BFY7usK5QblrCJhc/fYIqPic6EaTp1g5GwUF
ATa44HtvAHeShsVryiz0AupfLqQ2DL6DssI6ehysr9vvVvrszHkcYhTdG9V8D6zReYyqyeyqsxK+
aPq36sgEXZqDy+Aj35Fo4nlL2Nrly8NgdppqLCe1LvcFB6qcib90R0jgL/2cdIlpHY2bjMQJnjhB
zeCN2YOmqSO0nOmvxpiXbfCGIL8FeZARTHRDMMoHlOpNCN7dqoee/rmljyjMnIKYgQjAaqQa1YB5
rP46GjBTmh1VVYb7E0fmOpZV/8yu5otxV/YfTiUYzNFEP7Otm62tBdrshY9KuUrROdPNZP7bZaDt
y7b42WiNyE8FHDvw1IbagHSjdGGTKpC3nF0LcZ2x+GxJTiFKZ/+DhPdNC2IzUVPAhGDAotqgRli1
h+Et5czFP4uj1iBdN9fmVDDwAhIfSIlpFR/I5vqm2kclhQ5xwcwFDKd2SCkvzJEH2/LI5FEaydaE
pH5P6/jJE2eqqBkgpv7SuWFAnhAUaufrq5tE09obOYXu3+54wZsgwIVMFBWM8rE+Gzrky3C8miCC
QIT+3NTPtcuw7Xw3QPEcK2d5ZtYNeuuwiXHUQ+SY4C0D8C3PY2FRP174p1vx+E3k1jdkO9oAejO+
aPTa9TRSxa/649Q9poyN5joiA1kyPaNu2/WU6ZK20A2ylgbDmJM8Jin3aKOJxyPrXhisLRJgSy1X
Xv2PyaN5Gb1Bn4JuMXiOFzzzsbldfeWFXwgb4TcFJ9U9XO99uMRzdrfxxD1L6fVv5l+h/0ht13Rs
m+e+eCGtdNkA7X99cy24VP86IzMfbnlnRn/OjGvVw6m++2nxAiCqtBuvqoPXu1KKQ+uv6G3Hm0uj
zYOsxli6t2M0hRAFJanSzuyElnzorssdA1HupJzP+e5zd7+7Pul8gA/uxdDDGFLb0ruUUgC+ytcb
2RhANJ2cV1h7SZ2Z5TmYdTC6/qfnLENMLWhTofiupELAL4ypUcIf95XBttiPqE7UAN2bVd1BSrjM
K/ytjMc+e1fJHX3PYBMq53dde5wK4qHPv4utcMLog7TpDJ6Iur7vYYtijomv7VaMrYjKhfBXzGOC
dXRhkOo8HkAewMWT62m0XSOmvMb7sto2VSONofZTnoHyokyyQAj45J9XAFvtbpwYy1Jcg3L6ZHHt
EUlpBInC2AcAB5GOyEx7czW8FQLEd5DYy480uS3QC4H4u6QpUqBF2NruFOm9Dyd2vSxIAscHf7IC
GbNB8ULNOpgI4yuhMijVwxiGwUlWHF6xdXoILneB4oT4TIeVAYI7Qr3nfm7aAEIkO2zOvtwrwczH
+x9sfDIuDcZEdm8vEoWOko5znhvA3wdvcrGisxxnX9g/XVFaK79ve5BtX3Lz9IcOzRIUCekM7Cqd
A254T2q4uF5Rx1ki/HFbush59TojGpMKmFkjwAFBVhi4TxYmSLuDEBno50N0Jc20i5S6CMf/odDy
z2g1pMCM4/1nKg2x/iSEOhoKdoTW/75d7OY60ttXwaIklghwR9EdaiAcqF9ndM7rCn+AG3FiM/xx
m5s5RCtSd5iOWeSm3UEbx6Vos/bmrfthoY7XF4Q4EsZgX7wLlE3V0a92PDHk791VDqP8HzabUQjp
HyrdiDzGfmlG5cI0qI1K51eoCHWanyWn5vIi+tz39YqyVH/ZDDGunweuQA0wgWpk4HdMzNU7d/16
DwyNTmHuzLvZM+LhybyR082AB7rBiReT4YQLX9GUBHEmqrlurnUjT4hxQSH3Byn2Bevz2TWk02Mr
nacBTHgR9dp2ZhYCQSoVMwk2JJk1ZeAQn2nCnUxUoQTzVXx31F0qQpg33AYRYsX2s9HUbcy7WW+N
BTAOfB9RtQhj6W3XU+Ovegq2mSr0w7xG7XMqEXJlnInLljTirSZ306QKyqwBhWDKlRhE0IsCWDN8
F7vZ6qXzhccGtXX/4U1FmMgveomHgqerqJgSAvAN+CzOG++XvEuPy6wQBOrCI48+Z69GC1JYwgaf
8WEV6vt1A4PoxcXZ4TcEGX1R4ADJdysEIlulhvUCbbxqsU4+1q77SsrjyJO3svTop7RW2JAjL/gu
xrq56b79tVcTIV5O1eLaPyU19zFCA2vrFCDFP43DmWUko0apGKamwWKjv+dpJH5XNIGeFRWh8kQw
4DdqE/3gwu6HDKh8NRN5rwjBJ9kF85Mswa3y0ryBjfPw53FGDemt6qeVtBOCvEsRAaP7vlZefcka
yo+8CEG2huzxP8+5P7TCWptT4fP4JVZHsrMh7zsx3jpktmgTBe09foIWeKI7rewP2G+y4vdgSZ5v
OMcN+XERC/bxhnXC87x7gH0Nz2uJOBrcxklJQuW4pIOMuHIvBgmMrcVzLTLVzMS34NBeOTXjnq29
CXJs7RCL7OcVO4I2d0EGWu0yEIBDOfwiscXNYxGlYNCA+VqGbvsQ/+n5Y0GWSmcOL21ttPMBXAkF
1A/FZJpIXtnA347wgsjuCDgMe+ND3u3xNP3kVHMdAZa5IX+6DrUUpRxsMBd/SgF9Zmv6JADD1We1
RRRqQHmYmGl21LpsJKCBJz6fZbnqOHvmpZyvdb5t6I8C2EKfTycc+KsjzSV1xM+jWaFTjL6CcXci
FTxQBL4orXWhK7uh3eO1N3SDuU4wq+n43Xy3YJpwIvhggcRKLoWbVB5zkmuCjRVeFtHTGPc4EIJn
+Z8kfIldd0QlFikOPFbPZJ/iZAicDBMuUN647G66qPp+cV/vAFWLHKlX+KCm06ftaD1c/L9kNTiV
GX+ZLukCCKq/ejlkuCNiWb3Ame2+oYpUno/BiMbiobVMhH7VIBoI4aZmnuRFCNA88Ouk5b1crGAw
hSy/Qa5FHDIWjb+jmr/+88WszfiXQgy2lzs/L5+ZIuoTlpK1jcGGNukU2RZMcaSrLA4FlZGwkB+N
0tEmr94XlGqpHFv6KsYuWg/Wl+GVl/ip2EwJTp1lY1U8Imu2ZW6U9Eb3itu8pZT5uNClZPS+x9j6
uV7zGVQnLc0+cx8bI7mWCIoXedLavT5WmYbndBkQVt/BNmAcp+OS9LHpNmT9eDNqzPpfU4Iwdrls
pNHFvrZ99xeErcfb5uAghJVtIrWF1A00CME3ZhWC5dqqBab7F4myrXSBqNlJBzL6D8apU3MSFNDH
5iI2zuu6VsRY5fXl/0Q3a+AYjW2oQh13u66ubYb/wfr8clJx1Rm9syF/hOjBXs4HZSQIEB/kVJet
B6IGj3Kw6oCN3+uywfSKbDUQsNh7YxtFrJvWx3QHeuDEwG4xr+t1ZyZWKezGt9RVbPkzCby9kGlO
8g65XCTEQMfZ719BG99xfU1vJ6O4nNHx3TK/KJuCEpIa79jOHm+czundYiyky85z/Mk7VpKJDaLz
oP0URy/2J8yEn2hXWOh1sl3iBnVu8IMKbonpFinI1ljI+kwuxHx1aKCGvFUK+drKE4imSoLyV7FB
4eIRzM54LqIvuozUKKYSSioztZwqO/BTljarCuSgb5fDZ3vEFN9mLro/Ud/w7dBGQ9u7XpOUN5LC
NeonkTixXW7/o6lzRdNSbEXhoZ4GgQbq3lv8BvflwdyFbJdaFQR86VF17R6070ikFX07UYrVeA8Q
aamy8VJR5s4dLlCz/TpV9YMtDOrvhaPL9v+p/893MnSg/4Z3YXAKh+xCkD5yyZNWwhqPRw3IqgxZ
2VorhA827mAaiNbemtndj/VB/WFs5/xjb+aELIRSQPuH9JILnrzt397Z066jP1f7xw02+XVedCMP
0ticDulBkPKdZ3la1TnTPm0DOP/ss4SzdlJf/LbXRTzI9hjNEKUnU/pX+Hwi9CCOsVuVbtEDZFdw
uzCmbuKlUFR5HuzDEUkFuTic2dZmH3jljNYyOpBjD4hAEF1iUqVaOXKg8CMV0Lpq/DcjcsseMWR+
s/57DZ71MwjKsNeEm7FUbvdLUN/8wpFte6PqVixqPt0YxW+sFWg7LJsMHGw2i36m+uNVzJ6h3qx4
YIg1lFRiAHc3/AXyKZbqAFysscxQClTRimMhLShonHheMeK1xDqLcoKHV8CfUnfYwX3rdCGBtyE2
ptNcWWvPw9soY0GcxviS7Dyd063y7c2IRvFG77eBnkddrPAkYtGfxnqDGfJ6TzbQkvKGjZn5pl+5
YBbXkYbv9QGkcYxQky0VZSP87uPqkQZohZmyn2/MJcvs28CqwgoiFW5WH5ZWEP5UJCXzXWtaHWie
uPldgQ+NpAw3kz4j6Vk8A3mGyFXHuVqSVzBAksGUSseAjIulQHZnV1xWWBsHoCh60YDELX7j0X53
xqVMJ4NN+KGwXuHpKvhFy8agR7i0sh7/OVys5qHnokbvXe1dvQq0jNQLy61C4bo2ol0W4WlliIAt
vAI4tgKXdv+8WSu3AAxoHX+SyNCi4S6HZI/phVyZfWJQGnbR+9L7tYljm80LBrD/5s36wNrkCy05
zVD9XtlR5D2p570FfZWg90Mx3bYP6UL9TUEkyB+ywpOENswkTFJsW7F8RlW/+gxPdK3c26jg7Iqq
YW4zvm26mGARnu+gFDlBwGziwpAeOzd7pHAJ94nMCvAsDACEC3SbCPd9seMn0Se7XIeQoAB3eFqo
IrUJ2EhvE1VnKNeO7+JOAFdZy6IL6NdNmy9aDSAID4i7TFvSIXvc11zsjVnyMYHeDvw3xSEEjvLq
O+s76t6zuUWswvKyVx4WC2vYUxtZCeVoZfZqxxJFGR3n8hGNnS1o0tDa6hSfffi2GJapZuiqwfa/
MiD2xzcvPL+/QQCgddrF4LlkFuPBa51HubqaWH5VcVeassyrl1nRg+3kFohMPSkfT80FotBkrkKI
nyAJcXzsdBj80eSGaVDMyUuVqXVB8a1GXHYRp6ER9/D6FAOwlSS37ju+PYMhYyHEjS5vxwDjUD6i
xub62MKAi7fNBd6s96O6O4SiT29ZIfNElmH0bXifSKQhfRm6Glp7QytsMiYTq2P6t8GAxc93c87B
QIvmEdQLFoeCZafCu08HEP+c+ecKjCd8LZH8YsEGvCVBzU60Yk1GB+JFhfJeZB+j9mZ/4TfoOa1M
MY7UbSSPVBKZSc2nYQ4z7PcGxcr+QEJmKhoi2znuycU0eRpyYGTmOR5Ft2cgLbToBSB8NH6L7sUx
NHGsUTkPw+tOLl7V2je7OrOCpWzsU0AXpzhJ4ctjwop2vMGwo5+yja8ERIRKrcUNAkPkCBKXkRAl
eQzbqi431Z0rFS0JJ+TZJoUAHKBJysL+M16DcNJxVvuP1LckYvdyMuFplTJDHaj3EpqIN5crojcE
94RQbKPc1RhQPWk9ujDqwYQ+c0Ks6TtxW0o9uHBFlwzhhEVztK+DPrR/PkxkI4Lpb69w2Qjr+4NG
r+tOrjLYk19flECwqeNpt90AG1D2BjFEeBOYD43nc+D7SCCQlKvM2C3baEJjB5Y1NUhp/mrqDOTR
Vi36dmKhhSqGEgB3q3Ln/BJ5DSaGwBVLhhv1Qf4YdKibXH8BRvpNS4lKJdFazcopG3BCfCuWdIwe
iCPG2I4dZpHhquLLDUJOe8OtM44/CDBwiCzsbMazavNAt42zY/uxjFOJZ+sSVmavgYkVNCrqH2KP
WRm1M9cODXzhDK3my6ZvqzkSjawBLOF1ahUlcBsexP358yLf3RfCXL6YG0hvp6Yx9RvVswHFGv32
mKahxRkOdP9ixw9l3ehqnHcGlKA3UMyfbn7aiDR9nXGJPUobE987vbID+b6MRZMtqmjO6UMje4Js
JdG8rOFwbJTykyuIF1KBU4CHZA+WdgOFMjIZzsoGKHC7UVRfnYrT6THa8vJJHGJNCAuWc7Yqm2v6
POA+fI6Sv7VCD+Ol+f0t4/sJrz8YzGYqsauVPGYv/FvdsyDbALzZxDMeXTz7khykzuP28uarK3zH
h1aKU/3ifc2Y1bnUkb0Mjd7bgtquM/JHlq1JET4x12GhT4+gBARjKd3EZDmevicaWl/+0GP90ktA
KykfwQt1hAUAQYKu3kgsa0dwt1sbi5yk4dTKEcLvAqjNJr5nef0SUeBI/gMT6yjEQFUvkB6L3qVs
ZJChzm4vYSZC4jn4b+aZbZ2L45Xv3K1gwmqg+FmifFA4Q/1FoDFdFSYewew+zpDwkvfnAOiXMEv4
FUFLghGgK/iZ9bz0n7fSMp03ZoLKfJaTHyDVyefplcvhKSGe5+Mgc6ScGVo0kfnh3FCD3ThhaT/1
WfYr3xAocjLstizMeaBioOjZ7s7Z+/OQZqn+6GN1nLfi6K/c4TMEEMi4JNQtsyhVSmzTl4cOJNuo
m5fpN6DgsCLV7Ai5ic/ol7fUuWicWuYBdNoDiTr06IsgRlSDXepxWS1DU2XPBjSSYNTwNS05PT3N
JjTJAFvmCQ1kvmFpUnJzlougmcJF29btwi6ZRrSkP1Z0b1iXjBgYPd45IRrUG0bsr2QRkdZ20vuo
rPkva8SMjZ1KmU6VxGjj9Xa/qij5cP5Nex1S6g+/2Jdv16pnmzCR70Qh9xuJfepmxl0Gt69mp30V
ekiPaYWmVjjWpi7w5T5Lyihhz38z16PPJT2mki6x1Ce0wbeOkxWMQ//qmCtBEHxA3+OdPpOwLXNw
3T+Ro0jWH02pZ95kGRkXu/kORdZ73+tkJ9t/uHzD0oBynHK9/xa9XTlOLrW1aGp4uG/FrLhVkEMS
cu4CFpu2RMI5dG7dSOfRGi081Bl1kVOKHLK6EJpf/YDslE85ay1Hx6Wxf9/RPPvVoVdEuUZZs6/m
jsQxDy3MHR7gHLVFUJyMZ0GQmgmlc3rb6b919G30GlXJxOcqnZlNYVhdcmH7enOk0F3J8xK17I0U
xZdBUF89AZRnsl0kAQVyoyM204vozk4AAV+i7nphGpq00pAdbB5gjtKD+32KOooaK89Wszl4dcjr
PQe+78otV5fmuCdPJ8HEwdaIB5WjqMngrmsJNt5+B0b/h6cyZ4Ox5Rqs8zlmciz48K2LReJFZ5Ye
SFcj/QmdJFWKuGaIYELJuIu6Q8cKnlJdNQMX/3qMFNc9SokIpV6I2n3evpKcsWh/YArzRgLPmyoM
y/2yMKotMNNBz6QAnKGiDqF86iiYQO023jWeazdI5qpLcs7dZiat0UXDNNYZ2g5RzdGLxL49IHRS
cnbk5ZUugjC0YmMqHyGZS/7uKVvFM6HXB0AbHcjWecfV/Gu/+Mg4zW/L9/FaDp/iqtyR1LnWJiOk
zjcgDSxPHys4LKewp7EJvLFNRE9v2zCSP9Iw1GG8+KOkbAObnflkJLnLvrhrl+cfmno55ORrNwe7
ssO1tPebyvFxDbA4I1pdLAIJMhmKHw9YIkBqMyCp+GCny1BAWWOMZW13aS40lqC3WN5y24YK2eMe
W/jVzjV92ZsJJ9QUUHJT169Wk3ZXtmgU4sI2KTNevPEmos9xUaYp/NrO/lWC663XKF6JsL1Jl0sa
1+dmSnM8iFUFqu4B+Ha0AABIMQRawcb18uZV8BYo0Zo6YbhJZM3Ht8I67sLea+5NK3nHEyEDtXXu
aWwl8vELSTjnTE0n0LCSYOXQsK7kIxERBKbJRGofKNPhFApo/Pso9kHqiEilyYkO6gHGpAKpqd9r
Z+aQrAvYQUeUb3BaHblHU9ow3K7QnVXq1Uhe0JQZz4Yljq6wWqH28EhzhKDwHUx84HP2rdNy6ukA
4Uj6IjM0K/25W1qM2vuqqvpKADqYqKtF7D2+t2ajtrthTdj49JZLc5ldWjcw6nkXInXSlgzhvpiF
bDor1qZC/5KYXhbutpPUzcQ8xU/oRR0CrSntORXo8M7UYQ325fwXcc+elNRUPXiIQmf/fs1ZrEKF
42sVfeZlyljagGVgF/kLcu31HTZVP3ImokzuJBbTesvumvrEfStoSWxB3Ehjyz2jZ4uo1JtMvfJA
Azd9/aTqvegJi0maMhl9qYNIbVM3RXDdTxIINcvtCBuSXnsHrS6l1Z0STvY8gckgPCuDEXnBls1m
A/jZeSYDwsoV9S6YWpSmIwZp6h72ti/65aS+jgT2q4vU5nANfweSU1XVoAIwHA7VlO4wQ+lEETHA
Vras2QGuFmM+IwDjTHQwVX9CoT3ECArCbcvoBcCsBYwg2/9+ndZon50e6Ze4WMzOySjpkaUUp4km
Bq0s2egLe6V0uz1la3MBLRnsrbZD0NUbv6oazXPFlcmdNbYFoFl4FCDQesHT6zfpJdmzCrQ7UXiR
JkNdncrMcUIFVeafX4Im+nxsv1AZI80NlUkqqjfOF2QS7rPrfL1HgqIttQEAyChK6JbkMHDqlIZK
XOJNu5x4uxzCk0t6nabAItuw82USd4klLsZOGKTgnP0yriFnk7LIYBvGYu3Z3Kyv4yOPAwCKs4RF
9ni06n1H9rhH1assB9Ze7feOBDBir0jubJ7UKLM5PuSgqRcYd7SsBPXimKx+bjx1AjPfYNHTTn/Y
HDW4evrxBfWNH7ALX++9HAG5NDRQMYb2A6nKGV/+g3dKidcC2r//JhPp2/q2AAQ3fkFo5THVKKYg
OB0qsQ0tnu0Rh8ydnjlUj87XJmM3dsFS8qHpPjSIHx7OmCOnU7KX1bPGeV0jtwrp7e/awKSZlPqM
Hc/90aBHZ87Eqqt7Xe/0/LLhnyna3ctdKtEI1M9BJIDv7BLzdrtAz/nez1sDmvr1qJer/PtYUQk7
N4ivmHe2ZlkxEM+XT/+9kJxy6XPWtLRre8roydTjqMI+8RiLn8ylhvtkJqPRRjw1DSUTKeFUfum1
ULoGMNNaU+W/0Rm5RnnE1m4b1D5Vav4wOgQkNn7dvY8molZm9tzMVftlmMcl2wsRNfzXQZ4HCLfW
sUAL3qGuD0bCj9iHpq3l+5CZnRrHfOote2WFcA3a5rF+BtdY2mPsPNf3rdu0TlWleStcsnkY/pWv
1UD80tNmcT/F5KrdtB3ezOeDrOS1j4hZ1e77uozeUEPGvJhFuxEBpa5hh0SmC+Wr7mebzLHMJAlr
k76UDL18K01fn+eq0/qNvT9wz96AORS/SdznUjuE96UWhwYxBNfk+npobHBdOX8B4mP7mdYjj6sG
EDi6vxTsi9ykgDxBJazMYLHJjx2z3UDfkRxzMqBQLy85AWEsYX41fa4fOdjwZ6khPurGy2BtLRbn
JuZ/F5WELXz1nECrKr7WvqkIgOTc2GyMfBHzpBLDEYIfOR0PBOhyy1ge8MZIf7YymgEfpWO05fgz
qOoFRIvv95RsBRgV+SkZx7XW/gokDLXNNZTMRAC0qOr3EpB2jsvmF073rkFYTJGle8qHILqNPFlI
NLjKDPJffz2Du9NPE3Xf1YmZXWpcS76u5DOdn5TJ3JqoTSAv3SGrbL/1xvXWenCsd9IZfUUbif94
Bkpprh4kY+ECvi3B11ktk8b84NADEbhGHdQfmy94p5WfNMK0LgFGCwPzzXI5qJ3C1tVeZk89nfbW
ejRXGgzFwJZFHH3YVQbDfUpsmUW8k0ZQ1GPdt0I3jJJdvCT3XsNwTQhZP+nqrQzTMgb0+9NPoP8k
KvzFmSMHDNq4lFZyB5apzPMbIHmypu2QLPoriATDruX7bTqheavvS/jXWYmqlC9zTKn4ugC0znI2
b1pFj7nubZaEQ2pLuPxPq/7XfDc6U8IYHV3hNecUInCeLEaBNDOBWkW3jYM7SFFQNh8fBVARABNf
+kjIsMAUqVpe27xmRid9GGGtPzmmagptet16yvFVjIOLxyGbz+mhk7U64SM4keS2WkhG+Ldyj/V9
yGWzsNRHUoBAL/2IoA+nNeeb1//eXFO2i5ZEby0DXweaV+UifWU+XPgE63g6MVVjr4zl7fc5nUjB
PQ5QVLyLvdH2JF2FCSuaUe2LP1nn0LUsMYr4xxASZ3d08AAa5hWBXjYSKdtt4PDBBy8045jPY/J/
4EUQd/Saj5Qb/rM6madrYRyA30/yK2e6M1+yhwTeobluO4J/lFW7EMIrdU2uzNH+uqh5gqU0OD5e
xa0DbiMFKovsubtWWR0IhUVePlEXxF+nO2bEiFNpm3U2OUXD5HIrvoCubTPM/wmsaMjx7pMgYPi5
SOSQMc1D79ZY2MOO9z10Zq1xntA6rK8KVS2JTF44ohyADORe14xtGM1G+ebNxh5ZQfW9CVTmbLQl
jDuSmSfIrhqEHL9XHT6IlHcJ2enq1aIhwkS0sQuv8pbWRsNahk4f2KmpJhxOh1Tu3ajpWD6veMTb
lKga8RPnlbg8xPexJmoH1thoa05BY0vnr9uSU5WAyeosFD+7Vb38O7uiCTYSNTY7Utnxoe9tzfcI
IWImIOliPbYiRXf01hyqU5dXs1bIz3Gfzb0iMCPlJrVKp3P2VsAEryp4d7ZKLvtezzm9txJcdy8d
PW2a8vMac/OTA/gb4mN/sy3NjEsU1GrJXBgONFrUL6B1T3c3zLcGMWCtCRWdrU+jqHD8qzBrYwWA
+RcCrCAsGgmUFHqvdOzrFI7SFd6uwDhmlE77/QnAwApuhpaNXHFEJukrmLOKRSRsChqwwo4gqMgM
QAOuuLszSEpp2H1sdjMZFpNKskoAS3TpALLrhkHbZG4K+ruv71mqy+yzLgn04LSh7jvOTopYj0PW
G3xcMIxloeqDe4lMN3UN5kCpMjDkgfgzTOWfG1387lPwMVmJ22TmOjKGUjPENC0g2koJk1xOVY38
Aiu5KwQqyscA//QIbZQPOEKHX9te2oDY2Vne0TwDfgvA4MWJR2+e8CVakJobbJpmUvERd53p8yfH
tKTEQKHlCNa6baFHLSKeRsHee4ZN+GBi8lJupHSs2TYLgGp2h/lWg8E+RXjRd1JeGmHA+PZGeNow
4DDTE1Dn/5vTN8lM1wVQepnhZRvqYvYjlRNG3UdSRh7l2n9ziWHtRVLU5qMTO3N6lobK/ABrYx+e
SAHhmPEPhof1N+fvVUSfGMAV8LXpStmY79F5/Sda8T6rDpkuhFcPCWEmkFEWahyQBTUMb2WPXGwy
HMHe1JY070xlNZSMWa5Iawi1+9w/aYJRGFQZDro/tUwkhgeDUfXR/dEsjaejVF1YTAMrcg9m/qi9
NWrJW380xBBaJSJebPfTnMFQ5nISox83uAVWXqLcKFilaW4bXezQ1qacWPzpzwDVQDo40Do92rFG
lRG5uT4elZDVQ5MyZVmeBFeYlCakDb/VcGOT5PZJhyJUzMFQczW+m+JQGjxMrYCJMaA1N3+GmU7K
WclqEFUVVHaD42Z2MK+fGexZXNFh3FsmBkHxfBL289j0t34R5C4N3y7wxbMFCTsSbT708BejbtA1
GWGBZjXXF6DPYb5JdhQSIgMRe3xomrt8n0LJ3123EgCCuUnbqhQ+QxbrT54tJNpybWI3tsjkZml5
dpfIR9vScoNRsLz02gd3XXkYe7TpBo7ezvCKbePzXtFIXkFInAR1Cklms5lCU3KQ22V/uGDd1eTE
s++U6LpGLTDn35UsUFsib+WCnvyLBmODsDkiDE2CX6hfpoPffoAbN/4FyOylv88RIjZ9gx7VbXPX
TQk8RjEmXn+rjkmOVSLK9h+Jqi7RHsaAJ6PWwJGmcxjn3g4hHzcOeDjB01Uw0WHX07Wkw5WIpd3k
EoiE/dSIHtKZwUOirV3H4qmesYDMU8MS29Es/+oDRxyX1iugRNZIbgU+mjfWS59s5S7Qtn6tGoRa
InlnKLWIOI1meENg8Kp0t6wu0BZDLeY1anhYMyb6bLuIAVenuqewD2pcDKB0n9efclYSsFuTzCGR
xXn7ee+tSTuxqTHkXYbE2w4YWlu4S6jmz3NzPdrACq3JXqNXUbO5vxeQO1yGaYez6WFGsK78weI9
99hM+h4GZjfLCoBimvaKuhbg7LWW0k5ngqm0Rd+WBnSP5+fhA7WqALlhuRUb81+nf9AadAHbIpNw
K7+eGsphJ/n0AaKcSfXPfYlGCd/OT4dHty1dTAM+t1Gd16VBpjP5FAMQI50QJ1ODQGhVil9nXLJB
dgvQj4pUtQ/yygZBs3HUfJTh7AQu1wmJw3/PI3XiVLr/Dciph29vT4MS8XwUH+/6aydQ+RBxgIaq
R1xFL844Oh6DC7QlCvx96G8/wa6nO/s1ytMXBMRKewZI9qrjlUoOXlfjkGA+KabH/AElQj7HRqbR
7hxPL4HDJIOGiUo25TLjPoHC2sCecQLqDYdrW2c70Au8ryNPT0MfVv4pz4u9Ta3bT4Lq2/dvRrW1
fUE0m0l5gqyfxN340ujR2V2pmsmWqOiXwR0ApCd9zckyDypG9ROxFDAVT3UGfJf+IMNIPlnVceG0
+AFWUXcIJ+srxa0eVFJ8zMfQMr/VwHg2sKYfhprNQnba96UUoDPMh4XoAdrbLia9UKfsyZgu97Qs
ez3GsfCteLGLhkNVGzIkuLNmDQ4oNAX1dAbNol07ojqsRP3LX7iboJbOkuMHAw0Uecv7toB70QhG
Rva1nXqvLPaKSXwF88Vmis8EvszZiqwr+q4+f154Y/6nhRzKMIGAYiXuhCmTY3VaVLbBIAGKhd+n
FOsXyZSWom7h2CFEopPP4isEpcaE43Owmj08WT3SP7ZwPAbBaFOTtxaDfW5JZAmJIeImvV2AFuq9
XGe7Tc/00HTmBitZZv4RtYdPZ2fYNmRrzr6RbELCwqnuV02bUknfdhme4/sez5qSTb6j8MiJuYVz
ea7g5dNNHS8ySdS0BM6e+KPFrqpUad46x/0I+dwaGriWNOi+ppP6VSYbveFouRXlm9cMrAbujxj7
mHcREMkNseDSJ/goydP+6Q1n7Ank6dLtAjMoVdB+jppjhhBsfjbyRs2L/xzacjQuYuYiyGRShrut
JQ6lMNI/sm8kcn5H9Y5QYWfSN23d33QX8+iDqPkbOE6XVHSidrJvrvCaruq0S4/snewZk9/Ny69s
6gx2XeVqzHc313vd/Z+vH7iSgyAR5ZOJCw1zIJfOFaycoZR0UQa2y9xZrzk5xcajjXADu0W2IfuD
MBKN6YZbVfdSZ9st0l2A9CtyIBGeBvyM8q220EDG2l3JCefzaUo1cbUqbu44AIIJvuGNBiQc+oI/
HFeghBv3Dwk64CHTlpJfg/9ohIQ3cDOtDKC3q3qTItcYJR8iaWu/0EfYmJ1tds5X+iC7kYmTcMLH
H4QSh7Sy5Jgsmar5PXutiJIwxr/Lt+1n1SAeYbhl7FG+dqdjMsIedXwsKHiuNkSxq7LVHruF2dYW
tNAZL7ThKWuSciC9T1Tw68X3jaW9Ep0tlUSuA1E+EKIOBlrRAeYE9yn73JiWqsKAlfiSneUgiGcb
MGlyloXQfcyCXN3kDlk66FPinY94REsKoWvKvnyehgqrxLgovQPm2pbxD87NGqMK9eIscO3sH+PB
f0wwMEgqeu5uKaN15cjnUR+gTd/r/HdsglF8eJoc9Zh4dL5AemR+0Vw4wEgJuP5n/tCGP/g5U1hV
f71Bq2UTfqgWRMZlQardFMgKnM1CFhl93FBjEZFZn7wsSarTT1jd08m7FoiaOBFXdSYBSILSrfnh
d7jU+gocyk4PbgqbLG+tHeO/fZDVdfC9VXyJw/6xY80l9DtalBcBHuyBAURJ/2czweKyaGq2Uhnh
uaA27ePwXzZSjvel7jAhiCnI5DaNRySYaKQdQaDEE2isfCfidqIIK8cq9ZsDrOVKZwZA9XV0t4iM
V/TXt57M/aSKaK3npwkS2DosDah/xP/6O4SnCvGdEOXgeurVfliMKmpCAV6Cm8uh9O5xmRg/1bz8
DjBVbQ3CnCsnbVr8PBBEY/gAxY03pkv38aq2pGbL2deFIHZtAiB5APHb1pg0ffvpQLJzihgBRtYS
hVnCyKEEKHbWYAqeYGGnpnmMsmxWPX+EbPI4Ll6BnO9srFbv9AtCeiYUnrUq8xfsspgP28o/9kmK
O+NNFxIWM9pUE9uZmpznt6Z0FJPnHxjTxgGmBIwlmvjlLJWtIcCv4WcgvqAJrBWEajhmwSdRuojs
OCIkcjNwdAuyY62bhntOGnROX3bYFX66Dm+vnaeK19/XqIv1NHYoFfdDiAOw6Lucx2JHm4Bw5/5K
CAQb6XatPFvJwM7Wx6cU0CQii4kRjpTLAj/HpRGBiMuyXG/wRN3sIAbEEpWNczDeXeWP1za3rJ+s
0Y41fVoBtrSUn9Bpmm1cJDq5Q7GOwYow9aBfsvht23XO1BSR9e2Sij4u/pzAxWxx77S+32Gw4f0L
qgtbDnO+RranVmTYvfXbEXxuNVEn1XmPiyVAOLrXAB0X21UUa01yRXDt0pG639KgAZZwxCLVh7zz
51EeQqTXzL2s3m4qiJz7Hhe0y1QfXexUhcOtiEkU6EyjeelDPgOR3q+TaWf5OYibIoww88XpQvuU
0Wt+aXCR9tJ7GiEUG8BYKDabfe06wh71o5l7wxIkakP7pjOb3wJMqGXOJKUBt3NAxnunUeM9sBBW
zvo6qGjbqkpi2FE3oj1Zcys8qT8j7heO0eInmx/dRzB/RGsRcHhPcTQZd838JVXaYeJ7264hGu3s
jk8papE852dEhuVSihl/cqVy4OHZAwqkMMqFvvH9WZ7f8zm8Kv+FSTKTLUOgl3bttfS2oCG/CnhQ
58um5p3v/3gh1W5jNxj2kgHyQpdhJNJf2IrKxN34TZ2jDhkL6BNfm4Pt3l3kfinxFRxvM2wJZGDw
nuQY9HNwSsBVwIAeDJKn8zAdh5VYVpLhiF31dilM2DxEZs6XHDQ7c2NxLaLyThfoTOwJ0n4W4p0k
f5Njosmicd8cwVXwiBWC9ct/ie8yQIsQ7VUfcfQAHqlDhG4r/UeZ4c/vAZnI2Ma9nN8xgB1GYEMY
R5OtuFHixRCdsqp0XReHEh1Z/QW9OLLC9F9+7YGJ4oA/Jpn1fWJwg6owSyVkzVV2acTJnRftmgIx
GcoTqzqDtnh+RMsFnDqze1dFsR0iN8P7gEyib/ILI47A2BNN8lIhdYNdBz/HiIGhFiBiu3LmVfSl
lgqdAVU1Iofk9RYbR6HSm9hOlBOnqQtkE9nHXeEDX77pjsjOaZs0I6hq8qzODF+TuD+cGM7Cb8lz
UjY2fXMtSWoJX/u5p+d9iG4kaqsB963vcXD/O/BYCLUmF6Eix2j8dNER71RyHsSvz0+j2vEhRS7k
Wj/IyBxTmUSlUnyenUTnAGk7trivX6jDnKuUMEZMAl+SjwTMRxBOk6CxzkBA8/7NvMO1mYZFSXhF
IV4QWQCUsmSiznDFndZBX+ToSxRAO9FYAF8xPdC2S3b/PKp9nvcbWj4GHIqpzlAklrXb60C61vtk
u7zJbcMgzd0YGtnit/vgO4b9uXQd/uPNBl/6vyoirueZlK5jevnCDZqs4gMBqI/7ObrmDA0TnVJy
nS7+8v1XydnVEFGCrrKUzsrx+/WQLG/zoPTS09cCCEkYTRuDLiEligsCdtuIC8Jlb5EKoF/Tu4fN
eqj2y+rXMM2g3spLLiZeJW3b89O7w2/thJhe7ng8uD06WyOLuRQB5R9KGUouvdOY6BYPez0DzYCo
S7bzHZkEWYvfjVBEvIkrRCOBd0JdbLKAwbqZ8KOxJYR8172/2dH63txgzcYwUXV+1Dl3oQdWTo2s
jaKrW1yD75Vw1N0ee3kXzzKNQeOwrbZ7D7Ryjat9p9t7mhYmtRybtNeaS1sGVrBhfR3mz/cX46iT
826dUG8R1cNZ1vs2jSrlVrGIpvmc+mkKejxlhux2Muy56BBElqGKCBrClKosOdLj4iFeNzah6sts
jELjOeOOJgISExrsx5bufq2N9l86RQCbOCRWlFZoqoQO55lDSBCDmkSyjK5z1mfLyHqGAQuSF9it
rHgiPMIVrNq++OqUWbmzM3XUfbBEfWlNIieXj0W9Pml2+BN+lTylO2M+1y2XKF3PxolRIKJGzmGR
oC6cpFyoadv9EDshVLiEyrj76HPj1XMEdRieC+eQu0mX2+M5brys3ejGaqph8oRdmJKklCJXFo4V
VYv3RfhdvvmqVz6dsUsei1wmUzL/LOB6LAU4c4uDd0TeSqGmoPMxC46S64TfqMw/BxL6xpKK9P4a
ck3zIMY3Y90HTsWOKV2igAc69mk4FO7PZF4SBLRN/6bTfxKT7C/qvcq3o92wZt6opjegm5Qiz/AC
0gk0HHYeq4NAWRWPPFhbzBwKqBA3ZfcczzfroxmCv1e6L0bxxNM9VdhMaqTIj32NH4D9VGCabTyO
CngWufhR4+9eLpcIxlZZEvXXhXJAA2nSuEK4hNZm0JdsPH6QBtbRf3PdxXAsWSpR+uZ+PuycvZwg
TjmSlJX7maDniI8uzlET9JXYVBCRNnQ32c3LKMOw/h9Nmqc5PJqQ2TbWa4V6eu7rUkga7y2kRtMB
Kq8/4cbGINPRbo+x3k613ZSuxuCvTdYG4I7C1HqVd59kdNxwL1yIP2lxNlIT1PTFDqx3WAs1qooW
bze0wsciufWTkllwm6/UZhlCoGmlxdnTdVJHDflHy5iIVPuDQSPfymdz/wEHqbUQQkfIkGmO1wIy
G23UHF4IOd6vjJCe3CZ7r/BEkhggJBo75B/Ozm7aBF7ueGKpZp1WYSNy21UUNq3yms8yUfZRpLbs
+Gi+NyoPvnN4Fx08MQxttNQGNngUYKxNfUtTm26Kwg/MAple9DAGsCiIw0EYYEUDjTIC5+t7Fq0z
Irzr5J0JTunCNdtT1c6ucitxDcgWqzP/VscFTA3zpch4yJjRh27zu1BfRf3CsOd+cqiyr649OuQ9
hPAca+09FKD4uTjzyT/Y/dikC6YRLw5wuoWzZQLREnK918bmsuGuLhFj8sxXW14M5Sc1dFJMdPtQ
6ll/NSUfIm6bCoailXmQK6YuN7KB9k3m1wd8IeD6w9mniig0TgvTqomy/tDyzpiPz/295YfqLvVP
csN13qM/iC3n1Tu+SjokiqXr29z6mKM/WY0ijhb8djQfHHZ/wfQf6kurdq44wN2l6BIpHdk4rRaG
v+mYDwDU5MyICuE68Ovwjlh7YbVKBMv58d1W1UvETZbXBFNhQIvFVJW50TaCyyVOYrGzRqIjDLsL
bLkkGofYTPl8H8SbOgVW8kpUJpTj78FGiM8ThESoq4HJSQXO53kJ7Ow66tpqTnVx5hjGq2g4HyLC
KobBPvxTqxEiv3ODY7Rag05r2OStaUgWuTZ6U/bEbVnGJL7sT4X+lwZ/ake2m3octpTGR/HG+3ET
NPd+klTW4xUpaIuHm2XaitJuF2gqvfy4507WsbypBiEGD7Xvcwa4WPgFEUP87BWabkN/QfB/aF0j
vErQDJpGHWxiulfjJOiUZd52hMyspsCg83STaig0NXwpStCeq0kuMvBPTZV6QFV2ami1AvQzescB
OA3cUFJeWWFFwraJPueNVhuvb7mQ6Xb9UZvShFgfgI6iHWBf8cyO3zwGGq4OP8jL/fh4bjCUPq1Q
B4ZErYigtWQRfGzSu/AfvGXgw/Vf10+g6xyTZd2+RhyPUXi9msUpB8L63mNJmezj1xQmOvX5Zyt6
pKSl/Saol4yg7r1VA51xJIaaVZb5gFZPZgniZRyhvvG4EcE4WP6xCFD17WYNuxNGsGh5xqs/xZdb
Hm1cF4KFhk24oV0T3FVvtEHwWMi0wy047jbccVmyfWDPRrL6Za8PEOeGIDg9fMI3A/4pwZSYe+VE
H7g/3I45Fq3riZNbF/pGnqRXgYArQaQuqGlHlynbKjkTMNw2QjqGfWxHHZKtWNdyMW+Gl8cZrxse
QI4fI9TYXmTvszHbudaC3dO6CvFGEfSRKYKk1VS4k4BbUdECvtDzc5LtnnWgkT37ZrwsniinGtVx
IdzNO+J2xQH0hmRXL5OCXRvs6EnuoaHRW8vEr52KNDJtAQXJ41G8oHq3Ep/wof/EEYOs+c8BxhUA
kR9Z2Q7Sk7Vu/tgbLAXdQQxtOwrAXBvcUASIf8kZP/XLkYGighmIZvCgVIExTX8MQ6mlfLdUZ9AE
tKnlBvdFVCh7yPP7Pc3ExQyjQN35BuU8J3b+Z0lCxE7vH6hBHeLrAgKUHrpX+r2RsPjvDyRnl7qk
7MGUEyEnxmxZ9szMWmRpi2NwxCoQwHlV7mSi0mS/IKXBHoZweArVnMcIZCXTQcQn38GwBj7pScHS
dP9QidZaYtmgAHy2pyINZ6bjsp9cn+39JkQDMcEcbmckNsMMijVnOIenNbahEW7msWXS6GzdFW/g
MK6ynkkHQ2cYRcZbSwe3Qpae8GhLdPbUSlrwN0czcNN0F1+msWr8FBz5dXmQyjUsCE9o/g0/DZth
lc7jLLZHfRgnwfHL8YvPUQoTcTp/ZmEZJew7GLlqROrrQPpW4LlYGz3NdGzwuuGB7Q4Mu0dfDhSB
ajMlE+lWg575FNujzLngsqsINun6CRlaVhXbznk6uEY38dBj2OOCOcxCYqP1gi7IwZvvEAFXBooO
NyUaOUb7gwq55djJ8slWDMB+FFTqbYTCCZSpjdWJDYuKD4957hsN5lY1l5OHyK+9AU/dOCdt78FB
PmojrKFEXp0fLtrX3y/Nvsa65fMwmdO6PRMtnNNUNjGFNRv2pejUyoyU1UVJ+medTTC+KqvGX4SI
dGTu4/HfqE9pqEX8MY8v70OdUr0GvoMPf4Jk521tKa+uPbSx3BD0h82fozt3nY3bnM/sJ78KXCwF
pKalLgLklVYuZg1eHEWKzpvVBQU/K6+D2tqIXw0N1QU09dcGObjUSRLAayWrvqjJJ9PMGYra+1b6
LzaifH+4iVip2ASTN/wl2bXKQ88nUBBTYnB4NqzPXKVUCU3sk4RyHQJ1Gw4FUd9M6DnxMgdwlyLS
eOKG+cElza3E+ofe7zUpvoMv9Or9/CUVU3r9l9STAlBdZs0q8eIruaQMn1lC0LdTaK3Mdlp4znZS
D9vl1U8X1rnavto52bo9P5gClfGWpqYd2gQFCqF1PtAsG6/WspL43OchBt+CpetBKen4GTQnop7C
j9Ck0Rnb2qLjlRbl9gUtWIWZsjEsRgJo+0h/vD6+rCijbEp2hgPBo+IXeJw3KUsYuEp642A3n8zw
h894FMUb/6ubMDDZ2NmSBaBahebfF+5jMmvXgSyyRQr1j6ph/KY9DeXSGtvE45izdGdZNnEpayWI
In/Eea4TQhMGK+wdGOA3K5VftaM/M/LR66BvTnj2rh8CUKnFeUwqRLeC7NQoDpIY1BzrKpsuG/sM
9vQK1oUijmrwu3uDORNHvDF5l7sGkAmRsDj21I/HoI+vhfZ0LciI2C2spRNphOQ6704NFDJ0vknL
0tNN7Jb5s1onwcctWt3U8XcZEKrthZVeycL5ilXo+VcY5KypEJF9EeFtY/vJk4SWxJnxkNwGabLC
6+U8O+e6MnU8kyeOy0OuXy+MkffbcwbkNUfcH2/FdfTOQh2alRZucVKT/ywYnaKnhXgs4REYCtIr
/oEJNwoGleVUS09n0BO93wfROzakAhidbbVw1F0Z2QgUzRg4Puafi3+g5lDeD5Hj0rG5E3jenZ65
Na4BfHL/CMO21N4gwFGuzRnq7qOM+5jnGrJGJaInH8rzBSZh4cZ9xuV7V9Yx/QVfLy/hK3MnAgmp
qnCl9+cBWuLjGZVQe+9jB2SH8UwkpFh3WNIfV35P/uBANlWk3ktEVpT+Ujty/C7WPRRKcZs4AIgP
g1Pp1/cNGE93oeL3XzkUUPwZxjdEGJG9Yvbrc9ghUDzHsqhXEtpeD9zatSxhAlmhSIPTLF4rMLVO
RUv7o4YQWhfGsplB3hyyqP4Jc2+hwiDVD40Cc+ezp4O74/rXlCuBECRHt2WU+MyRX/kk9puV6Og6
76RgkuFiI+noAxd8aKlGTIdUpzjayVU8U0gcxMYpfHYv+5YW+416cm+7mpbpP80mJMq5KG6HqRHE
gbUZw4LvH9M1P8BTBesn5QgU4jancgivYQkY4u3vZwgPRRCxUeZV9lgQdf+FaWbJSZ7/oBdxz3KF
TY2HTGgfqvJ8/qDOisFcYnXQejDeUxxOHXUru9Id8EpTcoKjar1HtlzctY4bHqNY5g4mtKltsKUq
/Ci5gHmQy5RzEG0ks78dKxYT1/q0QbBy+Mz5zLGHpFb4OjciL9+zc/T356txXNRs2gpdsqGLZpGZ
aNGxcQPpf7TW1PqIlzj/2+nB2fUa/s5kujJcZpeiwwLa0xGztEsb/VEQBVuCg4wOpzIjfdxNDHbx
JIHNGv6fiuCtYXtw6v6LTXvXTNmQ6Qqe1xqZZOH9Mi+nktnhCejjy0n6RdwujtmUdUNn3Ak+huKE
flw0v5IyUj43rJuzpyiMEhBaFXF15VogDESrgoOXsjd9qVdE/3NaWYwGTr67M8AZfrM8sU/SrIs2
rqv81QSBYNiQ1gXz8Dm1gcM5sHJ5seMyinie7yZtwk8gpozWb6dIGAP3qrhw0hXD8i+SoFgdrr+f
4qZzlL448Da8Y0ZqKu9D2CAfTOArOvp4aw874c03aM5HV+R1TsAhZVuy9pT2yvpty5KMpdRJi6ea
2SrRAEETThTuSRtv6PPtp7yRnbM4vLognAjyqXFJieLB6SZLUhZuqFmf1Jhp4qv7OEnQ+mzpVVtE
ALaevClWvsVqUGOOKzk5z0x+6cbyyf/r/yX8IvEEiP10MQk/bs7miRwg0zShVQU0M8AqlPs8cBVd
iZ5p/tKD9MIsbwU5voE2R8illVQXX0Yaf9mYOykUR6fZT8xUQJYDcdKFoyL6RB2qrm9Jg/3xu2LD
FgmKGq9uhMH/97HiCZG3NhHPmlAnxeiRvvSdJK5hFVpnfb7TKHxp49fuSVQIXqh/HUsXj/0fPOPD
Cy7LjYhLMjBq05YMTSMtJroqn87N58oQsodbPxj59Xqe22lhqmtuCAXBgocUrvMJBHzEONY23k+u
WFe4wsOL9rkg8JVyy3N/bZbIhgEnow5tcoiiu6bWNQwiEFoNj+ZcW7KoHAGHfBQJbhscprwg6DNb
OhzeHBZxSsXUvoVwM5KtT7jGTOE8pWO56Wo0WWMdjMMVbdrbzYMzAegHUpWeqH1Kt00wwvbMkoZV
c+X5y3DKw3SZV/zcCcJh7zPqh5wzN3BRMRkhhRak2lghiRJ0Z25vKUcq+2DSi29bJU5yk0hoUq/i
M0BDh9woiy2IasWPsYvPuO0V6sybe/vctUIYIPyd/BuuHG0fykTosPYnvHR3Br2fO0boTug5FV6F
f9nHyWQ2VVKXHIq5kO7ZBhzMvb3xja5JcI7TlOxKjVEwO0Fi7bremB56SKxvb8qK1HRX5ntMFcQ9
9pmqqVG9Om6oeUOWiyvk9n5RUQqnaBX3vM7fCHMpDh4ROwDUDLdVly7qPC+E+7Y5VNnPgW4b8Jyy
/LJ3NLeS3N1BGf43B+ojNIyAa4IFtcBGi1UzicMg1ev2Aq679Zv63Q/ySy/AnaChgOZxtIDbqjJn
aIIgmMRpfoULmJZA9VYeeW8FinPbYeYLcFi53IpUtAfbdwoEoy86pN0Sj8WSUVST81unXezzuDCb
6u/cwdmvollFqbMq5mS/vfShLLNluVeWAFyNk7h2t7SqFIcd1MUW1tb0HqjiWll0Ui2dXZIayv0P
sMH12zYyH9auk3co3qaquwj/6icHJaTatBGoo/v4Rwc6/uo8Rpd48P7GEMJzksF9mTI0sFTkrJgE
zEc/MTaVkJ+th6o02XRryrlE8lVbsJiLCHUeSrU+9tGWmdpcQH+x1hZo1I5l9abNyxyja974jgBk
YUgjWW8OkChfIx/u4lQDc9mjVhbGdc1RhL/NjSiodUtPOQHDK5UpBkoT6+LNnOeKS/cQeBVXX6hs
tSrGraGOQVUeURpPzLes6oTXqxKS1SYo/9+qdxw5EBl9dr9QBb+0vMomNb5c/e5BQXE3FcN4rP34
psDMbelXPrIrGlU1n+kQWYgyh1Vktf9pZ+JksJvgvWsWoi1lRFNzjsh6QpNzGqUFrZnGEdDwIqL4
gKKitr5/Vqb1Ifg3jkJVVBzZSHQH0r2VfdG2bhGyyjvJiGoehfi6qApNiVAqVLKCbKQPz5SVWPEt
YsiEPoI+6ZAoZlPcIefEvwrGsZc9/DcWJ5zSawewBaZ5mszGGea6HcrBycsZ9nuLNxOuxq9SK6Ae
kcSIRlCkawS/uOp7p4OUqlHrrF9NO+bFLOznWSNjhN5bWN+UMPxEXnmqkoS4xXeMobf0Vm+c57/q
0ZYKNPC2ghm+QMbILp22x9XJnNmG0N2lNHgzknM/1D26AwHkRTDlWhnfYL0gx0ywAUrfi4xa4sdP
+TLN3TpqHlAigiLXYUiN74ttvqCFEWvyED/zBjx4C45L1DiG9p3wDqp5ZisJ8ZU22GwX2P2CoQJr
sAIVFcnIidOjluNqLpm8kooQ4ZyZJC0aTbIWO7VbTI7vip9f1GDkPhHYidpo11E076CZpRziJ5R8
3rmXcqZFLccl7ycqeJAY7czFSR+0cXBvNf0e3dAINu+Ui5UPseQ/Jm3mKnjdNsukkyUJ3ZUC79eh
QvLXVgu92L9KEH/4R83lyXWqnRB8kiGwNleH5XAa37pKIUw5YaMvj04Ep/S10mKUjmaFR3ni9lLp
ZyvhQlAlVo0trd/J3yiXrLyRG1NdvhDtxY4qNUnCFZ+2c+8eJrSDq8VClrGl3av3qI0FToHBY3SI
+LD8pPsP6lRXdAk11ZsK2ZDaYi8IvhXAKzFHrqwnie/J9Xf0pXGtJ9F4DFRDz5t9dw6w4FNjFH/D
z52pssKjn6clZH+FeZUSkrv01MKzn7NtnxdCCEWp0jcoXzZV07NAD4Ii8JY4YDW918/VPmbsHLgk
iAcOSUWNv7r7FVqV1DOsZZngtRBc1nhT0DgR5PRKT6j6frlBsfMLeruMdBeFO03gRp3OwNiFY+Wo
el4q5ozWGXPOa1UAVMVEZJIOegL7nohlB7xLezZUfL/Hy4iJ04N6fu55J+8/YlkQCPDQs2ofzr2j
4JWoyU7BInr/EbUna75qJgsz/ZHXy1S8/jJLMqLVNvTKjTM63BV4Oz+ghiCa3bEaa8h1ijlPwicf
tCS9s11z5xLZhBaw4A21vnhsnK2ZWXmBi1bXjLAKhQiqEE+8HY+9R00U/QxuHSScmKGG12EeYGUb
TTZ4kK126+zt7VK7Uw8fLi3LCsP3cP7hmysaqWYDzGQDs5YMfqLzvdWWI18qmwDSefebBsnhkp6+
6WagPX8igoHLZkNLT1EiZLYHViEIjrI7K9ybbIcR8WKq39+W9qCQ9mvLFr2sge3+bY5lu0A5MkOy
/q71+096ANiiRWUfNXCnqtO+DUVbj3F21irSJqQnlXZnoYWKoJ56xGUnOLr4wlwH9w+ziCYnm/aj
wgH5FV2YNrwRHuJXYG9VyG+dpR1KTIfEB1hm+FKhNRyblWDiPQA506zuOboHx1gHA7nBLypTGvqL
O8b+Mi6yClL6zN+WLdQX6rCHonrEwSWCVMo6/Uo6lMIVmCkL7yYA8fnUjkPW/bmw+oI2Kk5VEr6b
aywDtlG26ayFPOdyraQu+TSZ2gOnvhXnlEK4z2RM4fTS0xGgWENdhURzeM60n9ZcIo5dyFXxYcBw
7om8JGLVq4KEdGJ8SBICB1MBRNqSAvDCUOw4/GYT0clvZlBRBj/WE07b3vRSxMwc19JLOJrJCjna
Z1UM1NSoXk/k12HVmUffpuWfrEeXHbBGrgkk3G2Gs2z48uIPOcHwP28mr/V2T9GgqqnddEaOyLlC
E7YJK+EsDD1UNYm72C2mLPnukQxFi1V5YlxzrF2SCUTSNBJOvsCqtXLOnkTvzBNMaSStULaTCrVB
OxSJRkQf2/jhj0/zps0nGu8zQbbZiiS7adaZgdWUUy1yaH/or6HLGR58/hu9kvgRnoMFTbMiLaN2
9UZ6mw7A9y/5ePGEaHCZuNUkkENmnd60lz5p88l22ukPU9dC8XG344CPb4PukofK5MBnNQrxy4ob
NkF8Dtx9GJtT2moVH7z8KFa0s1rTafg+LGTnBVM1H/WLvmxQQ867SgTc3X1klkyl7OJVpXa8ulm2
dLjNRwwB6IBmYI04N4697MIpH3UiLk6aAy5GMx1j/rp6qkLlNb2k1hvoD97Vz7d0Pmc4aif2D5xh
ndF+givyA3mRMGU69d0WQCDyzHdlmpHd1/qYykFN/EZIDTezMS9BFLXzZLBL5FYB9LVVW7SJyPCE
mK2H2jlT9HYsP9cG1fpf+zjjlQPnCoSdXDSGyZKFi8RUfE7NXWEjKoxu5tAiSeQFiONVNYGYb3Yo
jXuwMl75FRq8aMqU++Ikoij/sW2px6+KptuzPNhPOvikhgziKo8DHQKxham913UBEqr6iYpuLuWs
mAWJT+DzUYZJsvTHKgcnpKuIigfamtjMkTjRFFJuNz/2lo69FyJYEFjhaYnSZCcW/bJGNIsJR/EP
7ZpAdwbYOM+GhZVZeBMQ4ZdtHNso8G7juNCbBEwUXsmgBGSQQorg64rRyZfJi/xTnpoAMzy43H9j
Fs6JntNWFTkNrflXlW8HUG+tvdkms8VhXxURRCNBI/BQ65YIgHMFjcXWiUrKXGechtp3ayV+l4EE
L+FXBeYyqxi2tx58FwtSuxd21Ue7OHZkksj3enNog0t/ZrtzHHK9rEW9rpeSWo/fBuAx4OboVM+B
Gui12Bi1TH8w3dfybwzTbCWpOjOicX8Dx5CbOck0+Zup2nOb1wQNQOeoZe80pr3kh2HdnQaJiYh7
gqFkv2ccEkYay22zKwnBABCaTsoL8JkvJgPwEJpJduqQAHubvJbKZwEYHoo45bCA4VMT39DLfrW2
jfC1/Ybzp7DuYb8qQfK0BTFd84DaSe/vGXeKAZyCn7OqNce7o6cUjXDnDDrIYXJDACdCwniLoBDp
bfb0bV0kPhTTOoa86qkYuBE5TAzPXsjka+LbsqLDg1AjLqzIHzs8oVC1HqLN278QI46zoAlVZvtA
dpkUyQ+CZD8KjxQze2jDmzxhQKK2ggN3N1FWDf/ORxWUDPi11SMyF/1jRNkfkcmyu2waqdOqQjUe
vLWYeW2+KBEV2LFOHro0J+Hrb7Ux/aN3QtWy/OOVXDUPebKbVaMVHhxY557S8iFud2eOkDFMUXEf
PZuIlo5YK2GvjR4aGYRZVpiVlXJSLy7lhgHnet/czFqzfR/4aTWhJFO8znKWmwfgUOpcG6+1J9HH
xwQBxk/wtBRb86oLhxVYYQtXwtc23hGZwwWws0yyNiMzlH+0UbTOhskKLA0OniNWAlZ/ADwlV2xH
29UTKEn9VC//Z5Na/87hep5sV26TwwRJfxl4jR6dq2nCi1M9DKscrKN9h9meR+cnp+JvCgDHsWzI
Zn7Y+gFTKQ7EmI43AC2H2jMcgP16btQ78S91dnL9AE677lDa1fPooCXtQujChCgZhBk6ydQ7Q+Rg
eI0rltBBy0/bVIEyTc/6uA9VfPrLmBrylLavPqgC41+9a1UhqjxP6IIK1OPpFb6v2X0V5LxFx5xs
/TOOWtLP8MevDzrRnUgEyuNmcK9KO46nK7WT9AqEiUdAK9yW6U60Tmyr3PNHZ6D6fYPOvkrsoBq/
vNRbfu5ise3N8IrLbG/qVj4YZPICanxT5KmIE8rRQpv0aYmuuC4DWq6GiVjhvEGguUCb5KhQfP2t
bwDRv2OVYGshpzvjlV5qaFC1K6wWYJloUKpa4PzwGo+P83xmO9WOouacEBlBiv5snX5kBeLeGYiQ
wHIQhWW3umqfn/A5zM/cspxeeDfQq0nvAHL9ngTu4OZblgCqPPT0ZMzTIVGdVFi9bZEm7hBkQK/7
qcbxOySAF7eXQH7A6y9fnOiCVa9cvDXe/vS7/g1uhkpJXv+c9SGluXeWFQ9UsbGXZ5mx8xvAxJ+h
SlYXWYSPQMRvI51C7fDbcXuJdLtS6O5aPufplKdC8AcjWY5P/zsPriDlWeTsDlrHm8KmnxaVztNu
f6BSAgvdtOzWLQ3kpcpTKdIw8u7gjcibAd+EW/2j5XQnLZUDBCqF0lDtFog3Lm5Xt7brkiB6woVN
oteX8kJ6d5KYlJ15KXl/g1/OAYrBYvy1yA1U9s5PFiTiYnyZtUpXe9fW+EK3D/pKvnvWr5Kk6mZw
omcu21iiYkr3StolABBRUswj65VCCJ49x7w1h9dUgpGUoOSVgstWuH6A+ixTlpWhBK3/KrHHdxNy
5ztZUN7T3JTIXXtrT7d1alZuXkcAdZ05MAFRD48N/5OXNvH4f2oOVkoLQ8cYjFccyg4cUKZCakaI
5nE29rj3wo/Ni5LM8DDS9OE5tuV23aI+qA17/kQVDdGAv1WL0KxRZNy2EgfF/jkn//YBvWF4oCz9
aWZBdY6XePErxMO5z/RTeii76sVZVdz74CBUo2QSL/JAZ9SsgzSq2V4fdElCgrILYznDY0y3+x35
dO11K+QkvYFEEpsZG9ziqzK70F9w9hPT2ls8kHjpiKxMKhskwKRyLjpX+fGjMy4AJmSlKtAPNVVd
LhkNIDM+OrBk+xYCcP2TKA9A2FqHufNq7bKyww2OFSAr3+Sqjg2R6pu0w9JXEqYZU7Z0qV+MqzhT
F83BcyJfBaC5+a1oOY/M3S0uvYASJXCfBwfqDAclVpyvEOx4R/xO1XY5H9Mn5JLSIn7ukIW/ldpX
WkSgAYXUkfAYRTE/Z2TH5w2L3OKVy1B6gjb07WYhfLeCpoxutPDhtMUwvPfk5jONN5a7Q0EVt/j+
j0vzUxa+DXd1LcnWfMZ1YpNuEi8yR/5bjGH/YalfVfNo41vKAVCVHnIE4jAf8GfbhLVZsrmhyzqp
h2bis2+j9ZZNdI7gEiIk9WyCei5v5fSjYph0FxudJK42wxxBXo3Xcr5i538e6tPcVagREDeb537J
p59XL+uuSsyGWoGdWwB/fiJ5OWcjADFrAUKAOzxnoieEYXEuWR7dN+OOQOU9sEK6DWGLAqzIfziG
MbtejBTOwfnxKTqzeS7x8mlt/uPOZLqDXI9t+pl307qBEn3eEQvW8x6u5Kpjm7EyCETiOaKh2TkM
ZUYRnfVKIaE4EsGJBcJyC/Y87PBS3ApUNOBCokSl4Vg5ykmFtQB03dXI2pNs52hGtLO8aKNVhM4l
+nO7wGy9k+yugBK9fuhOFh73tk9PAoEJnPSviaCtR+hwb2zYwK9vU9o3EvjvyIyia+xdADmuptG0
UMnOtzm7OUEvtOB492QzKBsMoQVWrQvEi4CG5b6GfWEMmnicUpyWTsIUlLhGaLjqJBQK1JxykJAQ
CAR7o7tUH67PprC7uiQgGpm1BuyfjhivzH6a6ntvORVCy5eR6le+eTtrZteJ8riqCrTtBSVxRtQm
hScuZDuz7soBhg20NSLTy2raoDEEk2eHn/s2qDByQ5Eyn2Ux4Ce4sFySGIwNKw3dTXfRmzp+rTGI
Pzu/YnMgY2oArGwawlP3x7AhZDWjIzflS2YiZE9kPTHPj65o2KQOUIorZw25kaLXDvfQVjg73gl4
Vm9YoEBxgZFOl2VfH9ANVEYK/npHBR+NxINuscBQIjS6vKrxRvwEaOlHupW1ACVa5/WQ6fL0dVH7
SwD9KIAgq+Z4YNeVgTTdkXope0aFMbVa4Kqe4+vRoIHiHJ9SVbur2n8gqaZ0yaCVnajRBOCMbLUr
1nM2zKq7mGAUrZKdiEq3eKn+SvcD05xPpgkI3TApJ3v5pXQeJTSX/ORRxKIUaI067qz64ZKNoNfQ
8EjHT1injgwCleXGyCD3hVAH+Du/Omt8hy7YQS+iPLyQogspvMNyNGd5KFGOIuBwZ71OKP5PxpwB
EFingpFQiI5J6S2cZIuv/Dk7ql5YVUSVmf+iR7HK7ob1Hx6piHO/Fha3lHImHKKWliW4ftZPqkCs
3hfYzHOmR9KYNbAEhL2w9uq9+T4PMezKDR5f+kScPxG1c2evH2pEFVsJm94wJTrQ/nwcitxRWO1H
L+u3EYU2gr5jMXVtCPeaoq1+2E2FnzeuMTi22VNhGptItHrdGEwU35Xkx3bdGMXl3tTvuoRS5weV
TUH4P+X2lqk6tQKlupkhX9P9RXtnXlxcsgS4lxWufWuw0zwbkieC250uer1iFqydTaCFBGl6M364
Z+boipW0Wryncfh98Xj9gBf9gPk+2wIY9/EtjdSRyhtfXdJDhxz079ahjsGcjwi2aMTjUli4eASS
466eKUp13smG6G8f/O6eL4B1/oQnofWmMyUkZpkuEPPz08B8FNYPDS1mxCwVPj3+YWsuIm9zw6C6
s0noeDn5jDKz339dMIbZew/DuU6evH5x7P1kEl5dfMnw0IV3M9C1DCc2k09nNvR4/lhp7weGxaxJ
xJ9czFCTuVP6j/mUWdHWDsmfozhXJ0hJ1HNEw1KJ1T3Q3l2g6Q2O+svSQATy0J3JNs3CMnUyVbJc
Ui3WR/IOBltDi7QzS8F4mc9XhWs1RHYkRBYT1hATKI2sHWfoZxNkCLaVpf0VWrw5LnSIQl9hlSDD
fqoCfJ/8Ax/Xw83RQaOWs51GHjdLYhZbI1GyOnbXsrgd0SslH5aSsfnkbt4K+BU7kmr7DBs5yLfU
iRuqb+LvZBGuKj7vHvrZh1zLd0URvwnGsOA/aeDQlrj/oyjfYIzaJDMHmY/CUyEuHuAfMNaQirq4
TUI7LvCjtzdOFTXsJJYQNHQ2Gc3T3qYef09z6KEIwRAi87dfhissQU8iV9VbpdBi5uAWu4z8vVuq
ff7tVd//oTh2H6iP0OMS1VqUCpWyz6W57riPZl0GA4q7SMNcCG2hd4nKtDuXVpCBJt6xdEjHjg7G
zi5v8bW1o6GN5K0TzLPAc7OqLhyF50wNZ3Tk8L3n/6i7h19RWiNuBiJBVaApvcyaDPOeFCPkSShL
Gds1F5m1bFCAjnvt/s1xqYZEayMNwjWC4OpxXED3Zkqur8PKnc5ca1mjQqoTyNgk5Q1ASgZX+Ofa
NrRuNY3ORi+IQl94TD0LkpG3cfWTDHm7CCjdQ5XN5CREvNWSi1oE5557WYpLMBTd143YkmTHjCrR
f/Z0vj7rNS+YBJn9ZPScGcDIjMzYtvwB1jL+r6ImK8Fd6h0VyQO9uN4HyIKmaLQ8DbMqCNsa/7W5
19GQ5oUIRj6TajShQtWJdmEystrXlBfzXRn3KEP728N69FXDmAtbj8CsHdhUGPBmEw5t/G8T10Y9
ehYtYQ/2oaucwiImyzwc34sOwq7rHNRwUWDq5jEqtxCf6vueibbnZHxICXPNzARkDYymXvE2GOWx
Vob9yahhRHBLpU1BDi6z6Y5GCFevCi05R5U7Hn/d3kR4sA93MPxPBITwdotmKtv4hhQ1dSmzLejP
YUXpaIvrva8IwdrVYXLR2bUw5GCeqm02R1x+N0Qh21Go9T72q5HVkE4WklQo94rNtl9nesTxqCYh
EYLKsFYEwsa/s3jt1t3WpUX7HULjQ9HErT5+cO3+Fgils2k/pOt05CVihkXyv6aAjmY+emeHDDEG
mvYHGiAMZIoB25lYKH58uUZc+LB0MR+843CfAEr+YoD5OjMiX1XJFzZmj7Iv2UoLXDaB/0Hqov9/
Y/MbeOK4Lmi3+eZ0DKjaNGjMditAnO3shpKchYf1G4HxUt5G90fMdUJixAipdMDIlanL8Wx0dDCJ
0ud+b1D4FYFU2kcX/xWCi4P+l9Q9TQdGcFXAbHlACiaOV2WXiuqIGhH+vmGNXl9my9rV2HFfbjRV
QekFhO+/GECphU/xzwaGggH194L9gX7g+DWRQHXLxLe56/BElPrStMH8fnJpVgfEmHZx5L7QKYLE
sDt2fE3eR1FVHJKC+YlXG4YobPRTrHiGKkJlvpHCBopcrFVPKhfwDhbGbk9/q5u85ADM5rv8XfW6
gxQEoZxx0u0onDHBaF3Q234oVl3mP+tlHI2/wo2Yw8wmg4DHND2+60EhWtbQ/MlNfMBp3oBjY94y
d/3+ZaW+SL2npnapJ1GYbfA1lgvwn6gC4CggIHbqZph5WdEEOmEJy8VPe3HfPe4c1bXIPon0UxMn
TK/yV+WuXO1UPOCck1kKvpyTrwNoHTJwTFVqmawHu7NBgaSSC3UNx88cqaTeIootOh/1ie/2EkFc
uuk2UAHqafQ/WZAzmwO9lkUcpzo2G53CN0H0WdjJ/yGNdWtBM1uP5HgKvLkX6AhxGpAshwDkTgsO
xBYQkQ+iWFlX1hTb6F2YV02wzvL9ZEv+/MI580qZORUPHgTEmNe/lSXmZjxFTkoW/rUII2QaajBT
ChMQPOgwOOthYH+tbaxvdUS6x/SDKzUsRQit0EKr+g9RlCnilI7JYPvbb5NOo0gLhJh7QJxdeHuF
zJZ78wF768U44jKyNCgJP9qy/CxQ45QDj78IAQ4X6OjicHgTi4dIeiPSAqqArs4QOQml9fa6KXUm
xQvVb9xXOhTnJ+BLbTVfT0H8FbZN1s5yHAj2XJ8DICChJP5en0fxlmaj5ubFUdZfWeHx0odvYiP4
kH2q4AVLSgQ4fsqoas2kodzsFTU+iv5MN5tmzGDw4vVjHWykIjr2EtGP4i4VSpJMq6OlQJkCaI//
zCHcR6Dlsu+FnAl6l0dDPVpglVeHHn+wAx+g47M1WwF9nU8il7/q8BFWObiIswBs10+2k9vvVcxh
UCR89ekQesv5darysuMJLWiz6ezw79HcErBIyjQje0TP+ZO7u0R8TMjgaK/LvufWmLlr8H950GmM
UeI1SDM5jnV6e47dkTNhdRSNMxmwqdIfpLgpfaihvJmUMHDe7f/YNTqsFZMotvZBF3NLjg504bGo
mqZcIgM+wLwONZ6mcrURW0j0eI9i6fZ8gWLhCSeUaW0B/nqLY10S9fXh8Vl3DmdFeXj/2OtIeQRE
uUH+ZWBy+sAMO9t+V2/+GGSrt/5v1Wvb6YUtWJ04qHfFRYhF/Mx742xb10ymRcTaT9YmQEX+Ho6j
6SWqf9mPxvHwfvgWNHO30ucKbWCE3GrN6P6JnGjtf5qRsubekDmhCGB9/I8Mi3PERna8JQ9kjQUI
9eCeEgWUGMMMwD8EjKG6fi9TGxJ6BT8laiMFwNH2BHJ6TyBuYinPrTfo9WH+GHt2iEkkRfBLMzWd
MA/QeQVHqCRDCAtaVbNZlvwkdkimouaI50UrdYimaZStL6eXnoLWkqoD/TE5AveYFN7H93FXVlSL
/fWdI5lNJVUclnEokZj209MosoI7egDjY7SeCZk2Vg13ENDoK8pk0Fc2TpBvx1p54QD6T17bODMr
2tufJ++ajQnhl/HVE0h/S1By4/I5ZnMa45jpRKCuAG/v9p+OZZcp2/W2H83zX69tzxc4Nsr4NSV9
d91D8C7nYrMwg4Xvcq9k5HpQlubVm0oS1NLlOlW5bBX1RyhWa27ejScUoFeJj5D1kdMfp5KCqSjS
uPIddNG1hNPSG0viuCi4Th097BLB4rAQpN3HDSlTHCmDdrwkYG094p0giccs/9sdLjLeDbyU8sEy
FuqV0veYXMNGesfvtJOVh28Nw7Y3HWAVtLBVUY+RVX4IWudKa6ZEyHad72KDB3XvXQ7zBv9vyAgC
Fc4Y9UL8vJmfHcoJ1VVPjU2N4rIRQi8gn9AKmxukam49J1b8v4Aok/zfmESv6g86Nauvd+myAQee
zlJtwUHmbpnSL304uuHYgInJspjmf1MpCODnZjTin7tVgAODrnPIj8p8UozJaUyJekbNla1vmKRQ
fizjNR8GRux1qOeIIliSnAy5qaUhJtZBZY0IgTZO79ZsTpXz4t+Nr6B0otOwQ/d8TFxFn23PISpq
FbGAEku389++jvx9EsKYT7EbsjmXBbLOxEL6VjPfMKP+0AU3YeTJpmF1YEylkPtpG4OG4QhiM6o0
BdSDdrPMdhY8lVdW7f5iLd+faxVj+siU2mYYGdFgxy5f1ohhiFTZgLo4Xwmgj7wn74e3XG39bzl5
Q5eF6+ypxU84VpmNyhFqFAUo5x8ReAK4Ey9JLQA9TkLK99o7xcRQUXmQ/SbqNmY4Yv+cvzQOcqUK
Lc5apJBDlnhSC0IMDuSkP52zPbkFG3NPv3AFWxV26c/oS7h+acfWs7M7v73FO44zhlNnju5BtmrZ
IGh/W2CvIvHwCaFamaZ8MffmFZ4WU/h3BXVwPTdW9XlJnopzb0Zs7ayp9G6H626uWjljfx7LZidI
s5MQprs5L1C9InSPNK8EF93snT1uVfEebOckJSy8rp+mkalJaQM61i9QNrDviRZnlSgIyUtSnzEG
F/oeI57RqzCMzMRnuLTz20YhNujvi+NAycGNUw3KK1XyFwFTU8RDurbJxn5WPj5xo6Ps3pQ0+KGa
QAdxhGFeEjlfMQCkMuNEGK8HQ3UhCu98pj2cmaBqNkmSlCsSxkY2FnuZKgLhUOmtjSeKifgsM9NX
Zif8KQJIsAf7xFu5OX2Cx4mio8yrhSYMoEFKUXYWttQDkJHWixybTkKBmrdC8ZarWYou7UMhLuVr
4nhvObZ2g5tQnWkkR8s3ao19pytqytvNuzH9obtIwbnlbUkFNa8mm4tOWzUiIiby1iBarnj76EuQ
OTJhOqrxnPJQgsNDxjoJcednsBEF2ZurZ8EVcnJJT55Of7MQoo7IqfNj2iqEuR2FQJvlARKWcHZR
+HInoUvyE8Bi5AAmgkJqK9QbP3tqfJQahoP5wqpfeoni8pl49b5J4QixiuLwtOK2HsvEUnHkYTex
lyouFDJvSsGwnmt+FB38WeyDjHkoSdbX4o5Oa4lfqhRvBT35emeNL+hn2tYY8zpCatFJihlKGrnV
nnhC3bqMAR4/KPYed28xhGlJskDEeuLHxYl9Vfjn7ywf+SJzVYyWwnkpwGp8PRNHK1nGV0wpZP8U
15ys9v+JH6gNvLfafTAPUQGRhwLhaqLIAvto8GnGUbgNtmqnMGBc0mckAjYBj9w8vKtfxPZcRxeV
lbqrIazmdJYa9/jj/QvkuI4eOLgE/ZkZUQdyzkuLJd/nEfSnftJA1wCuGuwFJo/UkVKdIQQ579YA
GeTKEUv86oJqEi8lHOeZkDTNS1YW0bEmNLE0nCFLilGCaKF96owDBOfp7qoe52y8Vg9aDgKCsNWS
UBMXu16ado+u4YSh0PI2o1UICbQ7303tK0qqzAJXD3iRU7BBb+rvaE7XNMVNTw/ADjjhoAGJ+YSc
YQZVy6TMUeuSDVxcbpHBPdmUS8qPTUwAv0hjftXAAT6kmxuw9vTJbmOHKUHpQYzrFPtLvwR0XZdU
sk0DXzfPBgesQU9vh5Gf3UhmKwy1AEbdoC/iXyGD6bjGCJrl3SomktgR0ykqLRTCrpGLuo4Mse9m
ygw4xxJ4Sg1m+iwaXIucKUSX2WMUdO/mjZ+Th86FBvid+sfH1jxS4W1vsZNj1hLLe/G0GFB5uKO/
ha/gBiNDH9Gp9ZOhISM0/Y4Xj7VU1RjsDFayIjRnNP5kubPq6zA/VXd1T6Ta9ga/A3Tovjb9iQDe
YmMoz5zWGonHDCOqS3TkEN/cj+KlaOh0tG0G8MONnlBNcnfC8gQ0Vrr8CsbD2RhuXrMee1T5SYba
pAasrG/EdPuJjEg60Ys6hrCbQSgQrTawCPeFeZcxSV3RYn4YGE14Rphp8RYBohGgaj5JHPk9Tx/f
bGuyJ7GWUWV2pfKYYZqT+5CWY5EghOCGObcBU+f2OkwFKjLvj/QV3qHcR+UQbIPOmTMoTUKULKDF
7kSjR0bB+Nz6rm8nU8OHTWteupBnNHRy/oO+eJECy1ggfDbXIx6VmxFj7OdzXx4C7DU7M7vg6ukU
qvGf90o5GYynyVIv5GpXS1iSR3Xx9js8mNEr+8X6ihZTv1qu0epdAl8uTwh/vNDp2J3KiKSl62nA
9gFjFTc3TaO4vKoGlLMIQ3z0K/a8NZeGg+rfwd+v44iqrYOM+YcfO7uu3rJgZqtX2GAhntjVGR7O
PFXNwILFow1q0WjhF0b2bnzeYOnZhZwIFuej1OkFU4Xp6hPH7xK0kxz3X77zfamxKHTRveHGrKmW
SsUpu1pjasp6q0QY/1zEoEDdO/oTTf2p3/2mqR653F4c7VFMAjSOs7U6A0YQZt+mqWZJ3P4fIKCd
FnUcIhs0UfEaET7YTYFmbRzC3vCd7s8L9tQ8YSwMA5b4I8iuRKCunP05SdcXveGbfO2wLKri+2Y2
CJwBLUp28xzdI5kffacaHiKWSJKWa4X2+2KE86GIggloSOmtEBHjvFhWAbNUaZxSpcOUneS4EyDq
nOIGGNkyvQLJRDQRQd6E+rlLJoaR0bAO0RciRnb/Mq61pAJyVhJZ1fXzH6xnatar8QIsSP5F8rIx
sMdhtu5Xc5DTtx/F1wCaaPuo3suSBxLSdFhj78TCX3i3DTQUloNZpLEfUb6/OBuwKHl0DgmmTPEX
VFwN/85/eI3Y6GFJkf7StIxRN3C/4N0BVpH9LLttCDvfuuG9Nt9RLulCpmU0/hiJiI7T0amedFeR
fp7v8WZjdS+WYPDm74vi/47SHc00VMd4vmqI6Xs2d0tkhnQnLwdHiCM1kF0rpYCp+0Qhmhyc3cap
49KNCahDmtYK16LNe9hoKyrmAM249VmVVSQMCfXMmeK37kdY5SvoScTjFvRZjs/p0yuZ2Hoha7BO
sCxCITcYVW7RKDO2EVf1YmcIpF4hdxMKmBzSqcbWQYiLt6DC7/tl1mal27tk3zD5wvW7xbM/piBI
Mpih3hCThdeqo+NZpiwKn21S666iCmOrkhIpXruDrGZSgAzxr3RVcS6KK0XDjUabaR8nCUb/H1wW
VNtDenUnooSm2+8kS9dRhSoJPAvaOJcjYVie6Ehhaer9SIxxNUBSPxBUet0F0wx48DuY9bpfNEtO
GkIlJBj3SyQIDBZSVVDe+N+iZzCb6p/DDc0RpAT3GX2BaLsGewMecL+pDg292vr9Ci5hIlIPBpHY
K6wCJ/9QBgv1sJmArJja/6PscxMpvoOaRVelIyypNENWURS+8bs8nakT+zg0aHl6bgMFLnneIuXi
F5tvNwqrfzn5EMD7+G1RGW3VL3OawKrXohgzN/NPlnea8ayku8gxqPkOC9ZC7NGqBwkCQV+WL0zJ
BtCGPfrBXEOTsSSbyPZNT+VlDH/8/40+s68gbhBS7S35Z9AzDUlTjuegROlFV4N9SiBePzC7ONWV
f1T9LuscLRNdAtgUe8gQ637E3+xVspQqzXSpDirNjpfY7rC0Ky9fvXZY6RUPwjYaOD6PGmhHrMZI
p2p85FTzV8cuOQA6TPG6SL08LuM+1rLJxkEMwnF65TaQw5U5hwMg3OY4tn4M0QZXxPaMgbYR9Yzw
zr/uOJESTF01/Yp5df0V93VYrjULtTcLrgFSFOS5nNmh5ii25Bu/vJW0r1FUa0fr7cMIvmcCWPyU
32QGHXtyJYo1fSLdm5vVbPkr9yWU97tjM/waMjyeYnWl92ddY55RgEh2CTQ0aRqm+birxLrwQ1M+
WOl1axFZE8XxoAdzLbYrQJoIsApqBXlR4IA5a7EMucee+ndurePKlDps+2WNSY16mPGNws3jQPS+
oaT9ntqQVbnwaEWV6XnJE9B5qf4UYrrnJNNrBeCb3wkUxpOHKVhY7BNW0s9ttECSTB3rBhMCZxp8
4bo2nYUd8IVpseBJs5wbzXlesWzbjLFrF9SYZlxA8X3z8K1b6FHZmooX7RnQpEuVhq1deicOAvPq
vs5Up3VKIOXQQFhc1wWFGnOtYJHryYBqdIyTt6595/LO8AIMNCLH3+RhX3jIfjJsjRvxKY8wb9Se
b4DWOY4sHRMXAzaxREgRTUUPdfToc9DVs9AbAGF1yF8yuYhPJ7TXVHSo40JmgpAEX6Kr2SRrhhzc
fD9fP/Abgm73d/7UpdfRsFJt4nKOky18Qxy1lR5tjQ3hAfaLSNNhIZ1JEegh4tShVIyEtWTVsRY1
7dxemFm9lEel+5pHzipBwu7TdGvVM3SfJrCMt1rrwGkAxmRnQOk2SG3eo/4KElio3LZWzW05Wa5i
JiB8QiLSkIEaDRaKbKZffeyOsI3a0UhrIedtvuk+XX1Ojrn2+oFNPBe0Ap6LdR+R/mjZyy6/Ugaq
8kq8CVLlfEpHmW8CIIKrPTYd0IbkU6lgDBmAcZOSENkLbiKlVqU2CRHS+OBwsenraV1CzUl/4HyQ
ap4huimzP6Qp4lsdXGPtIsH11qt0XdZ/1NJ7BfTAUjIm58zWzaDIkFnqtYmzJdua5Ka/joIB6nOS
Xy2hk2zl+WLxmqeb00eCS23V1v4A2vrjsnTug39u3orqnRw8ABig7taeb7FDMypobp/2XL5b8eCq
/lPdAJDpcUnZYp4E76Exw47QGkpwCwLj058RhiMbkc5g8yHS5tOFWULX0Uu/cifp0K93/oW7F+RE
owLkSqeUH/HRIzvEW1b1vEC9dKdF6b0Se1wN25ibAdlBes2KMqLbJS1Ik5XAmyUqSrLa6rajpPxk
YRVzDxpJkrswQb++v8Viy847gGdHDlqpnoU7ND1hd0j9O3JDO8NKZpo7ALUIUyT6SW0mIX/Y298x
hMfx8TxtCB/NbNrNOe95KfzCU+4Yblvxv6OUolilMUPd4RMi/EPtNKO3+gTQyGn0QrMe2QJ/cNYR
hbMmTRZ/q0eUu4kRNjorRf8k9VRMtW9uQLAyVHGez/fGi6iPOmRvyFkQ/eVaAt+wBe166ErtWUei
hAhyLajXxE+mlWSvdJRP0xgsk7INij5S9qz3IGX0QlMgUEw3urSkZA2lig3H6JOklocr7FuCH6gs
+/hg6ahk2iuPnuGtdb2baOlNirksxHOc+eLlo9aX6ptGOFJVqrThn3Ld4qxM9nFz4j2g0sWF5PMD
Lhx2WG3Rprb8yOOczSsHrKxOAir5ADLXDC9n3/zSoATVlvg9Vl7UXSizSye/+gCLdhi8mqUsbfUG
L8hJxeLdhjVlX0OEbhEuKjijU8rIYax3V9+T5QdUSGxU5Ec2Zj61CbKZ+vbcJGdtwZ3KzFbJv8AB
ggD6XWEDSG+FosgUQkglkicNOD7ufbh/2XIQjkHeX3Nyur+oTmlPDphiPswm8L7L8/+z9jpWVW45
+0hEbXb43yZaTyGFW1oXeROyCLiANopqpNKTvt2GAumyXNhzZROQ7843T1hFZoMVuGnSkyIjSVFI
qKMtLyUftYNzoAm8+m8bHxbdpaWcTQuAUeVPClcQs+NmoLMia5mxl1MZ0lg58ccomjoHAnSEI/Jy
XDKdFWzdorrhqwa23WlSt6UbQb2+tsBl/uIGYekVPww3MUCPEI/o0KCdwfYq+uEN7jLUjJJ02h9b
V5KJwJwOi9goK4aU+F4g22ehpbJKeXXZgDtVRMLo/vREsHVUpJRx5Nz1rp3UoOSnHKYPVAEret0k
iOCkroYC/k9NuyKZBC1Ga3CO2Jt5c+uCwb0Nm0uTO0yL3L0jmX6gQzV38D7cSHlbqv/veZ9cxvk3
fxJ0B1y8WRKRBVHu40Z/OuIALRKJQYND4q+Ebh2w1F6zlkMHiPkhnC/IBxw2nzU1w2AWJf6vXx5D
0Ou2+NCYv49WqYJCcA5ioZ8qkyG4kT1mMm22Y8eGzrzwSldAm5o2I+DiIZX2nO2n2Vej9N2+pDeM
lwqpbKfOuihsXlSLHyt2ZqmJ8d4zl6igGZialBD0FVqQcDpdJGKtO7W50rN033oFgZ1axausZMEJ
aCUXI+3KoEG0MTAdobn/IRm3gzFv8cZtc4OayAJzDj6Z5gXOOP5vcR0Kux/N+iJhTo8bnwGHdh8Q
kZYAXd6FI08KzgyMILihIHO0FaMvcON2TcPafkBolL5vVwpzkrHiiJIFMR/xZ+XN8REbPzlzsThF
wgRDY8GAHN2tLs0yoOzoRVlXaUW4FZTbrp8lEbJ4Rbgth//MlM5I/a6tG1pzmqCK76aIuHJ0MFkz
Pmz9YYKWIuy6XgDESZx0KvUayjY/yI1JJ+A/D26PP629zK3YucFBdvV/4tbVdSzvRF54J55SGpjl
bjSkjiKzuefRewyAZI51VBc2ZHcNODxatEytILjGLvVIqCpipojyMalN3biKuU5cSadiyrziLKWo
EOoP23iIF3pqR4ygjt6T2TnjagXL5lJ2DP8NfzemknTwfXOMIh0tAhcTio631vLPbtFkMqwEmtYb
466PhoO7+FeqoE9P2lN1HnzblfFx7B23F4zweyDDCxQxR5+AIjqjN7uQvDjy+gfKQL5CIkjrr5HW
a8my9hNq05nkYc5qNYalIievPhs+V9Zlj1bp6/AKm49NHpU3Hcbs5WVjjJ3DNacEF6SJ2QRJbEiH
WNxqYW7Bgk1u4/2BfMwkVt2kuKMKOZeXUWnOi/CjSUc60pSCWWpPdgFqE9AitvBfkL5hSelzxBNW
e52EhA33pUj1YhWd5LY8N5RN5mZIWvF8AJ+DQd0RGMz+qEjKelEejuMVvfk1KIpwivc1kDoaWd0Q
BQtUCa6oxLbvshzJP+ipXQwLMVK3GEilfPAIzqrswZL0OFmo5AF3uJHIjxXmGTFOouUXfdhSlu/w
9fXx+ixQex+NkblZSnn2baVWySaaqjmB+33tqoKcc/oNRlXxvHXdvsZcMzYjWLR168miXaC2kSOs
Hp5UXTADdGxnZeW9/a15S1zEG6CCxi7Jn+LM5TpcybOvDqzGT9sbQVc1hIHc8t5D1pW3ZR/HV+04
oKGYfBfW99OJEDHr22P7lIj7lxzGpnBl2Ifex1zgwqi46p4nrABNpKxljntC6QYqTv8R/PLmcz3v
+wqNeWA/WITxHMV0g0eS3txrxxuojh0oNRTeznpj5EYP1H4pblJ2rZ61UjRLRuif4mDil7NDJtO8
y2iZDHGEaFysWx0BIljSj7cUP1GJOoe/evdJnaEQw4rgY3ImpDU34gHW//WykITOx1FvmAL/DPx0
4mky6BoKQkeImbYer6p4j9nFMFPUruKKbnyng0isQC9e+SRkAi93zJwkMUMQY4WHtAMavTlID8pi
OgNCy9CaEMeRuh66SD1FBEF362OyNdgkuHEXHrfasqJ1fY011gpShZNGgDxd97Ghbj6IlzLOyW1z
UIj+G5lFKZrDMDeOYUsB58EyacZtpAoidP47L7hZHNQ/99fQMEiB6hl6QrkSvd1MdcQI3RToWr5q
oPTBxvGte6ewROg5pSNBC9vlvfuO++dDJgpU61/HSU9yC1xFsMZPgO4m3cL1Z4/FgzFBWs0zWcI3
W/JToFZav/Zk3p/9D0dkX6YlD7UZnheSaisbhlabSc9aYYFAq0dSNs9InXqoAUvXYGsDlpGr1c42
qEDSLj/jo496iYDofFfefPQWJLwqjPu7eVVcI4GdHgNE1HEuJ9KW8r7kNp9IOXuGSJ/j2TCByC2o
WvdqypN1ioxR51gXGf4fAF1vI3Lvef86a7+nabHPkAXkZFswN1g6+0ZmKvOsg3NSJhsC18WASVFX
0ztCAZPbs56XNAILOJAl2nhn1bsxAMVqgTmjjpHN8Ci/vSIKWO/fIK4f5n3heifTScGY1RKHV547
s92K1VI7XVR/Hg3e8x6yAU8/PwQt3ALMnM6aSahnaWjNipBkbH/ZNtPlIMMgYf2AFUNZzRuzTG7d
RCXE1RP+5isX47/mzv8UjREQR3+KieArsUARf1Wf2ICh914TZPGcFcQ6vBYkJU1Dc6qh6sqVKA4u
4gep3viW0W67f6XnlSWMaPTZdpuxCdLiKCbGy3xULECEAX3vf7w6JUFoi0Qt8o7VuoN3id51AQJK
RpZM5KuMTMu/GpMZm4d39VWMZfJlh9ZypIfIiAbUgbwxP6cSE/hs43QHp3w+uqMt9CDZ0UsNgQFe
OOp8fMG3ySEDTZd8l8fe96Q95SGMQR/ce9oU/NbQ/XHCOPVDwfIOaw4nfTUhqHn5o2RqMSMUFe4T
5D4aXPh31cvtufWVcHOINyqRwdgYqE/qj2/UZw/I0J7awLHRS90Jwd7WshK9wuS/HHgKxM3Lzh7m
1vCxD5S7w32dww3q+HvZD9UrQLxacqmj3cLVh5IYDjyc3q/WlkjWcy7h/g7WewwvCIFxGZcvML4E
f4l3EZrji418rDtTO+Bx0t6F6cCBCgAEIYgZaSif+I3rRiOXUfEr4f9niAHR6SddjelBdIaHQx6H
0q2UWfFAUooOHdbTDLKlN00dvhlRAji4yiJDS1oVrfqj9eM8oWq23RpOGaSLHtWjXdiiv0E95cLX
I5dlammp5Wp7V40nyDA/e4kNYwudk+RZXb1Tac0GCM1s3ItXlbPbWJNkoSFyg8zwOetg008sIAPs
jTjDOhh1GdRphk2xjr/ZZcNMiee3Bek9rNy6cC3X1OlLf+v5OrAl4GxDT/XOUKpTZaWObCLjoYo9
KZ4YUtrsO0fOSxWyqkDsO2Kum5uikBNCHtCOey2te6vdm3MfNsM8vBdYQREak4vGAOmKvlOP8R58
ksI2VnwshPrV/dG0fVtjo1dJ8dG++qqtHIXhk+G8BxnPYnmEcu4ge4ZpMOf3L5yZaJMMgyMsLou/
r6m4Pw9qLrIMeJ1R7FxTyCceYa5viHRGrDxU1Pscve1IumPPla8PFaLGrqFxv4hV8Nn17PU7OReK
TMvgvnV3N4cYIkZg8AirBUpP+uyyJV6TwZpG6pakB3ry5ie+kY0hw6T/fugVRZInVrrq95Il2DB1
Ic1I0wMiYpZZR0mt7+XNoYsZnjnoEHVlD91iOrhzw7TrXq+jpYyeKGIbQdD50SXYD/mxzmEd1LAp
orFEiCYHA3EF9rCntaZSL1RRxmk8ZTYKk8WQmxoV90kmFWzY8eO24Sswcnax/9de2T638LlTZiFg
EDs+95L4BWlW7dxsB39CDxJUR0yf7bT3TQ9GiJIo8IX6LIVD6poE0HcF5SU891kLWC8xCmuskS+L
pCEzZ6GdWQ36HXgKMId07rDqemvMwKGANloTxuMWIXErGr+UYcGgNsruzMbJNJh9afdN4YfWqVWS
6s7gwebIRf6iu73hydNzZkn8SdjTUmgsIXtjEhcJskboFkNm/UxiLARoqM59gRvqqGvZfYBPWTYY
4Oxq8EdLGHbq6raCanQwiQVhlvdmchgI/2q5tCYkHDNfzOAbxGKqNlhewzrtxemYhyufdIl+DMgZ
6yJMeS3+T6Bg94Rwu55Fs27BBBU/uSOeflGAaOiRO+vdrIXlMC0wJK7ZdI8wPSNdi8ZAfwFgdM9e
C7A6yxYZ7S/+HG82aup/GXloaS+Tf309AcZqAh+CC8d6oJw1i1YkaZkce4lWhN5ZzucK3t7jSbnX
pHjDinCHdImoVz52zvJlZGg8v6ZpP3zcETueV/iSD4iucU6bjM2qi1AV/OadWBKVRrbg0KT1LRca
Ad0GTuF70xVZ0T12OrAyGwc8L3/fv8Wr3VHA1wFlTcPgen5L/JBggK0JFuCzD60rOOcLMlIBcd8w
RMICApQev/QY8p6xnbQw+tj8mFVRBWNU7y1ao78DDrAVJJhmIiBx90985fJvfgy33Bth6xvNuouY
4EWN9AsEEKYRLOxHPVcXBINKYcEq2zoS3Ghdr7ksNVeP5SntuK6508lSRlcabwXqXpQ7sNzwDGPj
odPKIRFncxIlwKtCdIN18ct07ZEwGrc+urae9CqNg0UFY2rpK9PCZQ2blgBHJOuHlKeEN6PLp0IE
jlPKnMZlhJS/VwRP4UfZBDMgEolWUROZUEopj5rA+eNpH+MKeQ+2PMvTa1tjqtlXK70sfIJK7UI2
niQsjJhgTzfEDe2Dk9gpMl2ZD3qsiSAbFtFukkzMqtu1yAxA8+jHLNdtNb5u91BMtlI3KGT1U0VA
wDTwNYJaLr2m0nrckDs6uAGRqQxYAmAsq8kxPuGHci7h6ZWmY2Hyzzfw5e4Rb7u2yCY+xSFvQ+Ls
5ATNJqIVfYwaHuhzf/KOwuJ8H9ybxtiuzyMlAe+ZrDzRX6UUp9DyN1zjuEVH4SSlTHbJteH2iTBR
igMb//DxBcgvTtj/ongF4BWsEsDm9AwY+qjjbPb+sKGIMpyN09koBEwWBG9zaxVBdjbs9VrZ6Wuy
jS7HkNnewEFFBELf6MXIHJ0AJCWmtEufaa7D0tF8VTg99TL2beo+EofXU5Cj9POb7CCu69s7dWlU
eK9cUCbfzqfyineygCBCaBnjQQbN+K+FtN/6ien6C9RcvYS/zT28t0mgrOqq9R+lpkDc96bEHk2R
2TWj0/i2SqMur7KkJ9IXcyxybypEqG/855ZC+Bbj/hrpbPCXuSbk6KOYXcct2JSQ8883w/CzkNzC
qVua6hrZtPqlCUNbNzVUQLSJyEdXUFSonvdgNOYVnuGbGE5RK1/ovAds4pFPl8sVIqNDEZhcwrUQ
Y5uEkX099Ac5jPihrLbinE/QTeHQmQDps1JTlgve6BLWJHDTcO7M++sTY1ad545iX9CHriprrtm6
F8H1+cIyeusUUm9LLLvCo/KU6X85tacyHNG5VZAoA0KBLbYoNZaXY33sZqJKZwFlWcMKofUqDm/a
+sFTowzNK2ZtIwZfEgEp8o6D1Xo8K9Vt6HdGH4UKLvv9s297uXHap1lHGWaT87ZIEs2Vrqxh2Gs1
mqltpjD+2XqKkIy56DfKOD33BR7RHU1gtqW3KZ2rDMpQHY6FlYzFdYVt9lHcG4Otjn/4DE+O5AnI
QMnBXSDqL1yTDelfSYMZKMEFAT+vE4PNBjweYljXKKkOJU/vL9ZYbg+RNQnRFg0ppTj8kle/SUkU
ybeCYkQHXfjq6rblIYQiegfrhgTTizmAtmkqgpLtIaBdWbL+/xKvAhDd6I4TsYATGUgXE3XIQDUR
sWyTaP+LA5XIacoDXzZQ2C4YMyXmtNbRRD25sbjEZvuwHgBFYqtEAuVskrDI5yPd5jMEYQM8MqAM
vAKBPMMRKcWrd1iQGkpNRbfv0r4ZNEbSYGAZ3DXhaEYQnfDeNXRDF+cffjkYN7NCXYTh41PjKDxQ
IqZQpQHySMoKyo7QvNeXQalZV9tnvUgcZL0rOcaNIPOYsqqcKDn0hk8MnfBNOPFti7ImU/qP/Mjn
6N4+H6OwWRPGoinVYzygUWfMzq90hyEee0z7VR9ELegeRGcwmR4VOJQVHEbPkNIfmdVGO5FwV53z
KpHSr6BqOdn3Je7GkgraqUIiD8cx/YUbR+U+5LjMOJhU9BiYnzmbXQKqOLsn+btiGdUm9SiPki0r
vM3d9/qsYArpswMdFZEX5ZviOfKnwBoIhTTTLZJaKPxpZYoyCprOsXyMGbT6iud8Yroj6brEGyvd
eYtQUxJfgyiwbR2x0axgw9mB6HxQW+wsnCl7Mr4VaIPa75GF/gsX06e1KXfJmXZoDLXtudqIYWsr
S412sP8JuO1wSm7UC1b0kE3KbRYUn993+d9uK9cgSCUdlqiT3TCCfqpl3yLy8jheA+5gUddoy2vC
lckmrMzwA+fNTq5/t//YhmOcjuLXEuJtVsrSRH53Y4nzQBRlmBT9xy/l/H0PP0e17vwvTu1AhjbB
FU0Er8uZBF/t/5Vztaxf3DtYclng5hZv1mkgkUtqUp0ttgDHUy/fjK+OVov+hP4OkDqBGC5MVlNh
HeJfdO5PXbMPluibTrWJpVPbk93uzc6Kvq3VsriQQJfsX8Quqmm8cHOnd+/vwEXNxJx9JxSVxrDJ
Xh53TKt66BBLUAdmCxnyHRpZMKnj2JnnbPhHJmbWNVhHgjmbb660D5CZkspZoXOhiUzwUEgkwwWX
aO3wUHSfcwvLKgoXC0cLqfFWc7xFFIzMQ7s8+hZj5XFJKcNEdNy7hMAIYcr+DISQcOByvr1l708M
/w/xSV1eFNnLM1UVbOet6DQlgSQRxa/GtSAgElpdzJcgsHpIosUIwBtiy3c4lEx74NmIgUhyhWNV
1x91njZZ5qADY+4lIfM/CzDadGieNFaWkNGBsCrHsBxpm1G+Kts3O+tYv0vQZlCgqTRtYWvdN6ai
JP4eiIaj8OY5zbYEdd5P6oo5zjAbDx09j3rLioRLUwKSxOyzD4F92R9XT1/YN54Y7ny6c1HGhjMQ
Qr0HRZLygFIfp/+YaQ48cmu9GFPLjOmISNHHZWsWDMIR6Cjrkn8i8vDl+qF09cbb7M/8U2NGsmzB
Na4/VbUniTA1+y1kHk3YsRO8p2emIgwY45sij3LMT/DAq4HsCtk1rbSNbKwrKued8r6AIznU8B7Q
60SMcSkmMFgPGxeK15VTtLk0h3W54Hp8eDQUSc0CTa5UoJ3Qklbg3ccl+Q6e0t48krlcdqzBHmu1
ZeS8i+NL8fFj4uZlZ1M33Ho6nBfigRZdzNM2657jwh8CFmjkq9Oml4ijKYVWyg0jDEMIW11lm+rQ
xYBwNIv932MQHh6vLFyLdvgzZxWKl0YS2oebF6mYJxMxEPDkZN3U3Izm2erMfGNHHC9b/in3DGSB
GDNOAcAVJtbMI8AWb1OiOB/qyMKluzSmQnIVQ6HZJNPFY2uaEEo9GmKnBasAm4JiX6j1wptRCsGY
K3TPymqmA1BjEQzopk9uY2b7VClD6krF6UPiCeOY+MevX+txGsFYZjmvEftZreRX0FJ6kwJqg/dp
ipQJqMBBab4wHKld2eLFElZvwpS3c8fv8t+vk4pzAf5A1qRhrKzmRGt28o1811WIMeWevZ66snU1
QxNBXxZQKA6/QoDIuQ9u7+SgaTR1kANivCy/+OeItg5SR5VmUwfczZh5yQSa2PCqb8Qf/5MhrSdt
9GEtYM2tBcuI/2yyPC/CH8BgV+7iaAQTD7It1gJqyB6yhdP/McSb9CuGtZ8zQQsYTCoTsM7tmWn4
mvWizxx468AY2DiPVuRyPtuM4TznaNdjb2cuZkJxtfN+oMDdBbVBKx218+Bb2nQ8tHc5/cPcMVl6
mx0slXIuaC4zgOmNd1K4PaJ1z9baZRfo+bwwlY6x+r1uQnWluPLs+K/Z5+e64WT6c++CgO1iQqJV
qIEulQPOGkvbqWetV22/nGVZWSjixgurkgjDYDu4sLg1tSngayXjT/olZeh/7KRzzwMIZQaR8x/n
Az3FP5aA3vurAfRRZnO0cgbfEA6JQvbHe2pvOoCuDsh+I7XDBcbzjhbm3iN+vN+GwW9eVDnw0RzX
ziac/OpQyLFVOKsqVQW4a9imElntYxhVHAHsCaSStsMoQZadCr/kxLtTtU0Ni+Xn2W7UGvkcwUAo
vdzidNSSuXF2177jnhSbTeJ+8Eqo+B/2sUWuAXnn20SVK4tIfTIA3tSo8rjXaYk8JVQ2WREIh4MQ
YKvEdEYTT61qLPO6o/LsjD37aKZKWXRkHkmqGAEfx0kUFXSKe2oKGRXFqh9o7eMMcOoqzSrbXGT1
AKdCCO3Hs9II+kJDSnqjKBNL9sFulN9biA02QTI70t7rKT0JK5qWt/J3Jzmvt7BjzBjbuBupFkuV
2g3RtwJM7CvjQaNLek+L8ENfTGnzhwS/gvCAacKF9B0TM/Oul6b60I38pUdF7fKZXO3TDlQjeF0d
HUurBTkLcXmyTrt0tyGGnGZkqbYN6zo/BNkX6t0sU9xB0mo3sedvHjU/auJz/kL6p4kGXgJXeuGW
5yu0znihduiE+J3O1xkn5hQ2YwlBhXFlScxU7OhN7H+gheK4ArAjMwTNrLKEC8RgGMSpoEcuLKRF
4MZQnyljiaGz93iE6R9ZC4l0HIsj9eA13wK0LhsgU9xdpjBUTbAELTDVjvZD7Q5VGWabZXELMF87
N4OwgirRJ8WPZ/MzDdA/hhNo+SXXFlXuRJC1PCsuPRHySycZry6nnVRMUOxxbsEkQmGo5b5Y7Wfk
hNXP9iUMaOhVU/R8/PPwtobaTUabYNeyK2eM6zn9hoZan2gd673oDq8JiKqmutTPiEi4ClMrLMX7
vcMNK6vvigAHq8XYy54U+OzBW55LpO73Ml72ylkOtv2U/nYmC1q5Vo/BKZ6m8HiWppkq+Ra1VWnf
ec9FxLFiAV26wE4itvQ8vv98ipMdnsrWi6ZOLjDh6cngMEwfWDrdppRyAhyQhJc/JxLAmpzWPSZj
OZP3Uol6BL9qrTV/ITNNkZAp3RfKAu9VBpqDQMGJEuHmgKDc2EFcbxBczVur2uLsSj3wmKK5Km6Y
0meZJ7rle4cMUxB5WGCGzqWZHEKEQpaaO2Z66/9JkSU2HW4mbqYTfbQgi5v4N9vx20yOEX7wPChu
JStprbqBGTUrlJRohVMX1f1LVXASCMvzdNUlF6ycjK1tuqkTNLJ9LS+8tZ/yai7JyNX8kK2kNFbD
crxeh37XUDp8YYLnmKx8ikSxo/CVTZ7RIcIvSfx18MXwZuWPE3CORTZV/CKKIqylMqqSHhLV4iQq
6FCRxWxwf9APgVJS/lgRas3jHhf04qMMrLl+k7mgY5f6Amv8q9hyicy5kVMjsN8xEC4Xb5iOWmI0
/WZEFVqL1ah3zHddbs8VPjXdjrebL2FBH/ARnaFgMCIIevMtISTq4vvpnIL+guapXY65HS0n3FSi
afPyVVqzz84Hn23Lz69WT9Ll8pUsgCancgyHccRqpFtmvzdPyjy7MCbzpcs1Heyqk8AYs/sMVW1Q
VWr3bWwgVUt359mpY1gZNCoIHEq1c0DqVZEilms06BxckSoxoU4zlZmU8Zuyi/DDzjVyhr5WoB8s
nxFvaK/bYiMAqAc8zjTffLCkYgicv9xAbGB2kKQ/gWR1Xa3wiFqrNSXJtNa6qCDHIS1T3zoZ42Tt
w8ub8HOJf+TdzV1AToLz+OCgI5TnkRxmUESBSrk1+OUdS6ogoecJGJSDr+tKReqrQ6A2wOs3Ru18
15RwR639UF8sR2fNsRYV5KCyr4yeCyeXQBYbN6MwXBnRpwEHYwRdsq6GMDzm1r59MIHJNgX4zH3o
lEVV6K3fzM9hWy/z0RaONkqaNIY7v9vg4kneZ+3GFUI5IZTgU6FMJSlu3j1tCz3ypZc6M1RQdvms
of8kQGRo/iMjoxh9ILoODSCEKxrLQtv+i7aFQr0qkXilco9UyTs72wKvp+8DuPlNrwjDziIRieAv
+xSNilY0ObpcmF1gA93NiGV5zAbkMZNWIeTZ+nY1dhiRCFaP/pZ+RBkvpAOJMOCHlcSx2eM6FNSg
TIa5JQeimf8x0pCOyEKFVoDgHRxI0z6+p6ryR/JUoEwQkUUPy1bhobz9R9NU75qxBTAyLc2SfFXH
yjowBSgmxqv9Aghk1KLlIQ+R4NonFXWw27M5vtv2XDsk7RSjIjX9iP+/rtwsC8lXAx1oktZkKr4S
/Jdno3siuTSoCwO/iyRmtHAVKeKN6LuYLVpIdHpRmbRoV11id6+2yLEft0i5IpEFUm+L3qNcI9FV
7k+0QZ9oI/f0W2SiTB2cV1YhNkZs02NvIOXGI+AL5l81r/fBq1qhusYqTgsWmZP7Jk0KZWVz2dII
kOZvnfZgYnzIqGuybsSfVgkNNOkHD8ILJNLbd9h2FnS9WKcejsDyf3bo2oQbKxvyO52QnEON3Gn1
xPgPxNlHBP+MNy3M+oIkAjZQ+H62XeKe/dFRrC4utt3UejGGth5Y7wYvQfiTA+6WHcAE48sjJCD+
7sHlH0avBF0FAngwmzUReyBBdOde0IiAeuBdORW/7UmEQox+R2uW+kCCJOQvvjIKBpydmxq36KdN
AG4XW28Y8oO2E3zK42HqWOXADnUwIz3J4BSaxZ7s849fi22dV0z/J3g9L8HjWjLJf81/lL7xG9R9
AUsHjMX7VzuOe68wKBSLo7cE7OS7wu19J83cvtlIqmisgkYI0aU2zbTIU3XBWYYa0iwHhcxQL3TH
VnioL/oEyldXVQc5Fkeb+Dp/Pk+gSv4yJpyOiTjUMOvZYjebLpZ+VADVKJcRgL/wN+z9Fcvj9OPf
OODljIVKMUwO6QwTd+pWLA8KX+1OwK3UvHr8buRNzxBdZmCF8tGyYNuRka0CZY8BFigBMrUpO/rc
HBEA4Msd9J7u89hf21brlRb1lRY9zbJtN05YeJucoxbK8tEZGM8lSNSYJXQ3P3asYyTEuTSA55Jr
cGGTEWTYfD52gCbW4y7k191LiBDQAc9+dbF50F2Bp0Wh9Y8AuZ6c5QWkVpI/c+8ci10oqtn11fLA
6oB9wYflf6sR6WB/vMZ3GqVVWTagysxmtmw4ZhAIn2Y26V6XbExHsZJHKTgCyLtnGRPwYt5oKQJJ
HdS+MWuhnki70rWIiSOmbhIU+oyS86FFiiRnHWcOAkKoSDxlZZvKCIb6mgQVrVApS5B+Q3dyehpV
ZlZH4wcachbxzKaFQJkkjA5xSuiXhlg2synMmtXCDcV1ZSI2K6TTnuIhRuIg/htC7EbYpSxymo+k
pPVzk/olUYqSd1cheY9FdRaeF+OrwGHKbAeF3GLVvgR+2HbNkudzKoUKsDRrZL8bmt/EhoPBTKEy
A/zZZCKGbV8tZp3Ca9UBj9cgPwBsYJs4BYw5ZFwk/fpvUwvmG7Qlny6DyuHM5iM70ST+3FCswret
XEKQ+VDGOUovn+GxLj8M+wqn7F6vXxCYHKl/B/vl2hjcmu88ryfuOyLqYAaqHN1ytEqHCxO5ouY4
L0AppgqZeTzHRXZXUjjOssYKPUnEQ9pDvyh3fQ8ge5EJvOtQd7ZTRLtOc2tEbgbPv7paVBbxX/jP
ztA13I6t5P2fsyrFLlvzqcZIZYV++OIZpSV0ylbH4VEkkTh58ZrC4OUq5Shr8YaNNjXs/XdXQfAI
EM6BC8R2pMHWtNkJh3LesnVCk4DkTOUSEIgXbRKEtIjHFS7i936WWCDA7kfFt8LSxfAbbXnleKFn
vu2RGa6AD7j+0avPKyu8XXbktJ2UQZLHEEJhs6cdkzj4p64yr+Q1MWlL4FIDMcS0MZNcU/inRGH6
tnEZDvGcgin+tFfvbqmxRIykw8tEToVZE8UcvbnxwQTgi47vbbohz7TAWA3tnI1Z6I9UkG2WnW/J
RMjAfIFk8NgPNjePdwQHg5NoRwEy5ODj/FIbFOKtjhesdJrvOt6J8Co/hC//sx7IWJPvxtzJZxsV
oZUDUsD+lNjWs2cqfsr4uZa0UFJB+AbvrTwgAegm4DT6OwUKw+tGaqtBQsQQlUl5QL1SExmxYu5e
/4ObEaCOzyxWPSr23g4sxvXG35Boic45xibHiFihror1+M8dJrGq7wfBLKVEgD16cQod+2lUgXj/
q1CRkbarhkeT6STnw60b0TYz0qzh0ZFDCKvk4VrfWXS0Wa1vfhwSE725Rtwss9ThyCy5yD23uuaB
MsQ60wUbP1DOtxgpYHGIn8DIzeEEgH7gTrNA3TRrCDNo391KqkD504GGTrjUd1K03WuDWKV80uMe
L9MjRSMRIJBtjkFe8/SKtAMVk1Q7ACbVF8fvgpiqEZPnh1z2/JsJTV91lgMfaG8fgEDLpc1wGWa3
NRtjr4bjAjQ/oPWKKCiuoscoqGgf52R7j7BlpinugrCKE4sNgu0EvuIwoKVAAyTzDvEuKryAeKHY
wKrlDW61xD62F4YVWN+KUnvGGld7jeXYCvLRA3vlQAUysl+/2w9F5AWTNgpxSLqyVdhvkjpqeqtx
aliHh+0WeN1xcssWWCodgEMnE/mY2q1hg7nvBCVrGlywMWQ7I63W+2GUsZGEII126YDvIwMiJpMr
J/zQMOUmkdfKNQztPJjKhiZUfyJCVE3LRHH+6SfcNFTg/Q314oplOa6ookOhAAUmlkeh5oM+JkYR
xw9c8zM7N+KDQlHW+ekQ0buBGP/lWj5X/ZxKr+GDMYBdlbqturPS8nKWWNal9qaQzIuJngC5FzEi
qQRQHhke8POkzQqfjOuINq05DaT81VaxF0JguMrUURzGkBPR4nKkHHmRC3lb2trsoOrQ+KC2aNh0
z97g7w5rytyVEYTjn65sFbuMH8yLC3xp402Yw0obm4rLXzpUhgfJQxbM+gw2mWaDgCn07LT1TYaA
x8lVcPOBVcUq1huSB05/viLX023/FAVEN+n4m4Tyo6BT/0VuYvvE0zJADWmteHU8oNtLEbE862Li
1oUqZYdlQ8z2AF6FMTF3LQ5v6obnRSPEDpM/NlYxHX27FVjhVBgBL7qDSnMVc4Kzgr7pDxMix0+o
ZqFntecayclQ08TxGR5JCwM/M6UmMdPUMVXgyUUsZjPsIGhU0ykLOfJsBAmnngRDwPeIWGJqFTqK
n3dIIukC/3jX0D+6qbrBhraghIUGdeucCAkpTCuDL9neVGKwi+4qst5T6wyieWPPkhOWeUVrigm8
u10D65zkd3tf5S416rJiOwwofbZLshuQvP//Nq9zymcINvxH9v/Nyj4kQy7zsakm8KZ7MG9e4+u6
ym9VLJF2hLX8rgSimOAWWiJRDDUaG7ZcnUokiNqwvELw0+NcY6gpb1+PknVTAtq2QDnBthIJ56Nj
mFfj3lzmbgye8yZrqznN6G6QCK/L/fbsXXjdeoQzigBoJODek33YD11Cra1rTgriEvT+5vuy+V/a
F93KiNOdJuI3/eGShq5j2VI5oVkqAyhPXIcJ9/n2IlqG91kUC/kxu0PKVHlBSnKkXq+lCrvwyaYQ
rJiPhpH8o7bMungfBVC/OUnlIeFmAWTA91YwykACHvLFgPxS1wPxawnB+jDCR+DjLwYJbFO+ZExz
WI9KfixQJnX7NqtodfU9zb3BHYlY4w+3UdDe2fi/q0ZxRceyAFPSlPoJjI2HN2c7Ee5ndYwj2in4
X8gZvFy/ccjxe22W00zOcyh5ftNm/drfUTO0q6DX8cU1DEYqRxQ5lkvi98JiswD+n8x4uOB+jscs
zBt/khG0cFVik0StuVdv4Dc5ei6zjqf2f3Vqrn6WuX+QFNkQEvThpRPI8qKF7DoKJC8tpmX/JsKM
FY0fUgLwB67MA3LcrjJ6v2wJ+6UN6xf3zSwkRDTiLP5iqWq6Rty3OgVA9UbFIT5JqauEOEq5bCjf
vEAlY2dg/9EQ2hZvwfoEbj0fYLFvLS6tyQR4HXqfLGjvY7EvUrWtfqqTY3hM26uT6Mf7b+inM2j5
RD9XzFh2Y00oAFTqTpBzlEDR1ftbS307uu3d/HSIJI11FBYiJfLy8E7CF8PmwsauDdKghp5sTvYv
aZ/zRiGkax9Skq1eDTL1ZPB0+IjwfQN3Hpsj9e+HDOfWjoSGiHk8HrmW6U0Ghmf2LCKAfqrn03Le
AQEvOxD8+8TiJN8Cy7t2aq4cfp+rwTmPjhxntcviB2mx5qdj8NzhrDNNZDD/+eB5hOEJZtpUZv15
41apPKcNUCf4hz+2loLy9acPUpi+3WzLYphWjNFqgSjKhW6Dvv/M9dyMMJeoqKSd1cJrWFiwNzXT
oW/+6yjIUzHNgCc1J6xuI9vKpCHB3GHlni9W9eBERqumaf820hdH6SDOSUtb1V0zZNifKByfT9Gd
7Jk3I50cAFegcHt1TxtNJiCJG5bWaNtQFn1gdk+CCWAjrit1fW+YFTpPMiE8U75IHSq/ViloaYJi
yIG11DkeM5CmzoUCkfK5S2Xlly71IsYEEtZjGB4QPIReLOncD7VD/4gE2HfVTkHeCpPYB1B2GNBS
rPs/D5unnKKpw45At2O8gfzDjSWHJtZIm7kxpeCDs9BVh+x/IGrwOKdLEsH5Afk0gEUX+azNzlxJ
DRABk7rdofs7rrQuRADM2fWkg4RrcGsCPtPGVxeaknVRZla6HkTJcev5GXFNxuERS5FuS2fTxfvq
6LyEI1Wx5ycy6Xk9b7JvDa6mjgDksVYCb5qtqOSkdiDzfE6g61gKD6qRoWkiloEZv/WYa/vTs/Dm
yRHNKH4g/DWPqbkJC//aln0rvE0oQPOSbdv3c4Il1LKB+FAH9MvTuIRSkim9WjUxWLAkptTdjBVg
e1g4XUVTIQLdp1zIRtmcF328JwZTvgXcy0uUsM1Y5T5AE8lEafZgfLzB3LS6DUVY4Q9I6UnHL/qv
qVVQrxtq6FopHyDLOalTdX//gFWYd7u7V4VPjjI1xqijp03EXXySIghD9oYW2ZG8sR91Gmw+OBd1
uL1tl1xGvQ/0lPcAzKDxTpmzRyg0Bq3s2jxPyAw0TvgRxeNunF392ulj9q82H17+T3C6QB0rq5fN
YuJEmSaHpJR7yPgVxzs+MlE0Nb5ohQC1HQwwtN9P4siQcB8ZJSu7mdKOchMlUw2cpPJQiQTyiyws
XuSuYHc95wNdzZAOvpN7h1x3YYKoPriv9z2EGtYvU3FrqHrDJI3n/0PTGNcnl0WsC59V6LQZ8g2v
HXrjuRxmy+b/x2nrSCOKW+hSA/TvV2fJbBgpLLzklmIB4Y8vRlme1GZnUxM74dh/pZeIu48Ie2dp
0okvGXlSnBlV2LsDEj+AjZjgXW9UJ0z3j7jjowk4+9f8JEMCAOsFIFkTuse32/MBVJXAhOgXAef7
FTSiesg5AkwcETybE7d8gqRr1Z/EMh6FmCE3DSvW7yzSWn39wEVaciVmNUh7fMAv86Z8nZhIHlpG
Kvv6mqpXb8TbVCu58AUz5IzOo3BeAQFBWr0VpWath84P7pfShmxw7FlZCgfCHdRXcsjEHy8LUpeT
vTx0ZLtTc0I4BTr/tHEoFE0y/3L+i7T89keqJSoJkFkOSywxzdQEHPG7v9akOAjpCUJYamryllb0
N6u5YMJnjxF7nMYfYvHTj6GMQkbF2N6MmWshbGPAa7Bs4tS2RvbwLvnt1Wf9xOvm40EkMZbr3MLs
ACpiCqb3w59dWjpCh0frbgoh8gkIHLoned9oo0mPmgkzAv9T3pBP+Jb/u0LTX22Xm2ka87i1MicQ
gaa5xeUbSZcFw0AO0t9RDsUzM+/9fdpXrsKGF+jjlC2Cna59XOtl9LUuGnWhx8pUqK2JVjZhoLnC
L2OO22WTDIuymldd1fZ3XKvODHIcB3cwtFOGpm3mdsTQJs2T3hRV4xdqxzyEemU6Fzn9YYnRtpfS
JGopCsJHDetiT6ItElrKCuAb8pc96gsnTLAzgkagSZ1OFP9XBVXiREOYdol2kZckA6HII/YHDges
oEBgz9WP3YRIoJ4CQ15zYxcjSGWI+UV1u0pRk78Lom1AbgbSZm2SvhTSPQiIDA5Sudj76f+E9si6
Dulur4Yt2wfqndWPzP8BLFTaHeobB8uHrsGSi7hWv2Y5g3Gx9dktPHbwlyWz7NVYNuQRaB3IIrQL
GYqwGIC60vdaB11lRK49m/YgN7L+tENbgWfRTc8Z4hnsTtjgRhcM4QrbL3c1qEQ1/9YgvfgkIk9i
l3G3xPmf7Fgj7RAiWg8U6xRkBw2yqXpDJdm6mbEEwR4RB8sBSFdLlQxMm3AD8F3AlIMdeQh4io7m
gFl5AMjU6ULkO6i9WFq2TOHy7kud3xrjCPn8urC3sHa3hi9S5AwTTgJnovbEFz/myek9FlaIKvZK
RlYsjRPnwSjCSb6AZOOEpAHR/OLhgR3Ff0gN64hiQxV9BBaeSu+L74yQVEKUFxjuFrX4mcLOcBB6
MYFeien//xmulxyJoouszJifhUT97hezLxAgvHuribaadhKi/K0Nhpjz4qSbUnZmaJcbm3lakTlf
8BRSF7o/IP0NsEXjiJwd/ek8D+l4HEGu3vJUpSxt6ttUYKAf2iBvvdbCJL6EWNgHiNg9GVJw/Nj1
DUaYtYev/NHBNLRSIBKrolnMNwo7duuCHNABE5HHLktUdeIkZXNF7BYKQcotMM4R2qPGeJkrrRut
ZFmxxc/c0kWP9wwVp9F5OEHBCXKcqBCfLZOczY7oG5QJNucee9I+7sRfIOqyu/sG1fAVSGyqbYtS
J+EETBJ6Ybi7QcDLWL+I3rcjYTGXOJwWBzATlxdDNa1UIduqYJAdjgWDKGTgCJEfWtMzOrkNkZG6
ezOaQ93cRneaObiDzGJrHqxJJwm+YUtuvcAsmdot5+VnMknOUGe54v3LoMmfXiGMtQdfqnlXnHw2
Yf7AG4ccZ7PDWdgSwynlh+UimzBDAMc0rct6pxaEMIDiBnYFAjeUJ9uuMyfuPyv3B03B1fBjIG0D
iyl0nX9cJ2frsPBWCPdXBmB9/cNkM+GjUeo3J3tajt2ggZ66BYr8rLIwTKS1nEuNWF+FJkPVUe5J
UYwrnA8/d3Gp0Uq3MO0RKc2QM1lmw6SFq3+Z5lFiE/BknUWYfpIQIVybwb4HXa2ivOpRG3cA1K/4
7Y9IIewAcn/hBtX2pae66v2IDTh03cj2i8Z6B2QZVAHhsO/qCx2ZM3kn38iqw13aqyw+1WrBgZE9
l3u3kRWSKowuun7kjUzRgGB+1amvL7D3wUAaJNSlgq9DInecoMjTNa7oPaObXSpZtFz/JONaxMtn
LtBQVoAtuDlnonqt37EP57ux77Pk1grAG2bMzOqCU8f0NZyFaQLZ0DQkk1CYPfvmp5f6LI1CqXAP
ZaGgZ/1q87Rb/WzZIGZe8J/Q/voKQfbUN0Ob49f1VCDScF7sA9PnogqSv9YRazMF7RfmxMw9ANc9
KNzJLeM5wURR5eaE7eqZGIFExNXaecQXkCZxzL9IgTByB1Zol55V3wtqDdlQ18ZfCu/JVt5UaOXM
WVdZxp6nKvLR/pE2K7YkXwUlv4xrGW9rT/6v4osrtPJZIfeYpX2pBux6+MDxmGerM4CTzNsCYmJ3
vqT8AXQHmX1E+wHHPolXX0KtqEsmo7XIPgeTP2+4pQWRRyaLK/oUl7tQlSfzFygpRRIEsw+n3k7P
1KE3zZVK3UUkNnEjPDRJ3nK94NMqns2dP1xmufz7ZHKiiH0rdROg80eL/QC/2ubRRjeVaalNUCzX
U8WSHG4m+rHYZhuvNdOeZcZF9vOZgmc7iRx3QMyIWftJ0d8YMEy9OlGMYQyqxi8Msbou/PTKCeTi
OmcrVOGt/ddbCC6nbPTIhu/vIuCjGL1S+XIbq9r8OYGS8qSpuH8nIRuApcG2B/M8qxYiRkSOPrsg
e24BpRq4+u491xHxmLQdPikFShFoz4k8EFtFAKN6VVo+bdkobMlzYtL3lmL49fWhz0+NLsqJnlrZ
6hemmgYvRxA+JrJq7WqOqCtAd6jQ5OlJ695sHPZ1hxqmH66nKZK9mTZgtiadzNSkppCEKhoyivjE
D0woH9cpBYdROP79WoC8YQ1CrHp2OEwMTWVBxnZs2+AUOuhC092//ITafXTyrXLGpiCfPoe92r2t
4vv7H62j/m4ODsKEaNx54Sgpo4yP8/3sMT1AmhBUJ0kez3dgh/VGSvHt9FejbWTgy/Ui5/I+pTBt
piznHV3mYioniRdUHhCFYs2KTWwfgoMhbm3fxsdDfZGuzgZAGjCRyRIp/NwfPAV2mCS2ZkYOt8hK
EnTEP4KrHtWxcQtn1S4JuvrbkGxERzM1ky5aIuGxHO1oS9enGlK2qfj1nGvKPPVifEi40UEDRH1l
i2+C20a3icgisJU4pDcmuM0GzzCE2P2fX70SdkVcxFztaQUyAub2/WIpet5H1fkOQOAV+eXEbIRi
PMhA9z4Wjx+T23+aVBA5INsJbXtd2DkwduY+3DnRhUZgcVpvMMcuQEDbznIyefrxeqfYhWZZQZvi
BlY32YcecKsS/DRIYyub7NcU96bqiPCvXMdSW3jcpsr1q0tL5bt6qzaAojlzbLLMR2JpFypAcdMG
spC95fkltLCOV2ovkvNYwpA3L+Z9lxcV6EvgjNbFglnawtYGUwJYpcDVtCU+NxSJyOz5z2yK9KCA
0ZQdHOW1z4dBf6Tm34iLni15TzZ/SBdU1o6bwQrwwGjgr8SFajOQ4lSFfT9Zcdq/ReQGHEtBeE1t
WNZ1H1GDL6fxGBq254cPWRCH3YKIBxsMfppCw4QkS3M1yoGH9meOrAPmUzHrmxbdvOM8mxQpitBm
MnfaTFVX+Bm/h3sjI/Plw8QZHXkHy1XJVAQ8R85YrSxbaw1/WKPCU1b7XOcU4pqdH8OuiEfycM86
RtnfyoH7EzhjnO3SIYAXm3wTJ9t8IHp8aQlJnJFfr0MBIB+FEpDA00AIBQS1KqYedar17X4Wzqfl
k1R7TmOFGZPk8500Wq0Jwog5hwa2y8eGagTn46IqLsHGIkWcai5pkstdcWCVQ96Uayb1IaYKMee+
8i/ht6PsQrsToKGEdpKQnZQkj02ppsiNERyDRgSQJyD4PYzWzYElrZ1dbk96Yi/LHj2yP0nlpval
vAhKfuwztYM0jmA5ekcvzbVQIPu7kxxaAWO9ZncCwb4NWFFMJ2FWaS5bi3Ax8WWzTWcK36wz4WPA
+4/32ZNepAGXBFinw7r+d/t0xKYAhqf/GYcliDNhNQeguFtbjA6OJllfH8jjtqX1BULMsXzTKV/X
zA7MG8aLINC/nQqv5Ogh2tnaiCy3TbFwzwpQ1TPymxj5icIyy/gB39KVqPtQsG4aAO3WuevoiX29
CewBJ9irvl202if3gCNggwN21gAqztA/tk2LdlQ41NCEL7EVHHCQlf2uuRu3A8q3P55SDMezWDDX
yoQzbEUFFa3xMUAWclMEjodjRJOkXdwlswrgp++6+PtyHCXesS6Cu8QvKqYqc2Hc4ctyIxBFCylU
4a0CwLuPDqpKpU000aMLh8xftG/QFKczVsuZ9VvxPNOFcEh9hwH5Tw/NJlgJ9KWZhN/gOJpkhDqW
xkirbZBdM2cp4yl/X/wnxvBGdMXkx51qe4TBryScfr21bmJd4D15bOAYQKY0/6MfA+ZbLpS+EV27
i909xc2US5aMB0jYFcveKWcew4l6XRUYeCPmnOObZNVuZRdb7c5kGPB6A7b0lyElblfuilTxB1yz
90qc63LOLwW8ucKF/rlm3BAU5UnFY91j1J8ZNSTVyGEdwhjBESl+a6BwevkpvRQnt2yXxlVzwDec
HgQ5VcluXFobMNQjy1Fwy9UG9kKnhUWwP6A1HTq8BgVRckNKsGgRr+ZUF0SWZGKpohKibEI53K9X
4KSwXgmQlS713gdZvFdgYSiu5TWzcFUOXpYEUkEmfvao0Zsbl2gH0k0HwAXS5pg14GSrr4TxY2P4
qWACcOEpPn3iNs9Zom9v4Ikiv6kA1hCuqW91Xoa/hzoH2mdzd0nMo7jvC48MCs1X2Dj8kn9p+dI1
lsVSX5xLKb+xwXZ/9ysv7CzSy0vlDN7erPrr2IQWVqKOfPSdiwho5bT03Pdc6ONnJIsLE0K/kJP0
n2OqDTfHsTdpb1fnDulIrCkJv2n77R8JL94bNfaQstBmZxM2luO7P+sG8tdfnjtP52+/uwmRkIh5
JCAWO5yhKiZJq6HddpWFEYEEfFdFOlnMT2UDVog+jECxHpcSPfOB5NHrxRq9aVmY0+5uFV5X4AVV
g6kCmBLgwIpf/6M9kdGPGSUA8tVybjmri/tMaWulS/PlNHR1r0UYx21ESCkcVSgnUNPlAidpbn8G
tXsM5TFKfQlUPUVnxvqcKi57R+9tSTANJQt7JA0yp0BtoCzHOAZJaaZ5jj788OI//1xi3EiBhWAF
f5Pot2umMVyqehZ2KQZvkeru7SscnakeVn1NcZiXh2acRrVGdvDSM0Ge+8qoCpURbqVLrGl2uU8j
5TiBhCZY9wO3H/AFVVQnfUznYGwMng4VPTkr+jMqPnXYOCNYckP5LwtDlWC35i0FYyaCb2fy16jN
nuE7JGFWsmJupjLZI3d32T8ejmn1wxWzV91QK/1Gov0b1DZXbtOlofiGo/RlJ5t1feghhS58UlEt
oh7dRPwsJFuxySYBrXKGHJzOBQhU929Yq6xTKOtVsvb6CqUGCGSqyapdq1phah7Qrb9YXmw2uv/+
9ywtM3rM+jLgiLmDcaMYuE7PNVGnBfpSrB0XIX+uoC/D7HpJqXXHn72d9vwNssAT5sPhE7OGbFUK
vSkW9mRVXWNDKX4Xg8F81/Qa7lIHsNWZIkE0FR6x/WdYkS1BXqi/ghb7/Q3I2+ZKLumfqFQ0elmq
XzFSqOZYVyM6g/RlGWrJwbBLbkQe2rBR2lXXhQRle6BjnWMO/WAD4tXWCfZ5HbJzUnooCZEVSqz5
HFo/q+KTFTQMuhAyOo/9Fo6vC7DsT3wUnQV1sW5eRST5uSMh+aVb9MKfsuFTByuGOaQIWOXN6TV7
singzpuZO4CCxDDdOFPbP5wKfrZErz+RerAGGaP/Nkq6KSQmeQYf3uHmGpzfmjErNYYtPG4KweRQ
N7IBoPkAaMizQtPlZwNOIb5J/hFB5vH8VUf6mckD/t3DTDPLtz9qa2uSGTT61pD1QrHpjB5KKMpc
wCaVq6dMiQeQbezR6JJwWqDyEy40I5fWHRe1pbCb0EIRnoAr/WguKJ5JNmlgPvWovt3OOuZhFr2t
8HHKSbJ4zle8caIhDZDuUR4k/wpDh6xUnDg3wlRQhh5AeL1/ZgOemJtjb+a1iC+nfFUbDziu64En
vDTivI4DFIDFVPqFBGvkU9rl10i9bwRZdS+zwlehIv5yYs1GgLCZlcPkVzR5W83OQKNX8gNrYW49
Txu8/RLhq7ixhb37e0to0dT78fGSFXFqEmb22ktBnZmoYSw+oDBYkyzoZhjH6g0eWiopDzY1k4Qk
Q76hso53ZPhGcwosNYP2BT0FgKCh0+7IKKM3Thv9pXY8wjkUEFGd3MDPiOQDRRxNAoptdRSujqhx
QZ9+95WWoP4fFCAwsls34tCZahNgu0EReoimXk9qLPKZzX3wtoITIV4QxYS1n3yvz1wbFd0fk4yI
z0JAuOyt4x2FCtNNjDuWd8ZkQPjV9jaVtG/XKjuQbQPRKzoZOE2ds+d6KcB+x8FUzOhmBgoJMZqC
VncYPzYeMEvE2WODvdPiVHzPlYP4T9CPjlIfQJiSgEpr17rJENeIhSJwUxAPujAoGS1ywjVkLFkK
tybbMKQRlZSS/C+rqRHgjCyQhiQ5+/mKNB/arrL9rt2Y1v5jFnnQDPhCBpJZxF10HXyrMtwNoo1A
PJQqN4b6FN/Azf81SKl63QsTzdt3y39WSHWO2uOzaMB3pHLbtwNN3NYWO+K1Zih0kDqEE8g94SJE
7hsHnpfk0UcB4j4hsCK0dOgjtv7IWTYRnnHpgcgU4TV/aK9dv54UCq7yxUN1NhaQoX/b1G8GUMHj
GnuSbjEh6OWzna2gpSCZ1Z4/TQSBgRFU8MapxeR55QNwY0vxBffbxzj/eE8ou7pVzJbKIh+agXCe
pQJ7xuq/oq4AqE/zsSzkv7h0UQGZnf+rtxYgqGINVTAgf47vFwiOXha5R+dC7OSePgn5DR/58Bo9
YWQukWFbrUGSLps1Ju+iqhao5NaYpaENAhlNMgbhCPADzMSdyv0YNH3ibDuJakbrgWpyMj1B98iO
WrN8w+R5z2YxNon6xpuFzMaIvkQaud/NLbhOAbAymwQSp9G5jnOmZV2U5TeO2BU96DBoBAk8eewd
pf4RV0s4IqBYOsKoPoIxnDHCOUT5QiVWKsqu1J9f1tkzZOg/D/vkv4mL9WsCiZsrR6PF1Hx/Y+OO
fl6Kih4qygqNRVZ9H2qLpQk7NjQ/WXDhhzsyFWMJvnegpEg9vUnua0lHAdEk8dSu7vuCVZFXueyF
okyAB3FFMUtHe+2YYoE5nxR1lhKUPgPrQSMjYPQEcoriylSienxu6Gb3cFH8nXxwh7g2NUyV9DW5
SxlS5Hf6SiZOmrqa5yAC8tSlIRbF8lreLTi/HkmqmRysuouwXrJbeA35fOe5swbuIkJrAOt+YAVd
XsrWqSz3AyjhlPnZ3QgRwS7w9FqprSENVN0Wj8O1M45cgjoeXnkMHdHMWexalFbwQr7TniXGl9+k
Mad2c/72UItGhIEm4S0xyoYxm3eqxNHBwi+yNza08dUA5J5q5LsftRsUTwCaladXPMdpLEQwBVVB
TBGSI2hW9viquGbbNlwr/rrIhOKDkXF9ZWY23Jd5nhKhfhsP9AUkTP5eV7MyIJiVcvFcBC+ZgLxU
K3LSBJZmEUWTGVgrB0ID+sm6e/h1v7vYyuPnPqP5C3vJJ+4XjsIKmbc9uJUcsOHviTRiTazKTo6f
I6kNZt6BgT8dOUDMGEkap9Lpuz3fe/5JdxGesN6dusj7iUrClJDjmS7FrdfRPaFolMTFVrAGTbpa
R+uI0No8IbjAxA8XTRCHLQQ/jEETVWqLBVcmmGtkp7Kj9ppM5WORIRk9aoNe6q1DdppCDBNqXrwA
gQ/xfrq3xUIkGJPukLeJL+7TdC6aaHIk4D1c8kpKrBsUE4ztcAsWcn3aQ65y96opV29P05ftigNe
yzcMcH08MsnGaDILUQkCTCo3fV3EjgqXPsTMh2bZgLog1Hyz/Ndd5bSUPiA46qcLudb8l/5vws52
7ozr7jRGUWHjjUpX4nYV45+1V00gir46PNVIa+eyIe96ksiW0pXqN0TUV29mVPTZGY16GTlzBCQm
c6seaEHu3lyQuAVhLReByJ4jrmlW5jhPCj/4QnS389xbNTUCTz8zn0iQTeQPBEbQ+c22u/9qj5PT
STqgy4YCwD+2ysrb0st5PBGelROSdePAneTOKkRGZzvLWq+D7g8nSjOubbiOPTOp8QPBzd37d/SV
OHDde8/b0qVLV7leClP7p8pWFgrYAtk4iiA/yVdPP61W9ndDQI2Ym8tl0TxgZjRjn9avO1yhUVKM
MdiI2gdo/OBLqWlw2sf9d6w1nWcAtcl95c3ya63b2K329Qs/nJy560jV3DBC1Az7ZgjjjzfYjSNY
Fh7fjOTQ31ns4upV5mH9Eh3MBwMj5KfLVu8n/mbsSyrzbPwrctNZnl0H4nc/FE+yS/vFHbkSRf0R
i4Dq1whFuZx4PlyHDUEOOGePnKSGubtUk9IbLN7Z4si4NIX6QW1ByMCeekfJo8LvwGEOtB2NcltS
sZaPwMmQ2MI2QO/HFCy1YZaUcX9CR2N92ZhfuMlM97Kk/qtxTd9sH4plCRyyLIMujEaaKpq3eCHJ
2HFiWTuDdhpysV+h56Q9LOdketgE1ToMYHdZV5XSifF4fZEKlHb3y0Jso69OI/KsO/74K+8CGSMA
3INpzvT+5yZLvEXaNdxPvrS2fLDHwBnIQm4p5DWSbrPXJNuymhEQ2YdlCpcLpgwbopbiTmyQg3Xe
YXAdCWlue7m9wEP1L6tcplF6kBCohY2ehGz2tsgFvIOL71JgnYJ78hcGJLdKbjzwGd9itypDp4yM
l8LLrct2vkfsJNTxI5trhabNPQNCotQDEcgrtyEQAykf4cGw6yJD4f+js6dK25cSvjIqwTmTPUD7
KYeg1YBNqXYxdiKFCHSDH7OhnmSQE3CSrY3QaOlChKBPBdA2yGaXLwoNl75LWtgE95qsnnWPMvry
N3J2gp0z0uM1hn7roS7pepjPwBgc6Ysp0a2+YyBzaMBQCzMyR1a7G4tKKxzluA2TFiyqWVo+UfNB
c5yC4ZFqQyjZ7sZB68hr8NUGnegr71JLyaN48Jx9iTUtz9/zNA2hqXmrCyeg9GmWUBtige1DiF/s
O7HXj3IgS8FTI/QTMzpJy2i66xjuEbdBveMdFhqH4UMsJSX5BmGRei06OFwjQhL3ThBaYPTWFby4
uaOeIkqlS38kQDXvXyd/M1Nqs/05nkZlStkdxIa+oqdlMjaMlczRao9k/bfA9RXy09opoXgmwp0H
IlrlzM3pHsC0a1SuJeUe3Pv/2NQe4fybV3XFhqvliJr7DAuT+h4kIrHUxU2j78Foy08l5d9HQ00v
mI6laVJ5uXGw7kRc/vf3HstH64J78zaTLTrjt+nSAIS+vBCVUUR60SDaaghJy0RafEq/YcLAbbBc
XjRFz32p4dFXa3zstKwwG4DdoVjc8dO18N8aBbHFgxbK1NrlnEaidVuVFjgF4gx9lkSr2Ecxwdmw
RKlJvTXhSO7KXfPqxB6EOSte2PxYC8OQ4LkVphz5LfMp2wKxqtrCPQAcOLFthox/eaRK73r3ll7k
LR5dV3evVVgI65wziuwI+GY+MMHcbL1UQ2a6iBkiLZNzl3mXZoe48RNr6BV2kYREWFcTDwl24/8I
J7+vWflssXhu22loJf2sjwPD3GrpCWKwWbn8XFpDgwZvpbMPb55H/9EzmQeWVUgZzimsWOSzwF/m
8QP3rKVPuntNxX5qdHh3y3bcPuhY6P1vyZQ0Cdn5mb4g45gqL6hIixjtBPQETbfp5v1V3xM05J5c
54D+D8itYbk2fqbnMxiYyOaHD2ntkE9vFC+JvQlPg9DuxdKx+MK9ZtjENcEfus4EZ3Xd/BefeRho
1CNordzURvwehslj8D4s2lgc1NiLq3CE6WZ2FmJI527HYalVUINngILYoAhSRl072XDYfBONu3Fl
2eOvOpymsa7w7jidiKyKqZJ1Rg1oX37MSF8ay7Mi+SFVLggDUDO8MoBTMi6kG1p0w3xn0207wWAP
B4q3yjwVUkGZrGfIC9GAltiYU3dnWj4kEPziUWmg3xmau3cKGqZI7zsBKKJZkY2wy1Ak7wgj2Jqk
egyqeU1sdjIwEdxVpRptAp6SwK3uX+5Jjv+Mz+kQWvDk0OS+3iyjM+/ssRJuNIEkukprLNX/MXqm
6dR+OcosgfPmwNQhRELDh7pi955RfWn71dYNqDbgEVub3gjp9Nnqzs2hbN/N8bcwnSTbGuGMb+C8
Yu4i0Mw1nQftapO7mExjXZFotGoIofY4LouidwAYl+W25lGlvFAv86a+9kCxzZriLWHnwZlH106D
U5QmPuNvBofVSQN/SXwQm+fIBIFFq3whZ7ZMY8UDfK5ZNcFwCPh+nhgB0+fPOSGK/13zN7Jlm6FE
3fjb6F3H7FnwanS12oNu62dSsV9RZ8lWmn6/kHDblgXNDt3Dpp4AiG0dwcn3T27rcK0KZxHpZQH0
g0PYw9bPYYrPXML9XDvH0xaa/fEpqmUOsTqW57zdpvZ5ZQv5UtYhlZxwfqoaP56hnmNbExXSRlQR
cR0Px+/+6z1OCprV+mGBHLhejq9/D5MN+5HIm9mT05caPIewCZHSPgS0W7YxpGem+MAACGZzG4oN
zeXxMAjeSYpHLpE+DR8EMjfROTkvhmfU/Z1pV6Wxn97B4aWBlQywIePLeHL+LYhnkNqWMBNRHVd2
wRZ31/Wxr9j82416bPOINWTnYhvkwO/DwlUXWAaJEjiZ/zq6owMn2vp0pXA/ebk2htXxsBWE6M9k
mrMht6BbAC1TjsTx7wLib7iuBXR8P1JLejF/nL+hktA+ELOYF8Oh0a6C7T9caYhEOGUctmWlQ1kO
e4fNB+wH9pzv+w62XjW2BW5eGB27RnsIdZQZRgy72wQyAKcRNO3K18ARNRTevB/s5VNVQ/IuNqt9
/0yHlMLL6Brc8VoOM0zliev14gElElCtBrXIuMzXtKsEIGxOuCVWWm/hccloP/QZ3Omxw5QZd2uj
vwhYa49Nudt7eeJ2D9mtjrloliqY+EW5WJiEccDmxkVK+5o/0tgeMvxiYGcjCFXoPktYKqi2Z+51
ZFly2Ab2tnuPa3lP4qbrGWNnY+wpZFUPoSM2f0YWxGvFDyHXQ0fg9Tu6fk8VmKehbpA1PryUjBZX
RK5T/tIDmfBRctW8KTkg3OBrUyJN1SZiWYkq3TJK63Hd53+6FxX18YSLsTo9rT5CGN5djkXJeG5R
pyefY/cEhdHqMl2XbWuxRA3vKfEGnxmrVdqg7q9zhJpsfQaZY61A55E5qeSpG2hJlPFId+pE8dN8
3AGcn0H2G3TevA18HyVbLZWFlRS44Hbucx/BC6RodIpPwCeWcUw2MUZEtiP6nXXsDIkuFIzWHV/Y
0FYKjy2jhTZcO9H78IxuB0OIdWUKwWG0qMKGVFHdBro5tX9vUR7JKTZ9y8BPoxCw2k/GTedjhLsa
Tkzph2apuCg2ApVriJH+u4jvEeWE53nVSZt1k0Ch+sBkGmFBxG4waRJhTfahwhkU1/uriVR471TC
duXGy0BZq2Sd+QaA7mhFCXYUpKIQXthaVvcI8F0BQlXldM2P+xR+wvhgeSgc3FW6ZGo4U20pc6I/
ss2OQonnT074xlXuNqIttJEBRWhNtumxgcKpZFjBssItC+pUlo5R+spGh23XakuAlaEBb/6WI8PY
lDCGiGt1mBH07oFzl18AplGTnDskKhQDmQbaSGKcY6lbbl6rBGjGqUVTg1Wf6LGCJ0Uaork7UT73
mCF+6caIClelBsnI1NxqmPNrTSsYvsh/zr/uzuCz5pek/2CJdUQv9eY83UJI0mvt+djVUIJwSyWG
5n5K23KqS8ijp9PnstSuKyCB+YQWyInocc6eLcEohb1le469fK0G2dd9RjwaS/pxHXoGtpEG/b22
EOrleBYYTPhCbp4jd1K7QJYaNe2T9jF2s37kY+NC7fZ07JDbwxCgU02dYw9fzyZpaO8tIzg9+rC1
BeMh1PMt4uI1rVofIELI8QfMJUNXJHSZs0AA96o5Ilcv1YWbTqarvu0JrCMy2996czy2KjmQthh5
AwmXs4BmJTI5P1/ndDW6rO2Eycptb4qGq/dIhH84Zb0zUpGYkeKM8LeMphzn+O8YayP9ivmaKTBm
RZpd2h+vRZEmR5mPTPSr7SnaCMIXn2hJ1DKIJvEDFBrxWgT/qNitd2wpwMJDvmoF0ZMz+zc4w7OB
8DkwL0g1Eg8zJZn0FKjCidAl1v/8T68kHdM0Vj3sQ37ox1osT+QisgpR56wyd55KWQb+2D54T378
6QArPKvsqWzZdqmAtS6o9LiKXeTZIMCg3p3bKHI1Gq97PlwBFNc0H1l9w70bOE3UdRfTZRrXPWN2
7qwr5CXdIynrgFaPIqeuoc8deMJWu+vq76glO9tu5Ux0iAPQMU745hTlVM8HeEZH9zUAEY357LgH
Trc371BaEHTbIU33GzgZRSbKIT3CK1YgaJxqySIlcAmq/Vbn8n4ABBHEw9Tat/clQaR7QotqxFzG
R/4MSQ2hUxvEK+oueAlF4PwNFlMZb9GZFuQKfaSXwpij7FtPiHXgFkm0g8BwFM9z7AXJ4MWLcyPR
OwyF4f3ulSunv95DJ2wPWVYZ40MEbVimvbly4hbuJua2ayfxFtA8JWzDNgQL6rdumYnIU8xyQoUF
zZCyhN67YxnmyHQJwVmnQR/7TAt49Y4pjN+r29dX7LBMlh5+DzEZMkLsvXrBfAeHLJGLXv5jD1KH
CZ44txyOMY4urN8SYE5S/JH5o9+Eb380NIkgdQom0mQuiTD6XvxsjZzk+DPePSMSJlwL6L4Sc1aW
L0QReq9hzOC5tJgv1P0Q70jxIkojmjgiOZUamQbuZKYnD1S8jcyOSyEak/LUSs+QnfRfh4Qi0AIz
oLC4jQ4yytbM1O5UjO1stBWUtATdpgDLf5XUvjuQNqYuUayq0v8I4qwArXBFp3MR3xMjL+IzvszG
RmlDDWTXwiU/BBVoSbrDuM0YYDS7W7f4ctdEE6kpSnL95q2ZV4KumGP6mu3YzBe/VTA4KeJnNE3t
MEwRlLrmArqXtOP9AefXWarrN4iwMTS6q1a8p4M/IQFk2ZoqkBAcfXnxNNCMsftUMZfOi7qKnSIV
HWnygp40naSiMl2hwZfl1hl62xZhLzdY5wWNxP0RjrHivXzh1GRIQk+W/ohJiNRcFEg+fKtyiLps
ObSqwV/c9gh5MaNUjLJkCA0eOkUJsgmpDJ8NxMsuBMVE5FKxh/iL4uGrViir1GaP8LZ100X6WZrp
EBVYwZqsxdhv4XTdKSRYkk3+K6yyrgW+70KSG9s6K4TJtLVir7gmAJ6LQf/HntZJtmz9/ULx9krD
v2FCO6L0M3PsMHIOavAAnyOWWWEvJlNlTlp2ZRkMAg7STbNQXmEOlSekWrlxan6R79+Ad2b9oFcO
7m3Rv7x8qz7nisJpRJUu+KLT1QxcV9RejPxY9Qs+0HvP/wr/uCWiKR7cjvbT7y5eKqShRMAU+7qA
x8KtPJb+rr1GKimnHY80YKakaNkWwy2DC8xkq0v7tpiFEPAp6ehYjShq/l//WIOzLY55I6C0SjYB
OOCJm7tU4yhUQTju2onx+J61IUgzygpRriQyc1QMpvi+LmqNAw03fPbTJ18XDQ2DoO0N6jxBInZG
ynvDnLT2extUpF2IiMlN6tguvC7SFtlAEL7o5tYhd7fe1cYnJjXTDHtC9R6j2d6bGXblqFom5ozn
5aTCIw+YU48acZM7CVMS6Ly8hiEq31RhCk4j1dOaUSA40THADs4gKr5ShBgFu55pBO+YwaJyq4mr
KbTDKZ6iiv2VrsozD+0QoKKlclQyPzrMukJ37PTUlWvI2pt+nSTlfU5f97IdpYWUP0CcOnYN93B1
Tnwd+T+IlDVHnh4njFM03mv446w0xcO5w96z/042ITId1fML2O9wF3hq+x0TQdRTNhx78dKtsoLY
VhOfE5eijrXXlmDSCcQq8jKypm5fWDP4zXgW5n14JNb73wv05JmfHdlP8dnOhcOr6hQ6F10iSiT9
xbjfFaMVV0R29pKiygkjK82Jvu3AsJ/5xJgrV4jEnwJCPBNwr0HqGzcCtm8H6jtehDFfVKhiD3wu
YALCT7BE7WUaZWjQj1oOPmQY5wFzQ3w6at6USYZ/GLVdZFKYImlWuGRdnGfW7huphRtdY/FUusWQ
SsxN+t6fx+qjbuycVWVgQawgrRf5Y6PQKX4O4PpcL7BIDOVJWHRJ2qrIbVRD6h56WDIlSUq4OKE+
M23k+CGSJmbEBCjfQwLTbgEtuJxAEhUbJoyVE/Nn3M5RN5tvI55P7hoxrrZrbxVdIlK+TmgtUre0
uS6z+t9ltU0z1WFsywaOl0Gbq1zN1/qlzFOB8ronpD9Jxcjgt1mXMDOC6KUJ+80MuZqqMQ9owTf6
G6uH76jxbBhtcrd7FDmfRnz4rNAhZVx873poq/u2i2Pm5trjs4yArOyMKB1Hgv61zNogwadAvPPS
zZI4U10fvLJQITvHN9dQPZIow/efXyDOfPDER9OwPWGeSyknoITYaabGtesFKbsf2f0Ujfo430jw
lFE5KM6ySCCMRnvLrIag0R7MNMz1QoAis01Pis2+ZFx3Eq0Z4/Fe+L0V/FgAHGcxhseqFHcj/tUE
Onz8xgW3OK+ALNu5SR6xhxulf1vlj8UeNAkQL9Fu73UQeCGgMQCDNjHcODFIs1h6XVA75LdCHmqE
ti9uymaxlmM/EVU4YkvdS6iVCuz43JV12KHsOmAQGCzhf+B1koJqFAOK6RxcnNS+TMH1+YCLc/Rv
i1ptj+CYB9S1/Er4/kFwXkqvv4dDIX2qBlSEoegEt3KV28wPmCzTyfgviOWRC4iAh3i5fEhHwv4y
h2x1iibxCbnZw1DEwLf+7Fbjuxwban46vBZO8d07/tzTE4qg8jMDtPhJTNYD0USsxWJ5Zd/SjMFE
mxhBZ5tVb5R1TXLUCXKvzKsl7ils6//ljkQktd/lQe0TK3kjJtqwDZAL1rcu90oTKOvQvtoqqsNp
4fhq55bYXZfZ3a40+w9TpAThHSrS0R27Sz/AgmRU5cS0OoiJEiqBLfFDfXcR+zxavRv2ljm22kd9
HYPfHHxcMdFMVZS2XB15S28Xvlj7F0GtsVHxWOPkPZG+sIOewM5ZSe6eLlElDyF9y51eB9L1QZu+
30RcLx1wlM+ZLouYsSmIvKbGSr2UrHQuuEf8dm2+H/ShIRSX3bIz5OZh4or88KftTEIooi8MJM7s
jEuZDSX65EhXFDx1bsjr47Wfj4K9OLpI8NINWzVppRpnF7++Y+ONtYG0/STgX4wwjTRsb6h9GXmX
l0KNg3AkgOJO18A4Wqv+I6mdLGXyjV7bE8YGToDD2acJfEWPUClF5j1rsw7+AuMmuvL5gF8fqyR1
gGWi97EWcC4B43gpNlqYOXDzLTAXWrxJOOxDmqM+Nznj5GTIg1D9fw3m8hj4aRdsizNtwTBdvgCK
AScicxxf3mgDjGxvuw3AUo4rnCn5nrSkmet8SJ/7EkGCxivRfznN+Mm0V8swQlud3TW9WZHit96Q
JI9bvyMJnH7ZEGu/eV28gycBh+T4L9Y7jB2eGXmFpCeECB37C6yEYAm6uO+rOrMhDnWbaxZV5cmh
NJIFqOgxb4uCHeNUnd59s73zdGhHdX4pfSvm9A6s/6cyGM3zCALWW6Qs/mrT2MRmhL51m51bjiMK
9RKen2xXm+nsM70OPLYZUQXssfxh8ujzNqqPRc51rU+i9ZD+CZhw9o82D1gRtf3XzSARaXZmfZxh
A1zXYHp0c5MGwdVtO5VNcqnKz2IxXWk90XaT+g9Hp3X80gUqs9m0qvE6uovP21rVXLjI+uc5o+fH
bJCPXPSlI3lblvAlTAumo0hY83+HLe0tIgKAYoSddL3N1fuoHrfdMmOnYZHyBTAnreY5sCxA1jjp
dDNOpwiL/+z3xNjj0MnuiLX1bn7fxM52rDAwnE+ZE2YIFc6WOjaO9CoRk2u2/20nSSgeKJBawoGU
uYSnYi0TjTkUzEIUQUX11niTh8WfoE9Ujo5aEbA5mwZVvbYisymE1YcYAIB7ZcvNiKJ1NDmsIMZD
mD7b4Rfovig4Xgw5ENrwzuN8eKTNOuUYxpAzYo/I1nWyhQgbAYUFuhkiH900vm4gnrg/blDtvJse
Mq+Q/uQXra9bj1GTP+LFXZsj93QjQ4fkG2T/ZF7ydNtqkmz6TssaxHWzmR7nUBZYAqFDBGGIiegy
hzLGxH5ymQ9SJ1ktv7wPhM6wcWGUTygqFJlkBQUXfqOpl5nY/9YCmq5XhoKevOtQPUPJlCWbnyFe
OGPs2t0Pmq/Bt+uLZsZqEZLxNuCZtajXR4hqZpky+pLfvhT3rwqBe8nTp4ZHv38vr4LZoZWJQlaS
Q0U8ebIyfgCvIWt/6W8ba3RNy25dxYOcMqAwKzphiAPohn6T5xBTyFs/BwI4KNl4TFLKGI6Dtl42
SheejTdg3uQ7vxZbVMrSg1isUU9v8Ig9S18BiD4mUiovVo22d5dD1lxjloAZyB8QLytZ8nGhNlt7
DU1dVZrcYVdHuH4kfZzBO4j0IHTPIIgwuJRwgbxHD+fJyoFoTi5eWHOpH/k+7MvK8cYlIzfGuvA3
cWO2ObJd7m0FvsZ4UZ10ybg9HxQ8gwP20x8urCQ+yLkdux0aU9q57JwsRar+gWpF/UynQJaE1vzG
GdMeTQ/ZAJFbPXQSSMSxaBxETPebLmC4r+0C0vMZfYGxPQ6Spge4ZSJJsw3PBZ1o0zl/ktiWwVov
DgiDV1LJvNTnq2teujDMJpbdUBCYhtiiszkwqsvTsqErzDxIxQRufc7KGD7yW+fbXNrP7N36vE+F
wk1T21Rk9RUybutaL/Y03QYz3xFBC5XGtmLxk72YQMgCYVpyO99n/K6zv2rj1RmM4Ode6GY6KlFX
UfftK3LHAZpTPSw/NHECTLirHJansU4BbM68T7qlu3k4IKntILhUGy5Onko5mJi0ew8Io/y60013
s0hjhtiPdzgm07Vj/RKowNM9b8THGH1OmDmeWO5yWS+agtqjefgPPBfVsd59GqdWnuQ8H2x7NxHC
sMJsIkzKukW4US3gAmDBGmgNRbOWldjUAhisovGRyZwdAPzqaGlU8oSwWvJw2WCOX6ky/2WenPaC
HtIvY90OqZEBI0/RSpDjyDxTuzQm00pYhHY92bM9tsZ3FRpzALzV1Zc8tiVHwekFjraq6G+FgaUW
vzWv6D2LwgM4ZnKCL9/V9kvxp6EaXXX5ViW2wk1n097kBWWbPQsOP7ifLoHbJMwSsxC4PqLto/7L
/CUd2EdwRl1KoYD/76kmc+eitc3ibOKmDhvf8xzyzvBnSg36EtGi4iFknP/+7a8ahwZK89lP/D/K
kIURt1IKbFKlRlTXeEQQ9WAd4zmJSQTASjgaFdUVBJOgJFIr18pqBNeoPYfzUXXiniYUUluvdOjc
rwxkaxr+fzIzaObJ+JAJqsnd/YP00TKRm0Gl7/Qwnc5bji+QT0Xl5sHY3Gn42hprFpvKW4jTdjiZ
DWQQfR9GoKLkghpcyrZ3Cdu90EeDoH16CM12XNwRls84WFI+ERw/q8HMYMkvUQ6XnAQpvSkpXYev
LpNR76rnQpSxLK6oPd9BtXvLbTAvewYd3ZBgOJcjASoTlw4I0/oz5k/0Njdy26DKCZY0q2EQCySt
n4NfG8iv4WyRNVcuF+blnP5XXON2lQjxwX0r28nmILKbOv7ylGeN0SKaDN9Ke0FVjCGTsVUNT6QK
Hpem9F0AtzICBthv/0ZU0r+SvnTVQUKplh3dSCuBluaYy61atesywH0oFjEtwBic92GCfqP5Ff51
5HbNdw276ONzgc/b5+WpftqNe3Q0hqfQABwLUQm54hWi80S5seIAmVMMnsbLCYj+tlzUddHypjEK
t3ezu9q25Gea35fQptLen2d1cpGlz7++r/FvkUuOEtbHjxb4ai4L6VqzbuXRbwrh5LvQVAe6hk5H
xjxRVmBkq3qOULRGzjfueuq5Mj3m1zBPMZvrwFlnepJDKRyuejg3kPaKWStcIVzScs/oj7zIel/u
RLhZimUMjsUVrgyqIWSvF7SxM7JElYx1KZktM+tnSMOUd0HRtSFUHl3GfZuO/QSuRgqHrs8veFzI
jj/uhgHMTXG9i+MwVZuE6mJpxGAd1CnaDY+KpGqwdZhQGAme5jabUJfOSr91YxGwc6hzL2KEjYZg
w86zPKaSRrpSw/YJukA3f1qZB80AMbNZ0/u+zbz5rQS2VwUWuv84SM0AG7YiKN1kQTMRIT9PKuLU
7DUbfK5HUG5S7u9Wk/QhTOs6TrjOeL6pgxHpINSamAv8xW3Eqf0PPhLs7DNxGD2tW6UQBQSRgXMr
zXQY8pkYyJPe6B63WJlQdHUCdnnOh5HgtBoyrLbcVoWBq1ofVE8MdFZUxusuhMq4jXdl7+gBSVwW
tIiA8N6+Sxau/yzBNpB1ZAXoilwHMB7hf0ytUuAUy2itjapoRnq5e01g77yYk2Qd0hmkxVF/GH9m
7YnwrlzeAGxeVTU+sJ7HcOwfkuY98IvroQ2kenKEx/H7WsV/7NuERX/5aLpgp0EveZ5bectetPR9
8bjOzyqfGypG49DjGkWGsvTPbEM13kSMGG3KjAKfnDB7y6frITHuN5BWlWnTfkZ5uI5uwYg8RVo4
1qVW9+znb0Rpf7AGGu1As+5mP5OC8/nSbdsv16zzexV/4IWASBJkCWhbQE1BDr3s7cMdiDpeJEy1
vTZs5ciwyrQEV1dL3H8sXGG6DREjkUmbXyFViteQtCknnWToNJmkQUP1Pbw6u621lbtpxt8ZykIH
78Q1OMlwnSOALX/41E97YwbQ22X7on+cPi+5mqQxjf7X6s+bfwx4Dqxz4jRM1nGoDIlpKf6xm2qU
2WKGmESuVSyqJpr+nDw7vKERzEbNO27dQXJaicdZr0u4B7VpROwuAB6o1YeyK2nn9Turz6nj3Pyp
Qh7ArqXxzbeoogQWEF+sV3cC3BESq7WdLgNx/EmGPHWad7Fp5GeKFZaxk+EFxKVSOk2QuZdBeHKH
8ahQtsMdfQcZUmOfMrJXoXrmlo4MQ3zCyw3lueBqS8E1Vo9hntUpHzCMKkK0JieHNtr9IdW9NMjg
QrH4XvLHWuLwzCUnQb4aTyy4lBqSv70te1lLKJSpjGAt6H2w9g1OLp4EMd9calsEt5ZQgOds7T/0
rZGL1TZOvhu48x9x6eHK3rpZeG/0+/cOcOj1eNgZ1dHhMssJXlQb8Hw9Wv4Wj3SqiLqF+rkJt9Xr
SpyvxPDOEG6qsNgOQric6IVoL0qWGOg4HeRUDBCGk72s4psLC8gunsfjOdVfkJjsw/zALS0L7D5e
Y2OWcyn6aqiamXGSgEcHRotmSoE6vtCklBn+XwdTb6oVJ5KviHKIzYJ4k13vNje0he1mmxeEK20Y
spxFTfQ+HY72GXfe54EcKdqJTpKsfqLBYT+ewfXRNrLSXHseSNT1WB9rjik+pDddGUrkPo82honG
+lP5iE5RGyXv0hha5wd/i1euk3LChZzbNWDH1VsHmRrVbbCyGG9OTDQOnYFh0Op3eOF7ZionS4iR
nfARp9mmF1YDJMwt4Aj/hZWtsmftn17Ru66v3g8wOzs83aovBgmyota61oWd8Zf8iF+T2Nu+38iE
si9iMprqRid5Z/W+csOXU3n7Z5iRRVtTGhD2kH7PjxxILajtLKqUcWBOBdyvdxvc8PRtxrHKu1II
HF9bwgf0Bo0lHBJ5Q+WAqAfGBzCRpcP8BxNg+Glg1JGqhEsJJDB0fQgSKib4AguovJbd8nly8UH6
M23VdMuqj/EpNkmhGkmMpj5PUMm6rtpqmEzrjG5SW8rnrLk88ihMUhJQR93x+hBr3ByS7dg5FCGI
UPpeXWEJPb/bjykKl4aMvZ1X/JnwE/Epf7SHqgJ7B8Hhv3uXERdlun6lvqKzpuxAn/6EKgSQFLZJ
kxhMMyjKbMPHacjY/HvFCNLH3/C2UT/ZoqoYYNVwBQyAXL4AvXX2+SkzZW+OFHQnfG4bGTyUio/7
lcQ+GEr7yJ/zlt7hLI63SV9DRbhbVsUvX2i0c3gZBGV0YEwuIyOKnwZ6BbLv+i94+6FiMHSokgko
doV4qFn6cM9zw3gzs95sEsQb2qTpOg/8tic2dpFDVAXhw51lUSRNUmTa+bI2JJs7NPuIXqj9DTaC
Qr2Ox6PA5SEFbj//Uu9IMqj1En1g0DbzgXe+2QHnQCU4iSy85KYEgCBPnoZ1buxC0ARV16Scrd06
q/GzP0zGLUqYXUvnEe1syb9G0y1ZQLLNBopWT527LI/fwc/SWG5Ypjlzzg30RCrmTx866sgOjm2g
okq22G6nBtk3mSR4GC+bBbJ56HFuNCZ8x0ZiZcJJ/V1ErT0roxd8aAtiOXrMvnZl49yileqs+IL+
HBpHk2PPb0SIO8W+hUjMTsIaHbl8sZg3yIHNiT3pnVeek44LryE8cyKsDqtI+D05CqGkcEOoXb+f
gXI0/h6CRmGRYKM0h8C7NhLuZ3Pm/dOLkNBrVWv4zbjdXcdfxlgBJDWezF9JsTroFtqM9GI3CvmX
15CoUPII9hlCwy+FeMHlNHqF/EnVdH7SrPkBCTN86frmlagJukuhjqR6jld6RQFI6Xh5N+xKlEtB
ymOYnUFET6ov9dLvRAcw1/hwjCqDSuCbYo/XHCG94GX58Mj55NyI+5DHNp8XWcUlQCNioKqz+uya
OljZFL5MFls4/csjjHX9xOhvxoLkj6EYgcv41U4wVQEfXUA4eZQvyNW0YFikhN7ghMHXNqJCps6B
wkZ8EeqMYEAlqMt6FLaAVyIvwC7Prgg0/EJH6aDAY8t29/pJOCDeyxXGtRHWVFHBWntCJnG7L68Y
hmb+wzOOdCV8yEQcAaij8QkGVnBUizO9gcTNf/DT1y0UsbuWItn1mpROAk0VIw7soK14ubcagrWc
PtAcuLuZAO5n+N0A2ziYbtV8B4G1mWRKZThDyjn6KR54Lv2mBon3a30qRePhwwWMO5+ReIzy/sSX
uBHN5kaIqnOTtfXup2EGRJwgt6b9y9NMARqh54Z62spEGE/1J8pcXTM38LV2/ukhxJlcFffp7Sf1
XcP63LO+UUKBZojRsCyROY1tQp0sdeJvxZPunXjnYUhiytaLYNf6Blr3BRVV2JZ/oOuFxGseZq2H
SIOLBTjS1EZ6lLjyu+Dq50l5LfN0idePxRYLJ5e8D3fiBanjz/iTPgKBFhnVos0hMp5d6BRe6rb7
PVPbR/Vm6CfksvAIgIFMAOuYbtWX2E8+bh8KdcnyPevRW3tI5rYSosNZuvQ4w2aHGVu8SXHPMisF
WwmqRfF22Z7J0dtJwp+sjAtumhqGi59njBIXZ99oEd0UWNNE2Z6vQfKfaze8akWfe8Ksyp4ZiI1Y
nkoaLUN7G9GkJetH2wDaOIE1l3/Qwt4db1rrzm4h2vSEFX9Rrx/pdi090BiSWKu2wrSwm89g3TXq
OQCfhzB+W+Jbs4e+nu+DmyAzhoxK8ahCYz4M5K69r4pdir/0zunwWJxqZsFk2/1hfyBDiZbxBC35
TeyMszlJJ3okAYaZAIGCwr/LoKfunI9VS+lPB8NLd5qt5TS2pYNrjtNIyYShbdjaxMOtlsa+SvUf
DU6GxcgJZ7E6toN8dVAIIH0g6am57VRqqqKUy4/rqkItaTGXpGh5/TYkCJ4/35cXNgWu+n2Gravq
bEHGk6K047tWhcmUsmTk/gGYDP8ffWOB7FNxACBjH4rqv0jzzY1J4F3z95FmpWhTF0A9db6TBPS+
uYem4fzwWqL1HDZnQVToIEaHqS2a1dN506M0o+/47yi+Qn4b7cmkuJrCN7NmfhWr8QmLfIvEPCyP
WSo/lYiCuuthzB2S66O17nPQ6rguysi6WJ1qbPp2yPzmK8yVLM++x7B3GShap9Td1nWyo3oVfEtp
/cj0ZIuf585+6HiDi030M6FGlDM/G+Ni4h11+C9rgkDf4lsms2KuNXmkGB/e2Obl1Kfio+qQMpn/
OUzh0sT6hiHYP9vSp2IPihajCdXssWIMT9RA9McvvoM6bBqL2Z+LwoJFCUZrFyMtsd+Xa1NzdL1j
Ul3diWnmLdbE9r9MoVsHOI/ABnHNcfhKL5JtwjNDSO4tPFhMsWZ/+re0tWga3cssXHs1dIQyqbE5
pEjYJhHgKq3iHLejqelFVJpgiXY5of7ACvvibtDf6Qq8ou+e+7OHdRJpMVNdyickgDYcUO2f7+vf
DpjQdiBDYzbMF1TygErL0nZbj1d0mLjTn0nwwzJiJlhKR2fWsLe+BSu+lK5HIzLAvjBYyhVswpQT
6z1U8wBl48HtpO+KXMnJjtBkNRUw7gz9s7uMjjxtc0vBfsN1QDUt15swhcbjKvLcDY5AwDd0wamB
ByWbCHj9TaTlJaRbjvizgYr8+HATl32VwbcU7ZNurfXZACaLEuqHCotAGVw8fH8fUIIxbL10wqhn
3l5uvcQgjdOnLQC4c5+wTOrjQhGww3jsu85057e9ClF3W4vWH9aFKNm7yfTBU/XjryjFSmWYGn89
63pgMLV0UHMbYJDHPPBHBLMols3sGWb74Y/cUXYIa+9unANFUq8ih1jLXnBYM8lkxXB6CfGmizhe
W44OLmkDANqmJMD5GArKxH1MUwljmG99ZqJZ5VZ/oDwsKYHpFY6TRsgkzZuXvyqXE8ZGN5Ze5/1Z
td1dy3TczVQk0tlOiNwaqCi/9QRRvm7a1vFfbJcpENPE/QQY+r9haOSqHLd1D5UpLeegFxVDiZWJ
JN+wg71SeiYUr7gIil0XHlEEUKa41hdE0KYCi3u6kslEasnlaYRnhclYnAs5DePS7+QFgoIsJlMt
E/10UvrRy7X8xIxz5QRotyiXASaX5zXNn8doTgDE8M+GzMvlrq488gEUiUB74c+gcelPumCR0Qoy
hEgFeiWJOM+CP5MduwbPXq9gaaS8XjUvDRDQOeNl9NyrBWvqhMnpKjcJTH5zeilNcja2fnreiQRk
j6N9OkkvaWYYD0tPcXy0i0bvJVhtbjKvDGPj1mLBYRjfj9nlJOOrtZNBQx+VCqvWu4IoSPzYSkwg
cismdlO/hiCYXBb1PjhfhRDYKii6vh0EAOMVFw7XQ23v7kZ8h2fwgcRvDgT86Gs/LmnBE4YJZeYA
66ypMWobEopuhIsYB5h6OsxhhAxSpdDQQB49UTBP4FjGiW948sNevop/hEof3zgqeHpaF+bjytI2
8Vt6BS8AgC+fnF1MUFTvvJjQhq6KOfy4AooI47/NuRJfmUD4AZp9KXIksYGO353fHIjA+C6O1qUf
77l4cyxdmhmI7B495/rgWhKJfMUrL0cIgXtYE/tPdrBc5F4ynrgNGUcHhbsgJQa8x9pJdjPhT3Lu
hzbVsl4XSpL594fxFnk6KLP15o/LwWiZxxzeABiK8Vv6NR1idGRvUNuHD5IpekfUlYoNUTiUOvBP
fCyfi6ZDmeaL52jz89OWpghC/E80ZZpmg6v/q3OFo5c6nE88/9bxcAQsqtK5/qPkt1DMiD5w9fJL
aAr6Ui1Y/pzIgsGdfMtjbBkxNeAI4n5CPnAawdhC4zyuKQ03y22kZO0N2C26PGvFWtGe1X0/qPwx
7tHsI5CFqfIY3UdPPQWAd4eMi488+3y1eFLAuErEzyR4UbLFynVS1msoSLhyKrgqDJHUxAOsWros
9dQR2YrQO3MI+mBx/GY9MEZZiAi6LL1sKcz88apeMMtVdaKNkmuJ2OQdRoJVqME+y0X1XKq+dgqD
Ni4R6TSKStSYiE7W1/8hlxGrob/1aBBFjwScBbGGvLdBFMPftpfbAMTV1ED/NBX5ESde4I85yHMd
y9ekJ80lAd9XE/2eAP0WG/RsVdXPhrFM5WOn+9pPYShuJwuYjYj4dgSwhvJAA3nNt5xRFC4SXebH
T2Z8ZQDinSI/xuA2TKHIsEgH/45I9Q1UPmToS7F+65tkqv8KvHNDStnk49GPgh0Zq2jQAzynyjEy
ymHAAyOnjrsGkB0BtiK67/P0np1lTKUg5hozxUt+Uygu8jq1xnIMmFXvn/5ATMEPuQ8Tb0Ycq/47
24PjW2uM8F1eUWfGMRr1Du9/FnB4gp1TAkXVI1h3rB1HEaaKv0pI1akUxx4eEqG9GmCmTNHqRkdg
DeFUIYD63lOIWtFohjoYET+pMsgCq03Iu7k7I1K3U+zPex9tQuzX0Xx3bW+RavfSmnxH9cM19yI/
UN/2qkXqqu3LlYbvQgaJNtwAou2uFplA27Pj9e+noCO0lcax0TldHa7ZITK4kwhCpbtIjs/JlvTG
3j4i3AOgdufhSbSlIpK0D5rokIXP4gBPWcL9xgSmgr338QuLDOcNbsb2eFaNo9kHkXhzP3rhQoR+
I1nArSnWzwUTZwVaIm/+LW/re8+A2pVdG113oM5D3c30jhf2m75bCmUGGgHnDSQNt7t1LSG36CqJ
B6ki4WChpxBREvBihWb+kc14Mc0XIBJjpy2ZlyWmgizNmqKDRg/ClXq1FwcuXP2ChYY0yLH5hEbq
dvouMXErMBomXl35gV0YC1s8WV5LMx2ZS052TFC8v7ebFZUI9JVlBqgONEmYl4M8SwLnQ6Yi3Bl5
e9EqQWpFyjnkKYFnrPazlRypMRjFXuDTbZeptxdOlrfUrtf6/DBtbeNRSofdc8UHNOcmvd7plb5Q
A2AdmyOfNtl41doXeTj9FNCU0OClH/1w70DQMp2G8u+fkQ3K7CJpFFWY/KXltfRSZXIDF6CQ34Ex
214vld9dFtMsNlHnfR/ukOcUuleU8GHSthQAP8OaccUjI1b2wXD+TbPx8w36ydfEweYJ8mYlqs3c
Q592Fus/jKaBHNbNcRG05TqZZbnPpUGnBQGE1TdjleVh7quW92mfLkPkzd8ECltfvJl6/Bb+hFkT
k8LmCdPCsdJKRarEobUf6eODHL6KjYyvXXnaPhUE7Q1XjMBvnVyoY0JO+Z5VHVWC8eN5FhsBmPVW
9xRl3+copeOfancK60/Q+2CpVuTj8GRO/2wdmE08xDWrMBbzwl+NXwXlswQEGa9Y+MkZACzhP7sC
S4mganHWS37VgluFV1LHuaFE8Te+bXyjP5kCHu7lzgfzXyVAbKDn+N8mGexdFOhxN40H+j0trvaq
b+sBekZWluw8laJi6+/3k0EUCY/9EYhwI+2Zf+zHzgKv9CG5jV1EEcg4vnp0tRsCvavbWY/dU/0r
tWIcgPAcno3PW5oFFcKBYntK5YG2IJmdp4r/QOyc2D9wvmSV3ND1GKNAnKYqXDDz7wdsZRb0TSsL
4o4K7ly9E6JH7m4JIuB9Z6GTt5cxMUdMsxSUEK5aIV2kLuclcgGQJDzg17x745eaknLv4YpCS605
M/PioIVNxTdOqRL5ZR5kZOEY1huAjYfTz7bbRgSCUxZddXlFek20Tjh47WSovxBuFWUQbhjhq9oz
Vb3JNsyKucgotg/gvCHJ+p5h6EalRDTPKvukza+7ACPPoqEM2YJ5HixpklCbYq8Ti5TB5Pa7glr8
ggd6lsVfbOu++96ap42S3vuO1JRaBa1F8vpUwgCSeHDWrmHC0GlceB8O0VFds2upZPs05JQhcWTz
P4SVHCfKPj+IMgo9Hy8zyScsCwGNaSzfOM2Rf2DWrsCekJOLpRBn8e43Zf/iobpFuRdkng0RCyhL
XZ40r7sbCq24/r+8syHBlwYkokayYqSGRFkKcc4T95cYN3KnJBzQ0njTkymZOWSTcjgjX60PF1Ih
CeiDcvlyXfoEvRMZ3UEHZ7qSAcnPXkMgKRxAofhS++LCoTD2wVe4MliIRfU4gCHYAoWVyBM+k+95
RQvVyQWsaRFEMhadaRrV/TBNQSwfCfK55vIb+obuqGYEz4DrjqnasBEiN6mo5PdXqQ5n7idGk3EQ
HkNLPTxCFYsziRXE/QzolIIhd0DYJ1xvGpbQZAABy44tWUd/KtsyW/mUJfsQitoqi9hdg54jp/K/
7iI17VKVYCSClf9Fy7VE6sw6FFeOOpEnWtD9kTjPLvO703nzlVlQmnrI72E/71hWtgIOKiRE6ZY1
WbjXlbMci4W4YmPqwGEVuOl7yRTgbDV1lTP0LOW75rtRD9+9ibk9ijJyh2Gt4sm2dwENQNf4OfTl
yUA7YJDr4a57EGIX75Yzg9q8C/tLuP1KOgpG7gEml+jljW0TV+5A8Rknuo05I2s9eFTEQ9EFpl5c
LLQjbwZD5z3FgSlRS7yjRLzw8EB6KhbjbqnZbFTqyqeKafJL6bC+PMkCF0rNZt6PMkeGCbeeeSE3
7nNfDehuL/XAbyY+ligQwx4sc+Yzr9298Swts1xAU4L1p5pys6rPIWFzCxcY61XzDeiMI00GXfDd
6EWpkNJrqC879tmjJ+3P76rnHQeNFF5lGN6WFvvEbEJZCGArLn1V4kKZFSsA74G6qaOA84XhyaTc
0vT5itQCmb/MLVuev3MkUqcU/WFLmrjvH9nj4ySFJLC9BJl22hn+j/1i0tOjkhACuOrPLpKTaKpT
AMmAww5rpgbJpCk2Vy+7PCdjUAU8KXqdmBn/eDMKqlLqKjZ3Nm+nWG0S2LBA4ggps2ll4JEXPCKf
iEHH6wzmATKnVa/E1ocSTEGJkTijOskLsvKv/djjlQudR+KVfNYZXi2TqqBekrPVwmPlccDyVS1n
LuCB6z6cI1TRzwneEWUL8isiVKB/J79Rz/LM5tchr7oUNJ40bavGs9jVWDKCg33DLfvET4NheKbp
v7BDdQnDqiD5ycMcI3I7BeAR4dZmdOo5PH42+5XJOgjQj9k+U9+0p9CxmC6JNktODuOZi0/mdrwi
8q4B5NOytY9VIIAul+YYe1okAJbGE73MhkUZLe/ccZvLBDQ8MvQNJXZN410KZK/qMIgWvcHzhjOJ
CpFHEUoHXrOkbSsimdb7s0zcsEGS3WbKg30KZZGUpnohe1Ed7CSR+xJjdNvtJ24Zy56BJs/zF3VB
Q3m1G5uSp+rBDq16tEP4cvpxR/shMvxkXoKx/DeTRAykf3uEEXCH6mw2jUhOWkuYkCXLXxkQoV8O
aHkMGfaFKwb5ndmfmw1ejOIHbD0orXckge9Ko2KSt2i5dJ9GhhHKrBGJQlN+im0zZ2/dzlrTvDHE
2FIH2pN43tF2XPYOvyvGJEM5hpmq/X+giJmVnzlYuJ/uFrqPJNxRAEjpJL+42F2MdMPJqsPuzDUw
On0G3Q7zs6tzpY31qUhNZG+Y1vJoV4uLnOY5iJN5sEgtx3wCyHWITXTlQDXNynSanR6pI3E9UI/s
xyYGkaM4DJOXqCb1hmA0czVv1/3I1n4Nqu5mOLlttry4AcNWGbg2UaraEXBlSE1qVXcFya0Ytzx3
bmw9LD9xlLQJQUQkJM1xDqFVTLZdntcik32vo7Khi2/+vhBhl7no5kY2Hiarp2yR1EFDGrg+jr3p
WgRN12YGc1SY6adZhtotQ2lThyTZf9SdpehfYlgeciF4j9q8WOtfd6Ps5YdehVuAXmH8ijwasgyc
f9/hgV4kFx2oeGuTPVzHZcAFsNbovy0XxVs05HE/juIv7p8+45JzTrJuQP7WHzr7ztIiUhIgm7y1
cNQ2Wpok2DF6/1F9hbHnjTKeMGH8JqnkH7Ei2onze2+RH5zsFWfzg17dhfziMBXYwRTXqT5AIOa9
da9/92nBdIFGSE81/jby3ts87/F90KZh2LDY2QFShBFdkF5lxLMMi65HlRrXlvOi1aZUz/Qf51lk
/Mb/h7cVdsCuonxFQDIo3/WGhKRgfcCo+SGPUObrmYn8Rvs1Y1LxxetUK/XvDwYSZgfxporetUxR
E4s1AA8h3H+v81fCY6LPnJtcwEATw4gSwRHokts9y1oDKatSDRYAc2N3NxHprXkxBPjFeyHgYI4h
K6qtWSZ3sMzNYILt6gJ5Ou7BKpAPCbJACYIfM39cyeJakDMWtWEAF/OzpqF0euvvLnuqeyNBczZr
5+uWoQ+JpnXJBoDszeuLt6LP3e815aEzvVmyj5fwMdcc5rXrLo7JFCbnhEy7uUHlu86l1wO35LR4
1LgfnzYva/GyGnjF9Dg+Ma6KC4f+0DXqXt0uZzjg8BFU9WiHG2krNpAcUyfT2ot+CoHBUIetg3VP
AtJS4+bTAjB5n7JyCaHzkvo2t0Zcq7Ms1yxDfCcLDDtXqqfrFrUh0qHyCurV9j9Fm4Z+88qIoJda
icJ58o5FMIihFHUAlyXB7x70BvMB333dTUm/6PX5ZNUl6eqNFtTJA7+CfcIisRWJPI4nJZbs3N3z
NnoOpbKBQqeuf+s4vztz0ZPr7pMSWlo7TVYLhqLdLFjGMDFSJOIw2mztBzHuGzQQCAxPAtaHLjb8
S9AvwiY1JtJHQnUcgECmdizI5WPLGcnlc3u6eZ3twesmzsGywV8gVLTAT6Ul+0SmfZ/Fx3UOfXlF
mz1qbSjDDMh3DaifBXPqymWJPKzzECMo6jDHVyNo4pvayzx1kXyKgHksvyk0wzKu1wxawnBcCr88
eu4vqmCu5ScCp2zCRdw4kz4Rd3hRhvvXYlIMpu4XywLgyrmKh15JqRHuQIGXjqGJYRXtpZ6wyZVp
sb2Cjl4DCXWeLWROUPXazcKdLxvU+xVQJXLuv8AlfQFXR3WyheHmtzSuh/xGFr+NplElejX0TEFQ
B8qqWbOwnb5zXqLwfUuTW0djZRaK27jmuWS+DdhBm8KWnSTd5L3VqHD8J5qTgkkOF288XktyUHxG
2k0tB14H9jqYuezJJuC6PEZuKjnScAd1GP5iGna1P8T0mqzmeMqb57hVdMZ/opYO6Oejn5iVIXB1
EBrsXwi+mt1yWnmWB7hKVtkPHd98gAVHGvA446HUXQ3vShcoCQBiocfsCRV0Dti8fwsPfLL1Cfcd
3QCopymzayzmvo3qXDdkPjqsVF70/2ukJYJZh9yUass5Xee60Gd2oZmPfIdvBtC3S/5fQx6Jh6jN
iVoRwLydRs7g4mnZgxtnsTZ9/SaJsnAMvGJuHDVkFDIzEljatWsFnedtPSjwwc7YeHFIICHO+T6L
fJkJrw7Ll36eDbQTCPZzdE/sRycQcjnbEE/joNBi1rZDFxw+QM8n76Cv7RmdOgUgbn26i7vgnia3
VxlhVAo/NA/s980OSlftx1huimBYD01O2nmsqz8QiG7ovGzbq/HbjjCU49cmliKONr9mGWIVPXby
ut0tGNZf+5xtN+VpTDjIe0N5EcDPVeWpp3c8a/jmPNfu0vtycY9dKCyNwQZEa7GaUHcWDPDdM3NK
/m4zqW3GOtqHRp2b4pdYfubsqktMFr5QGl6FOe1wHzcWkdYz/OGeN7P8VZJxHACaf305/KO6bzW/
OepADrfVe1ksUQCav/p3t/06DYOyd0pqGR2kkkvhHQNA4UOPcqTg4UV0zdj6OF0z9I25nUPW7tix
k7D1agvPHKRatVn4Upz/IcxCou+ZC2SE8EAaEGUohSY7zLrwbZm8mNHL3fx5etBx9S9Yqp9DjGOE
/u3p5dys606RDo/+guQYW5soXfj8+VczBc0B2mp/qCWtj+PFWG07b2uMctE/FTk38aMgBCj4cyWQ
LGoujX9Rvy7lDLIhOIQqocd0pG61E/UP9D3Ok1NHijVZpVhYxMBsHPjw1CKy5bYjz8gr72Q0actD
l7/+r8MHk+7z3ORP51sdm3ITCn3dcvkyQJFYinTn4HFqU+I3V7EjjAlk66IROuUQKE9syAjLufSA
j1BoBiusZrmnccO0YorI25QN/V5nv/zfeCUzSMPi/HJ++6TRW3wpnq9VLny9+E8BYyDOerebvj+m
xJ0qf1oCLr5RaUj91LbQ21gCQb+rysYoMUG8oN5EBPC6b7sZctnZ0wGTK+FcnxvHDb99DKiOANHg
+qGodjvSSvA233myhzwkZk1ks8KJ/Lbu0r1tBcc/AfY7igaNrDobp6SRkzIKCH6MkO1FaZoC7uAr
SOCat4Juh2UdjfuTSc7QvL6tqcUpFOTgWbts1pqKwRv3MefUiNXlz4Mn+X++LzzQ8o32Gpy1SIyd
4PXvYQZpMsCEb0gxqLIZNi/96BoHM8es/M3vT61SKaD7ilMT0krRAN328kdVd5QYPv/RppfJQn/5
PG9FWUKh47ahtwZx/oRIEeBm8wjaJT/R6BbmGDccYBAwmiiR9atU9hnOKkq4lpYF8NEszXtA8PQO
x6fQOOCAN5wbfOfVWtYlWsK4dcVdWNDvMQA3YnAST9O7UjnYFh7zHBHGApCeAFxmTFz6PwM9Kqku
ml0594PcuN453QzFXTS7m0Bop7Sibcn5WiHwh2upFnF3ekiACShh2oRqqQqy/IZap2/YIcQrReJ/
kJDKD6flV9M3kO+AEtkF749AMvKt+uNqdLU8DYUyMyIlvCXDjJnl2DcD1uEthwxOMiaCw57ZS4RO
9RC39NU0jyzZiqzHVDPaCNKTEf8kVy2V0odZpjXKhrb5IWYirEz8i92HlSKwRNxuDgVIb6xBNm5Q
llEtpVBsxJSVMg1Uspp14L++7wrpoPQoul44yuANSKU0phnH6apD9+faRkoTBpiaPGHhPeH0p3Dv
RVbewSHJ+HOutyGnOG6Yx8DTSbBKyl/SLAClzj+N86XorMi+Kf7IjIY1cWsPzfMReUktygX5lQPy
hmdDKcD89ODJ3Ok5CQ1hIkX8R5B7QPJ65itjxrge1CvbTdROqIZZxDwKq3Hxl+kj7+5WDlLREqP1
CSVLp1Fj7vnBkV7MoccKgQhBCG4thcIEo0IStAVDUUj27MVhP+557bdlWKx8/l2idtxamhhrUqZM
vzMisbiw1cI/GQCecbDSDg2c7zPdb5omGf1Bzq4CZY/Eas3wb4C8v7KlfVP4WJv36//u1fAUpazY
KewsCsgkLMrU1u8pwN6sYvRtWhWRAR0IZ3yJh1wZodID2w4Xuwm+utK+jgfHj34PK7CbmL5uXa6P
0971MmunfdlH21wCQ0GptjHNmhbM9PVUCRm4dT9GevwURQVy2afoQcv3R9VRvCbmTg3hA1PAeoBm
aYc3elC8pghCgBT+jlQvPS7wPqcK4fNM41ElFqqrlC/jYMXMrQjJdHcRqMi6bImC/DwZnrfd528b
xh8RJHtfJIhsyXkzhXDYf1wnSm9/seNTdQW/s5mYHMvkgY0Ct40p8LmTyPnMTZ6W1QLwIPFqQap4
Ef1RtuzqNVadE0XlMzXFodInFO8ohWctuO5wLQEHPWCXJef5g8vdB2egVJgj5T4CYd8GN3akkuyy
Xe60OtdXteO/xIx/8t+tbSVK5XN/ta+MD3uCJvBam3poDhHWEL3uvMF2y4lDZnbxafVaUqo90THY
WzxPGhaac7V9EMtiDPtcRhPRSQoPx5OnVly34T2oSLjIH1hNTosRIBhyIalLK5ELGddUIcx8yeHt
XeCGgZh9h2tlfxNFtLN8IixsF8Zib9IXCu7/c/ihaDIkEt6EUnOn/oj/la6sSdYkXWUlMmELybT9
VmSgj7l5XMFhkkCZH7exb0tyx5LfQd9C3VBCAE8gffUmtdbQTKlIvjXRcBfjdleXqhdMcLutTiiB
lItjBu7vcbI0rikpdFUEvBDupvu+xheqtYUkvClTL3Ux+w1XsCl/iJRQ51imZNW0qP3AspJg3zsa
vCU/5yOKbknhKf4DHVTrKQqJsGWj028zpf/+TKeoyRS1Vjoi4y/hwmSmFy2cJI2a0CKQun6WDRlf
0hpcQWZdR5jlQAkhNFeSlabMper9bsJgTXqs4tsARQLo4+WcuKebS2c/rtKRCMuxu8k4vB+p5nVy
ad/Eyf4BEpce0p54ZPaDILD6E9fGi9nQmxC67N1mjU8AhfWrNU2NpnqoXRWvbyNwI4zEMT7CsV0A
ASKNlLp5nBfDKzU41hO12B0HuuHS6E3NYqwRV0YjAzpN6t2uIueLL87UIIiNAzrh/nEzbL6ZqBD9
wv+K3fmg7QWCdkxum/x29khvD1MjPWrlnGLOBcmT3ozXtXVz8TgDG6Du9IGFRFbVYzcPpBya/Cfk
QJlYF2DW9J7ey9F1Pa8//MS4kzYAbEgcYhl/V2JgxloWjIesmM5V4DTpZEYNUvxiXk+OomVMOURW
kvmfjsJZFp3QaeSabXGRfMFxHY85Vk/dXUUcn8IbGWuVkpu5K7DIUo9IsCuSNyChaUevkI32lK/P
8O4QDBYatqij96wFf9k42O5P4f5DfNwqirkZzrKTkaRZYccXUArS5ZkKeEtYRUrRutT8RPPIY1b0
9ZMSPjF+dnYScq7BfkjDzhn/cS+vX+6vvtsWHrsnDjWrtXjPNJVOPl6OqxZqkzbRNRKDMq1fPG1R
0wEK+S8Hi3bYSjYZedYRJ8NPzVuYE26ZFadqKG5GcCBJxDe8vi7/NIBJB6/XOTeCklSKEtAxbp4d
hVjDMX3o+2WSi9Z+qaB3+KHUcQfzGl9OmueQ73hiifTCWLhkskGi8IpehnhUblNAygd4D+h3vaDl
77otYhQg4+wAWrTjPeSDv8mHsrz+ZOMXkgFqGf/cWY0NjURK3BxKhbGJfsdrIxdtlc++ICFAFE0Y
L+bLThcMlhVMaKuE/hlghw+6aQzcF9a1c5+j3UkdEqFZ+WzSj8JzmAiNavc4ky+52RqrO+pL3wwQ
YOzZaqgLiL7P1HF8kMq4po3iWyc174qYcDq4uvKagElq8zn2JGqG1mhJ3XNr05NbQ8McpStBePjS
276rmCLb3Y2OgY1PlFey+jXkMttt1GVPxpWCQ19UbplQ9SlurfKlThwmo2UIjFfFVfK50tapJ4S/
WLJnFr0loM4ef6mvNHiKp/V+XL2Yvl/cHO5NCPwqnOOG2Ii41L1fqCNVHgUthtplNdJ8tlJSX/IQ
p1ZlvmJucR+3b3mCMTg408cdWql952/h7ZMM+aRcCQ52n9vfiLaSjfipHco8em/rwyhNLAbWg9ne
XVKNxhOUEiRCeB+EXu429b8pJmC3vm+gNBACQL2KbVUOTLZf5OyR6zJII6FpV+j0ncM5Ju5zqgqm
BmEpBbKIamQApu8mUC49giyE2wp0Wq4itoA9/37z+gBD4qoTAg6aOm7OfTw6f1TufTyxHWu7Bpgv
NeiRf53e3SCNfDFl0ED7Asg7QOgt7KTicwBDM2gS0jIJhXR04Tiq6Ok+DpCAwyS8Ss0AbUEjgUd+
S8I5+ffKNQlxguGu0xziYKsyfEWc6NHC8IlcAPgL1p5BIX/4PbcgerWc/FpcmMpeRFRkQxcQK+U4
ncCfbTSLIFizEo8qxuDecvXW5Xd6iL11b9zkCEgayS/Qr2bobpzxO0hRKY1C8aJ4QFRlPpo3sFyd
sB/PEYDT5mc2yh0xePwB9PEaNOFH4dt1u+ou1BhrzV0SAoAyI19YlL4igln26KwK9p2JTOHjUQQ8
GOVlhZI6kkTQ87BtgRtG/vnuPqFw9zHrO3JUvtj4igbi+bJ0l2aQeHhnqmrIH4AgRvFkocQ6jKDa
rWZvj4HRgg8ryU9BQlVnkfkEE54bPiVizklgXt3otHwsiZl02hr3v/BNhvCLWXCE8XCdCCUG8DmG
IJlo7OM9iKForqUG+NnR+P6ID9/uQdzZrGz4n7UkodFlpL+qwBQZAXzZr1wC0XdCiJ0/8KVyh6jT
iMftk+cI9ZZHwBLujDr7qB5mhQixE5yQLNitJZtwt67NTuF0owNbEIvokhOtBp9dFmOUHZLTVEZS
U5Xn1rUbqQYL7HQJLwklaCCyh9ZgfjaGdJ4A5btfW1SaSd2ZBzYXagA8+WrkLcynpJo1XFEG9xNU
U+H84jilmdD0ZRNWle5jcHElYeOu1tI5di19pTaj/+4i1nkiowtoorVtyJAEZ9kVJPvOGeWN2M5U
hwItwi0ObgZWGCwaBUJaPBiC7B+SslbZ0B+UxxnhA6zLYn7bU+g96llNlpZdGqi156ewqaJrgbBl
P7gFNVhrmkbA/TmiE/KRMBNUGpllxMj5d/mHTJzCctzMnuLM+o9vl8yGqXvaH1Q7gNwgdtMFPN9C
tfSQltlFlT3TsPGtqQDEFqfYLk6vHz3hfGRi8bw35DDnNTM8At63Oohni7ytzOVHgOxCKNhGhWdT
aY5JdAT4YBhRkshbJ+OBSclHf0yQLLr0woSm/s1kScqmnYFcEZyB9o1w0wt6Z/jQlSI1hlHy7y/1
tqsieiYQG0+cqwmh9ZfrNfSvqX6r+6HVMgi3M/ys188YqRQr00eUt8LqsagF+UrdCuvq6Dxf8/7i
UCRGAr41x4F97NCgl6d3TslzZXQz2odEIVFEhpXgxK5aWC8ZuWmrxzua5vv6OlKpZe34HYRJbpMZ
re0hOj41/pVKq/oSTV9Yyu9Gl7HJqCxAY02GuD2sEzMBkRlVqVX8VvA4+VXECfn9LE0A/lzr1pR1
vGasVKuAf2Uvu1mV4ndmC2Q2ce9w3aO9XwV00TncbIEITDuqvw6YV9DY24qhMziRdsXrCBJ72SHD
60/cyiGt8Vyl+4IpE3x2x6ZLXeHylP3GA0ffI27FdvU7P/tQ6Yo55smpUAX16ZwincEY7hOsbjlY
epbNzQ5Te9s/hus/jmgn7BtDTdbbvbRAHZf3wPZjuAgONYDJOwNSvewtKgtlGt9X0fJZsYAF9NRQ
Ejv9TuaFRjlSIL+zn9orbiU+KZkgFoXNeqwTzJ/KGyW8e5RoEVr2S0yvhLOfn+oCqrXTHSjAoxkD
/xDMB7tCvLuMAOV6lgkcZKliecfpkEiTCpx818bSaO0c9bQ+4zu4eOfUDQG6TVOZQRwZfoZgXAx3
7QsWt+ab1hOHdGUqkJ+fiVHJWTiS9rxm3u3yYJxuF2TcVffEN8I9Ris5SjipvxMA7Gbv9lc2QsQX
0ODgxYyAH66fvCf0SE+AlC5+tyIP0Iw7Mbu04FoQG0nZa76eLWgumgk7BNpTM04DFb5IlgPiylSg
najM1hwo1hlSyLVJefmCNmy8ADRVSkf/xEESBJCs06c3mEnX35Kjh8p9q7lLJmGkja4Ozk37hOBX
r1/znGnAsmBj3m78mqpJgrtxMf8PpUv0+I8a3THVgno5OOl4BSnIeuTkBBjE4qrT2760irJb3nv2
E9HkhHn2nFZnMkv4diOft/da+s08i4TCa+esgQCPlMR3UQc2kaRx0QVFgIfPpfEeKTKdjMdinKvK
1xBFPiQXBe3IxJyrprhzO9n022TfXU5z6hvtqzrJW123Gzs1keQOUFjbvcBfcq5EgO80CfX3zDdS
+6FJm0YW7GAddS/hGDgs5TVaZ6orAnM/m3YUPyIxn9SEa4ocNCaXblD8H9XX96qWN9WPz/5KVFsV
IL4JlBvKhQTZ1p819gKRjjZnWJNDeBxYdZAoLkh3ZUmVwqHdZDbxArnnhkft7UmOeeKIczXBX/Kv
czkrM0Z4ha5CPNjqrx64Es0vcBodREDHhH7c5jYkn5Qp/5APFu43KDKi4rJsKWO4Wemr2Y0/4hhf
wDgpu8RspECTOABV+ZjdveXnEk5cc6Jdi1PjVrHcZdKL8sUCB3lLQCUl4+sETYIJEZpp2y1NTtoq
4TPNyGdaXIXL1WA9V5yZXLryEvDG6GfXsEy9cqni8kcIULESHn7d6Hjf3FSN81XrSQ0ksBvo/J6c
4OeKc7AbMSjjaD0HPvKXQl2zSK0E5o22f3TYPjRRQpI7m8jiFDlCYe6V7V6xB7y8G0+oqsRZRHTa
YrfCXmshGjc/OQO4FL4fL0eh+vmbTjtM4TFcZapxnwu65q4R0rcrqk64fczKEBpJ/SYV8EnG3Zx+
aJfEtO+MFyxmU6jg32aCACJ214JyCIqUAXjzOQqkY1DB1eGHmOTTwrELPhGxDmIBGJxHhF5beR0D
3ujkB2CDIIqdCGuyRXn8OP85ZgA8ue9l7l4TTb0N1PXadsgKOYsKA9o+/JumsReNJ3oMAMy+8T1+
E4xt1y49uZTDUUuQ5ABgolQVkOwDp2xLg9fc6RQ+YNpFJ8IBiwvGCRcgZZ1+eFsOr9U0iGvcYdjK
sjK92ix5FeG0TH6qyKaAKn7eAXUhu488/a/+9cA/qh0TEQUQ1ef/PceaASuGQaBJJPG7gX47d9UV
WHmD9VLn7PFVz4Zhv1qQdqy4M2g0vuAzlTUFMTlL9c0VRbWmNzBfqE8i7ZFaVuRNux16kuZP7Mhc
0JjAkHsMtVPnMTRePxxNa8EfL5C7F7Joia0SFx8UhfEl6VfCj6ndKrnPsM8Q2V9PkqE8oilsWix9
MWlxCAKYazHaGg9mx1rKTltoycfDh1vB+yi2mLe++cRNMdL3Nlh3WOl8xcsCQKfhrdtm29fToK5V
aRQ1IBe+/PbCF8Nj1KzQm2XaCDrljnEi5QgQ1Ha1lrOcCRrMI0fdjzyXLd9lcNWzF7KAn9GzR5Yl
7dlxZ9kUmmrw881hw58RhIARIrISDaowcOBsVKQARohAyEGXqsSxQki6VshRtB2hUbZ7O1YIc6ik
ltDmjWgrdRCEjXmc8Sy650GXblyy0JdnMTIsZGu2/KSpjQ+57kpoEHQvBXvcWl/aQKs1epo0zatW
96+nWtBpgAT7nUgTdYr6DOjIJ/aGf4a4JgJRg9DR1ehQLziMYkH6lshiNfLyBeplXnlljGAI+MWW
SiEVr5uPs4ggh20UqE1kSCkTUwQ8J3MUnkUhhY00hXtJwbKDsW3ADbyh4rydu/cMaMfahg3+o9wf
vXl5BIaDfF2H7q0YM1CdwtG8tzDtp/HpbtXrXcf9HkWgOx7DbWgXU1sKv15iTzvPtKkJFE7PQz2l
VXuxU7bxwd6TJ1n847xJ6ZFrct9FJAQh+jvR4JXfg7EQPXSeknxM4exT5p9kgwP76MUs7UJUob2b
yJbK/p4jLJVAsYN7lpZwuUvvJ2nSo5UIpIG4VjnB7kpk+lnmobDL1PBydh+C6C2sfn7wYO0aohT6
MfNu7UvbVAgBvQY92M4539fAX2pi723WIHZEbPhjBtKjDxtz46pQOop/Gs592nd3rxzMZoP3HC2a
bdVuHnYsLXt5s3lpEWaFyIGZFFpvJBzQ1seV6jtZa6KFCvIZvA4ajcy1IGQSxmFyVv7JKXQcTqqs
gqGOKqrrIsXEp7S0uepvVtRSmYSoKIvYBSnT5QwWKLvvqoHM+H1IizqQS/mdfwHp/QLGRTRWlvL8
V18cXWzWeSpGw/YvKAanJsfy+2nTrc7NaGcnAbcB7JWMquNpdkJqvLvvplN/P4vNqgkew/34MiC/
Fwp5xPbkBgsKROXaSQ7sWpibwGm2i007Vbw7ePTL8IdYsQmYoSJzF4fxzmgUcvUP4py0VNWxww8I
nUKzSspz+h+HJX031ZdAEYFnVf+IpwOclBXk0yJqPJByBoS67SVADh0G5a7DbKh6A0twZ3OhOUOc
4KneRy3Vdbfz21ve/GS/qwGIcwNhukaI3rPCFQNIbkgWwytqca8gUSwlITWJeVZoY8gOpXrDB30w
jHnJ7acbmEf6rquv7fovhBsLkeQslCnvyenInOwYK6ax7FCDA6Vn6eSEO5K6tiwu064rI3OErnDo
s7nIbNMki1howHgd0TcBR/JwmoqKcxd/GlBU42trCq+UUMQUYcYw1fzdO3tAQBORzVqw8WKHyLvf
QBI2dpwdCmS+W7r9cL6iz5XzxqpliAMrTtrXqvKkPl7Uo8Gz6D4v5qXe0fvOwPE78UGbeq07bjjy
5xE/5HCFtVpymIEz4LnygUPeWCgxtjlIC3+6lmojwAPDXIeZfnBi+YuqAX8mNNVgcNb+7RwPCnyY
sYwzv7xDzq+r0GHLs0jfS+FYsTZy8tv/AK9fzzcOWLvwR2zNWWDvLUBlyGqgGf3+Yw0NO6MpK6h6
1sl2t4/+L0RyKtZPl8wGCR3c2ldDEw92X7GXlLoah4pBd2j8iLhoGSYyr43m5g4+ObJT/Je1Ww6V
2U9MTzalBj8L1EhFztbld1jQ+lvhV1KF4OuZ7+NdJifQwRnDUfSBXsbwJzMtgcnTQe16zYoxo5hV
AXrgDVPbe9tw60HV6Oi5YTzu+P3DkzXXOkuFy5+H1nSZjJvGmSrdt0vGYDk9TgPVNP8AhjNgwYfB
XhKOpB9X6wnH3TpUn1kmKdtCisndkDRZVZvICIJXoW7wKv+q6t5Bu+QKKwrllwYzUHo/l73tpqxS
8bJMXubrUNZeHn7kRnDZm8AyS/m0odD3VneBQiZ4qUDo4MTaGlXxDiOAxbdUVJ6dp2rpOMuHvkvo
ehdtlInNu0m93s6ZZZig2n/fzjt61BGl2rQCfwI4sVBF/aISzu9xJKwbHUPr4oCyJqA4ySpPbg/j
FomdK+ZPhEV78Uets/QVmZdiU4nMfo/GKho17bnf0Xb4g49Z73s3aWNbeQqaDEj7gyiB0+Qo/mRi
m6IlUde5LnuQIyjomNqhI7QzTwcsBAxvcSMw+Ccd4tL0uLzdLqQ8wbDia08ZgDOlp0ylJkr7qV1l
enMI4gtDgjAswXVIHnkjuHFdRrF8nPfUpoDmXbwr9lXnQo3qOe5whLPAabOhG+0vQuSs1c0xJKEM
rbkPswp9cilyfOHtZd4j28/Nj9VkHEMsGzuOzMUmzvwuJ2+HiL2v7AogLnl5vCHovt6oAwvFVzLq
NBgakQgB1Ur3ZwlkcXnXQBAbejhHVLndQT+m62c4iBK2Wo2+qmS2CfnK9WhJFQuQDg0eO+ONghKO
lH61lh+kV+Ve5jbk/1RkyBLi9MeQ0Ohda2FekrHghQMhyaxufVHI4bsliW20/aZGpkYeiZCn60q1
GGgdwSnaOZB/dyVOONDl7aCuWE2NIZOla3rZilqJ+xFOrVAavpVdVxQCCtqTj8Zom8y0J4g444Sn
8s/HTDTjoeItlktY0hmIQdnJbDr1TxSZ0GvDCDvKRDaScYowyoYr6YB1WxaFF4YcnxQVX+7NtR8D
/Cja07F/91reKti89YLaKwEkzWRFs/2EAk4eJIYv4ZYW5q2Fn3tbyimD5z1gYGy3eXD+1HAEp94U
hjB50cAHvdLhu9C/eojJWLG0Xgwld7bLnb5x8apCnpDeEp4rvayP7W4Zr5IHt5NQDhUytnPuclZp
NRXEIsB8fzKkiBrt/qTaejOno775lxjJnkICZzFH9hoVZRh5N8tMequ6+TdSdLXzDD4NiLCLxAZh
IescO3SpgZY1KGqbbHLnIFXJQi/+DNoDqMxo9Wrkd8KzqcOLbVmf+FVMZkrMkVsqCqtHFLZb3SJ6
/caqTmUUbYHMq3J0QoJJXzNmzdhFQpCPlbK259jW+qjqPs/DIc2aNhKodAQwqxaiV7KNiswp0og/
Ij5DtGaPobkE/QNDCgbQQd4y6DOmfNGrllNb0C31hPUHC27u57ogirjDeEmCzXMI9vSYMafPgBnp
xekWWjZiPsUWFQgpxTCRsAhsaOKiUSMms1DlOsmfy0bkVvSSUDTPSFn5+oqceAAAC9dGw/F3oU2/
UkhD0YhzOyILpdSPfNTceq7oVzbgmpo49XESbUTFij5Bx4+r3b7DlQ8RAzCam/JRBMmfNcdtX9mw
2aMS6ve0ar+vsyaT9Yzidp+9A6HB7HPFpMkjraX8YInN8XLlQN62eJufThyXFfqsjLgTC8BEEint
sgeHZdlBNgLCL0SkIdO6nIwUtNK+/MceMcBckFWzugCsU3GXorktLiPGYM38g85P5bwvRy0sUWmk
qmOBb/K4v7ZC7t4Hq5hqd4wuZTjElD907N3MvKhOucLM3tsYn+2ZHFQUramU/OiXS1DQhpxbNKkF
S/lqN3HHR9H+o4zJXTShwteUvB0B3nYV4Brybapub0cxcG9oZd3EX6nXm3Rq9qGInRDjMuwNBbe9
mzH4QhOBwIS4okn+t4CDnKzGNMmw6TuvixfNtTv4ovj6MSB6LC06I5kkP+6FC8itGN49+Ge6uiQe
JPiSAkeVJFI4wHpE7uWx1j5IJxNzXVxvZYeQXf5PRsqKaBZ3BcglVT8M7/JI4OhX7pHIfU/ui7PT
217M+jfvMgEjMI8qWSIo2/B2jC4GSksCKIgzVXbovD/fdf2oPoUjDE75PfT3w6muZZ2jJPY3ZjpL
/nzsEdIr2pBvuSkiLqRcX5oA3s6zCqJ2NbpBQH8LtgpYs2XZmfz74mj0Eg7k7TBtjpAfWMceki4O
moC8bG3cF4m5f/yrn9nuEF1SRNJtzO42O+BEzVq6/4oUdzNTZHuac5VbTp2HBeBXgD3UR4dOOI50
V5nFqEwQMF8+FBmUCiPQ9PobR/F9O+Zv/IstCcW+u6eERx9c0x5mGVEgFBSYZW3/gFujKe8oJaUq
J9WtGHlxJx0K2PXOBXUl2P4Y+NSWsbVO7QqineRCbxpA76QAghQ17juQVnvk6Xqq6X+6i0Ykk74T
LkJA8xImZUaxYEF7s6+C+BjQNja4DQqRjXBJky2aAcz8ZSioiLhra8c2+QIwNCPWqD0zdK6A+EZv
0G+y5D9XiIt98L8WVcEQe24zFmKvO8yw6/CqkU3FGDv2N2eEGU6lt1nnJrzhhk6+ZAPn0nEnjsrA
3aF2qilvBYhKHsWjJYrcUW/N3lvO69yD6Wtdyw7KCoEqimBk58+KrkLJj9V3SaikVlPlZAuMUfgY
VnHtZf6gUZqBrxmxq3Up7owZqoLHKGtSUUP2Y07xRV1OHesPoZpae/TvvHRHaH35WEUsdDmXubbe
CmdLL3RS5UeBJEGlX8pBolyFmW8FX3QdUiQBmweMAQmiNtO+6F2feOOmmKgUcq7SNlVKfBfiw86W
KT+jX0umXTkTeQTKYOD24OgHEh31kyfKQaD1FY0rz7TRLJO9QyZdQC1jtXHgr57Nnm18OE3hlTs1
Lr0MOm41G0txb93VWm8oF/WuA6Kf/CQVaXfRqG5SHQH19A8P443IR7akuiEb3fONjjbpeEH9IFK7
MZxuKu2XlnYd1auDpKBpjJ4qXHGZlinL/UIKsIW8EnpZ21f3eLGa06ZPs2AM8dzzJv5UM5OszK0/
MModWNCefCNkeDSJ1kLGQQi5wgHjcfpVoac/+T4CKHyyTHmUqURazG886CafSbY2OaKVyMwap1/m
D5UB/Q27BAkF7K2diTUSG029pwJ/BNxcHZb6qaZATLWRbraFgxVFQK5DMNu2UzhndtlCBBMlBrh/
KiGScMcbX/zihyjexSiuRLamWNapqzdRrTCYkGdWbRCP8uRk//DUeYnvGdzUohFJzQzXz5czeURl
4rZZ2SZThw6SX9t+KmQ0ULarYwM8/zNbbVVxsmcXLktyIH9Zn1zpbF82Gs/8qcrGbUlqY1BHWaok
5rzf2+uEhD1SUSkw1uh2yikh2zgxAKxvpKWalcDq8oyowfPO7f667obMYmLCsevdK9nsLATp/RYP
Ap+uwCU9iPKck24qnOHSM+jHYK7+zV6hjMzQmEtU/HQRHtFUAXZebLje40YZMqhCWfvbgTjqY8Kg
gEJWk6hL9wJCnetsQhVKHXkTeHZGMW6DRaIBRFTqUXMbDbniWg78Gvhak43OrU4wg9kJ8U5h9T9c
uUWLkYiFXlzwpKjA5Qbi75EDp4eyrPRlz+MfjytNfPRVHCD0VAxsKQcq1CQXoViFbWRswpty0ykt
o9IxZA4rhdvpH65XGqIwdIP0ARoX7taWHN0ymRWmLTmzUcwKCx4yyXFK+tLKd90Rc/fVx5Nys0tO
BjrgA9VTA4O/+a98/OAXycaXJtDVUD9nZwrE2Vkd6efSr1CvfFv+2dnMhcWZbs7fZHcBspk9dBSe
tl+K3VeViBXMslKsiD4H1VH+/38IlFCkZjbKLmvxFMBsPma792TND0RT7a9xAY5uvckdoo4sAK/V
JjivCaLWKinyhdRw7iXg0XNPcHlwYztCYGUkvIPXvUHrv9rJa3JfBfLIpfH55gfuh2SRkQm6JD0Z
niJJEqa1cbpZ4TIMl/Mby+JEP5EdHrjK+YHTuNgaqGhdP9AIqBwPgkVYQiiScFUkelABxNDL0SAH
WLrgaR0xI5bwkUrpnXO/v9WlVMfPKP6c7Vna4LThi4NBABMFZ3jie1s7JJwkRORGz0Y5Cn+UeEmC
k6Y8O0iG8yOZ2h0WGyiu7FHmjXjGfF1EFT9+vSyXd4cPAkHchxUbN1LAq91OUCmsL5kC6HMaP6rL
W9vtOrH9kMkv3PNl965v2Lg9QHjTIR6nm+hTe988DjkSvb7ka5JrSZhP2QwAqXS5T3LN2xMOjkqV
f1+oJKdq5ANeVpuXBP5MwGPJrWiACg/BqInRIRVk0ve5600fv54N51AP6M3OO0JKFufU+elT+J1a
Kw9owCQujVjm7cRynniG+ZGhszSLnWHNjqAYWvGQaWPPQIRZ/iC2lL0SeBuH/nLK9ZFnpjCsGDPq
eIsKHtVeQTak15I+LjYYHla31j2s9ao0nCrOgBQhgZh+Op/D9okgrSPcdrpazti/umTbDgBY+H1c
t3LWd9O/3U59dgr0aYuhYbeFkd39KIfvM2ufKilKLjLdwQ1X1bmVcTpQAQU3PjuH8v+RFMQEbOFu
PJoszQw5UvgIgUvSH2tSTN7zII5hprgG+NYIRBjg6utXzRbdWbwr7I/ZTZln3BxAQxhvc4Lphliw
6Sk4BHFVvBQ08Aaaj4LX2NdDsDyyyS+Sy1qQAEqMn72TE8EcrRxQiSRrX/Zfi/Bs87gZEBeaFxqz
cWhycQvwvSmuhy69xs6Zz8DjFiQ7xdXEtXU4mSJ6hCfY/I8OzZTWoRVaNFqBsLYUD3B3M5e2uk/D
+3XEYvP8tR0XFTBaiLjaE77yIVw7A7FqnEQ8ZF2YdY9De4ccY2rTw03Gbo8SS6kBBZC6wCnFvVjT
mqZxWj5pLdDDGb3hhdAJpgNZAJU7fhCCw66YXNoYLP0TfbZr3NHE6s8fo5sZX39Wg87t2O0J+Dv8
P5yADC2GSnbC84bUnnCYPrQnM+xDaJSQGNt2BA6IsPXqu1C0hKf70eIcybNkClRjYxXsyTuJ+I38
HDFip7e+wTLBCCUNx1mtcAQY9cv2lDOjQWwBH/jAaft2Hpt7vpcW6c7NHD+jscdeisApuZunOpKD
MZWmlRJ7I8kVK5zFanXYGQtBwYcRlmSqoZ5uear2g3tNSBfws72wifJAdHibLV7E1PPbZUw/AZmb
Ddkeo6HQamUqwuSFDMnU0MUvXZ3JU0Pw7C2v39T2CnffY6K5jbVqraCK7jh7WWvU+wLNHlW8oJHR
sMchUkX9CQT/HHGYrfjIYdgzAbOvLs1kQmz3enURGy2fT2cIByTd5vj9SQTWAeEQXwHbqKzPl9IR
wC4GXkrzSSHfDytkjJ6o88DuMTpA9Gd4hp+oPaPCwJktRqYCH0TbTXYdZUSfa28cQl35rpmS60AJ
kq3WCHUk7PkfG9fFOQO6JfTK1rwaI/8ORNNR3FrZBuiyBklxV9HBneRijMIxr8/S/KQfsb7UO+S1
9jCS3ylc9JZmH6gzY3doTI4QRZT2yr6es9PwjjRoGgr2bRKzAE8yr/Mgbt8B0lhh2sNBQdiJ6nA9
A4FLDiSZQViAUoWFcioAJym73u9iolqDpddB+vA9yGfOrKeP55V+tcWp0Sj3q6ZhUDqphmkG1YVG
/QGRRfrEhrx4M5CfeN1Q8sAVB3wbpVvBldhgxIAu4nMgEMzGq0SO24NBQhtIv48ZZG9KddtK4UQb
z4kr9xe3bw1tb1wPZpApz5anl9ljPqbtm8/vu9K8mAXNj4P4ndF2wquLSbaa3CvBfN6SbrNp05bl
kapxp8UCD6Zzo5JUokWlcnfmJCMNeXFtcedPVe0/fTxbs4VyuicqVo/ZFVM2BAQAWLfpcgc18LkA
7cWTg+UNuM8IwbhESd0VifyCH1WOSHgMwBoWREWPKCqOJZFPjD2MeVljafEsRxixbvFQageQYlM7
FP5c1076mpoLkBcn5hnqwka0bzHmISvPaJkooRsWDhboRDTY8k9RLHzGa2WgwfoDrWun+bsAa8tX
Fk60N6K7pK+JTfSysf9xHQmk60fFbtGUChe86HeuAe/esBT7C4CP1GfORfF7EGO0Z/5iX4LZPWBK
baq4EjDQn/gwpIHqMBUziRHxFqV9GSK3tfqRhfAZcOMcZUwOJCNmsltVWHd0Z0Qg/1QyZqU8uq6L
NG6ms2Oa13t3z49krORew6UfHcRahJJUsXKUgkSVkLmFTD6D30M3HoNdPIL1ICh9NsbCjuY9zJ+r
rV9ZQSk+07zb7e7QmpI2b9xJyWSaAqT0ziz3wtSh943x/ayKTDOtS6VR5Tuo0p0MU/f0K3EUxI9g
J/+eiEyHl/7Q3Ac9MlDfNZb0XwQlKg2WAlL9rrKZfVUxk7NDmSaXgCtbT+1z+z6ngcBG8c6Gidph
OShKsli1xZKFNz7OPcTBYeV34s6U8lsPKGfGn6cEOJmFYIoZrt3NMFcDRH7oaIf6q6a6az37POLU
G6YI9MnJvevyFLDvzH3I7j9wU+wAZdJ+8UGbU4E2i/Nk+akYMsDOt5b4vse4cXfhTYrU/Qs06JY1
VfVB1vBOueXCf8f4MkoF1Tkj76OF/nPeVyTqv9azrU/ELhq9RcCeQwW3wufVdVdKvxzeyDwlDKHq
8wFLeaRHD06ob9Os0+cWyJUplf8Mdbozzaa9rOwr+8NXNQ5JdXf3Y9nl9+P4q9kfOiLo6r3HQE3t
EwL8zSyGSgILrBm2HefwwG1Czy2x6a/A9T2fWCQWI8OKxX/mkwyxkatC6l+ZwCjM3N2WT5oXfHMy
UF0l0/Y+i2rjKzJBzdpDttqbOETQWBjNm8Jpc0Lv8X+/7HccrsTwCynfPmaMrVw/t4N0kXMIFCDP
xE+tEO19siBBFVeJ8Nm5pX6/Rz3n7+sc5PbI7aTuW+4Kl4aWtQB8wJrZM77GbbkeUkz0BwbDle2O
0VzJBW9pX3UUReC5ywpA/74OM/mAtAj6AqxaGAaFTrPg1PLjUs/5wGWP1hT4L75yCCvgFPsXKn0Y
8lxMKuRlCwPzWQrqwCxXFfVzgkhL0TL9uKQMkah/xjZnjCWnHyMZRin/OpDYB+OrwMqOgyHcL/wc
OMdl2gLyp934/S1QVZHROLwfbD9yEbEty/9FIv1vBehrJaSGE9gmT1XSkEonbdlZPhLAVgC2esEF
Ay7cI00UA67A2Cx2LidAL6Dsv0RyBU26OFdt5ufO3rmmq9H/xd+y1E2Qo1ASTbIuWKFPjDvYxDJi
0BKDQ9krO2+JPexbSxV0jbLpjkD7nSbMsttWXXNu6CxO/NyXVVS1W4VnKVK1K5/p0rqQfXP1JMPu
Ej5tnH4OMlLxOuf+i+FPGbOsL8UCJvH23Mn3omowtSt94wlbgs1u52jShZ2OuoFvMjQIr4sY7Pe/
g+wRfLSUcYjKBoCiyPZgHPdsIzOJyt0w6t4k43vxGchXBdOibEpz5r2kiuVZVX7gpH7Jc7RM0J2J
MQCuxsdtJ1Q3J3YIP0fKO82z8U99QOHkD2o8B5a13CoP+A8S++/2k/5Z7aMPprv90d99bLUDdsUK
G6dm7d5NMzIaCwbWHGGg8LEWo4vXXrH1r4Q+RVYVk49+s1fc48quSiOCZLDZNH4FSx0NdjmLh9VE
eZOhot1sAenAfEaDQMg4wbAOUsFlaNRvCZNlqpk9cyQ+phgRUuBOvJyk7LM0v1jWyLyAtzeFJ5gk
UCQ6MIMSxnhSh4NyukPRj332QXfuH2uTlLsQ7D6bLJ8aTZxXx+H02rmvq5ZBYHFDAdWozeYMvwdM
y6wlHc7AL1eWvNLD3DIWpm9wxs+qfHAGBygFLXs9Xiwv6nX6o9DkR829sYNeynHyd0WVgNE8loMB
a44rEOC4Js0WcaD1F189kDxBob578IS0zItClYVYKaWjuv13Lljj3D5izDetUY9xOO7ByOFIvEj9
6a7jGnGsKwPn1rDVic3rVuOEZjVY155VonI2ZXnpxGC3o8dkGYHWvOnmDSi6WeWM7RB/J1tglQrp
F15ks1TX4UyByP0qkUslmownILS0CfFqaYdmtfbz8evn3TcP429KSq2Fj0g7s9z4dq7LiRpJoeQ0
M9Itt1jM+7PwblPlJyWGs1MPFviQpuyYHKXQ7gy9agQJCD4k9LXxmEDJ/+l6ZCEtwBoNmN6nXkTD
sVDPTT2eISXGkaUG/vxz677sfHFt4s24PHKZ9oF14MnEiVNZNWJxT81iAh/xkeWEifMS0dTSF4Ch
PQxW2BD795bKu9KdHpo7s/1Hue1k+LFx8YTWlhzMkfr0Sxsp1lZh1T8+s1FFquZjuQUaboqDtV5C
Epble1ZmbG1bt14zpQljIqRM4iBnAbG37EsbhkxRgDri27z+3EaKJ4q6I9JQ0WlxKqfH5Lcq7syG
NMgrfk+VqE7FxYeivof+7cKzhC4O2Tfud4KVigM2z5PM46s3dB0W/8sN2Ev3cHKaQigW4xhi0uqX
wKaujD5K2ihdKs++OmdOPKRgy8/KkJFHBKOdz3yspb1Ip/04uks57YalyRUO653ey+kPseUpHSoI
aSMtt6n+d4jPvITpVWnG19ZtHX0ddWS7sB305cDKkR1XonhAxttu6VDI/KlqDNsqUEEZBRgSOgrG
TM36ePGFhQF7R0EQbGhjMpD7fmSYUpabTHM+kRF9tMnUU8nlWYpgdMIjGYsM2vVhi/IDpD7Use6M
B2HZUFuLiom62TxuGeX0jAriPHBOoIfXR/bF7jJGEV6Khtph/SWzH0KNiC1eR5Woe1zT+bH34PR3
GxWj1/bMAtzrTjakPpGVdmjWmvBkkq+quigdsLVbn8jUCmpWV5qhdgpCidmQQeGWGntFQp6qFwXy
YfGX3CvY0K11CPUpcQNW1D6ddXo3ymYnuroyYoudI6TvfdRmBRRror85y6lsHyBNqsV6hQcqmwa4
U9TIgBw=
`protect end_protected
