`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BeDk6slWwyJ7dkKWyaZdmI5S1xnQWnB2oiiYkvyYe3ILPohOGwb55RsmeeSbX1QjJu01hxqQuKng
/gQKr+nekw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ASzYKVAZmSO0SmC0FWgRspy8UM6oxvcf3jSUzSQ5aTbQcdQEmkCnyOPWPw5rhfBxgGmpUIes9+yb
Y1HX9gskfNW1iUc9hvj0/7i23Dl3Awuv9PwzU2qkFTur1xa+VTaDhjRdBkmelm1XEmzy0fVWfN3E
JrqrAgqGTQHZ2JkK6Bo=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oJBoHreUf2ZGu1uujJJM+r+7FZbqExapJJyyvy1o9iddxQis4QmRw6/bE0DAY0iOm9OEPedgUYiN
HJiQO008872laIEmtmT/BZsMbhdVL80RK/NlqxNSooHOOtA7Q2ooOW5Qroi6pqh15Of2uGz4EX8r
QzKai9gyZ1nNfMdTAvc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gXcd8sTNtxVLLLKC4rAjsRNsfX1NVlxv5NlbcoCN3RLErB2fm8TB5dri0TbIQGAb+HGHGVOVAHgx
uVooaR3J4n0jcKalCdHupCpw5tdmXAARWsN3+yNMWjktBvDZlREeBk2BplNU4DXuIjpyRlcW28oq
fXURF5uCQelaIUMgDwAyoK4ndypdafocPYsPsbB7ZcLdDX4H5Le9tBCnXO/3QcalHHXgUWKcLkyn
o62h+Ts9twP03kQwoK/zsw/Mj8ubV//CFoyYXoAsGg33zvV6pCpWjHcIR6qmaj3YFStAb9Gwjq47
yV9Y3uGyv5WU5KKhj3xqBA2tQXCqQY863nIZnQ==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZCOLBlM+DOBMBQ8zvcBqrtqtygwYjI0iydlVEAyokc0UPDasfRQj4taurJsghnxG4bETs5xI8oYV
0HnNJr9QlLNdd6mcJgJqN/c90+zI7I0/hnO/qlv0Pup/OiWbYiiAzYaGPmKRDqi7WYyqSO7I4TS2
AG2Q/zR6LKL+UR1LQcmMcJ4RgLFqPmMasX9iUCz5I9lsv9KntADfsOLwcJl5QoT1i4VZKbohe5Qm
MESQHJetAMfbworTVW5vJr8gNUaDSSpP+4845B0JGNCebeUUC8/1KVkOL2aPgIiLRFtWjAGp0OdP
Hgc1IPHx2d0B9ihxkm+YRP31ignQS302EQYvBw==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NrFXeDUSk0IEdKSAJNgkeyX3IOnuNIcPQAo5W4y9LavsF2f6Nt+rduqEQbagw39p3ash8XtbR/w2
nbOm3koCj/8C0OoRET7PqvN4QJy3y4VTXAZe0/S0IrLxQsNhhv6J/qZfD8QvZ356rQBjqyRt3tes
FKIyW/uL9wD45Iy27+yn385eZ31TEAWa3qUWjlZ4QirRNAT1OkORBDIQDHOOlrRwhcFvBqpmP+bt
dB3NdDgt5niwoonBSPDFf2StNdLHNsQCxz9zmE4Hap77op41g4Avc9CdLgPyKBKRlvYKlsU5dB+X
7VzJf8Jl3UhqXRVBX0i7dzEKJTZE1Bhvb5jelg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16928)
`protect data_block
YzO9pHxtvhOPxb1qQ4BRxhcexAT6MOvoLoMQ6pEsO3MmgUGxKQPyDpDUSAig0CKHe6C7zFS10HIf
z1LTktR+WQLgK5puIGhWBRe49G6eXAVk5x4XcJlcq5nbELFKxFMqyE0iC29t69wCWGtbAp+OxoXP
4On/waZTrarFiqYcS4dcxwamx2QIOREyoc2TvFT9vJlLd35QnK8gfmOSp8V+lczxWH432Nxu5ozd
dM0Jk7/ynbGqY0lgnaaBSlg2M6wqLqp/u57hgbf9S3UXnExl4b+4FDY9ezdz6zJx3T0yjl/7Ma3l
djyLgS5thvuakSPlsHiij8+fV8EpIU3516L51gqy0wUcfr3KM3qyOLB25J9Q3JrTM+4gTH5ebRV4
1nCqR2QBqW7I6JQBszWQ3ANyndExURqPKbWXvUyh4o/8ZVZ519e/XAiX60jWoEydiUFuUUmY6KNV
kPy+XHMxMPeYRyRMggwZfWvd/+6FMTWi4JpGz7jNTYEtnNUPP1oK/PudDJVkv4OlAJkz+oUJ0Lt/
Dv+Dje5k/4BxCmlPKf87zwgfN9oFTqKb8zGRFifF56QAj5xrAe5ojhchHTEu3lnWR36tgV+2hJFP
EjOgRtn3ISPK+1tQFXmP+N1qpDmyFtawycmDalYK3XK3D/ZvrNZLMv0MpTOoYu9fIE0P/vCVj1qn
eKHhuAJ29pZHbqNlZSg8CDxGZ8jaSbF7xHZcHPGBF3FghN4CaFuvnxH2V+Dnh4Xrz1bzD+ZqNZ7F
zYk0wERZDDFWmG+0jWRLUS8Fk5C41wqQddsxT02eiVtStv170cBIt/E3hivC+712vPXLpey7jjCK
3YNfKk9tXvmwzUimtuHE4b5MLf07BY3yc/I8CGlt/EOLircGKU+KeSmxK95aBi+2ucY5A6ewXakS
2nPb0e5RtlnBXyH191NkIfmTEKD5aau57JKyCkwEJqKw4CkQ9aWh5JIVRnBMSQT3LpsL8NLHUBMn
7KBREns5og4ZBVCbe3Pg6rnCemET2PKKBeWgbM/0qX6oFR95RpNKBB9KU4Te7KodHRJU0AynrVPH
V/gFjmCtsnDCBs3FK4pierSMxYJpD4Tm/j/MMNfR6Vo9tX3dwc3ctkmgK3W24CDll/ZhbiM7qhch
bKbZqAt57ZAyzkaxfhvviBmwkJYFD5+ygIAyaA+/5g+s74A3rEtrzLt4hmUc/PrBpgvCZCynJVfI
arbmNz5nA889Un4Rj7t8rJGl/1yLZK8CApLnIhhT3Gf+FXaewMXrF0wf61vzUfg1C3hR6o+My+pX
0Sf33c6Gl+2ztdqpDsKNKeyJfOM/qGQ3L7kzLhmGtLVOTB+Wq8Aa1sT5VLaO3psOcOvLkiRBgfM4
wngrb4MMThiNii67oG6LgeaBHisFbmEK3CaZZ5PwPQuoFPpxWp7RdgPT/mij0fkxwG7NPLrpKTos
99yheDl/EDGNX3X031/kmUWAhxgfR7EZpdAdCdMapg/qnAWtusXHNT3waFvKvUlvlQvbn0yX8p8p
JAzmfnbvbdCoYsSqlMR4c4F7pkYuKJotCCccCWA7HvLdGcTs4xudLT5wHBauV1FNAXtnthBJQiZu
iyIea9cM/qqvRWRyDM84B6k0nRg8LqpIAv1uzIh4Be4BqoY0hKw50rEbRb+964oQdCywJlY/ubPY
2KERfl/yQeofLP1uDXd8lniXOGIE2eIS4ymLNUXvAjy9P07QsfzOVI075T+3kpUN7AncEEoWCbcZ
TZsrAc1dccjdlyy/CZtyMGJWX9is/EU8jNpDXgcPErrDvPW2HUYDbzgd4An8zcfGkHmMDAofho6e
OOp1YLL+zbm0HysUnjsnAatDyvmsM423hCLWXB3PWlxOXiq9c081jlxYz5Y2YY4q2yZrEl02NxL/
MZ1w2WyT6pH3QlJ/MSRq3A5fZIw7d/4IrJLnnY03d0DH3MdlgkMtOkov8PTiW70NMSEI2CREG8FU
eJyZtdskf/K7r4GQMr1eqRx1Y4wIznvvFdB+xIRLp9wiVBnazd+TCptax743Sxwv+Xni12bfrYdJ
/gkzdw1JHf1kyG5XpF9lxHMJRzCu/07kE+6qvJDPwl75TLfwVI0yb9bIpIGzDeZximO9bkbY8uOy
hirOLeaOWmMXrnLHINkGbwIOOE1ZsLTenT8+T+bNURvadxK8BLbwzAwkfwWvEINInKjvWhK+91E4
PMpi31TQ/hYqCAeD6zk+LZx1Rf185oykNyG8Al4q9bD0HYRprgvFt0dXCsEA57r7QEpvipnTnbv/
k7KTg0Qm9exa1nF3oAYE/P46+sV/pegy8UjzTq9gPAPHpLVN+aThSUdg78KXc2uou9GyQymUinpz
Xhao4MKLgBHpJVcTWNM4Y6e0Bbs/qiFjz7h5wM+7mTKfHQZXDaEVTaxw/mpt8yrMN7mziIdvE6a3
jXSjyWi8YA4D3+hQKgrU1PAaTyBVGCv7d9T2RKbMDgymMCeFMICOom2zKxeCm3h29m74KP13Ag3C
dDUrGsHltOSnT/k3NPj24mqdHcoo3WUco2kSnAsuCjCOgpP9v35BOdchO/2CoRfX2T57/rVrgh5J
usDBCxOV5XS/H7mmU1xHEZQAo8VlEZ8R4SAyupaY2EAl/j/wePsYu7VWU8TyxgEGJy+O52yu38Qu
fC+uLrZ/7Dt2nx2HVaqGCguOJE0HYlvW5GKgt9couqwP8omFZGOUQwjW8WQ0MlT38vTf/Qc9exNu
V1ozGlMoSRawQ4o1UlZqypiCv/T5Ah0Im+IMfE4Lp9s9l4UOfv57T8P0h6lyJ4Zhm7ZnFwae1hXc
OUbwtlF+3BznRGZogQvdNxP7D15z2msDQnBR+Ki73RwJvwXrJ6fO+d9tuZrYBSH61s+DUTyyjlWi
4ofoug6VKFPHLRu48NtCdMwtKbDSwmljH4xHB7QcsTeNq1baW8WORwt4fAelRVzHhoxq7KC9zCAe
wAfHETgL9Bh/J1fsp3uih3MEfOF/s18xpSxnqDSs8Z0PRIyY22CEsSmFPbslViQ7XoR1hINO+Q47
Z2ZsQya2/dZ2jgtNLkSfhU6TFc2cdHKakgvWG6banol6Ai+AQQGCV5HIrcftByYt1EgWCAxhVFfV
jq4660P3caCs6if6w8r0gmB71+010pLbAFNfv5A2GSTJof/AdJJEzQB5jgBDf2KlgP7ok809dwfL
EEEoBpYGtwJp2b8r+xU0eQArkBZXFmi9pbZv9/2MO2w65tgiocVZX97734JOTYJRRdfR0JvkxTOU
iNStDMWK55nSYg9DDYI1k29t83ws9qgdYqgi+KrOA1TuLdOkHzzMoVSfO7D4iaCj48xG8afDmT6i
5wGOR5TxQ1u4+Jv5+KBORxgGZXXpmY2G+CG8QbJAlNz6b3GChXDQ6vwfFA0Hiq3+rjBx5Sr+1SQV
Ofqgxc6CLGnr/a5B7rqkF7tipPGY7bLHWGhAjpfMUHHZQeA2ud2dp19mCtPFEJrzfgDvrQAaR/5L
fnKBylZJb2h5o2X7IroEFT+BMKqTr+tKm2UED2d9SR6aoHxRqyvqhhdJ995UbUMEjlrOE3z5fNw/
REOGM2DrxEqXfzM1tKvb6exgp+35RZY/Bz7AcoZJ7bQyWrEZXDMV7M49VzUfVVosi+dj9sW/4IAY
vxRP3tn8x3dghdzhbABE21YiGrBZdj3AsdG32vccx2FPCEroFNSHnwcTYLTDxjso4n2abqjcHjZg
cphLGrkehkxYQ8DESFtBYWf6n2D3Ri6/J6jEYoCVRyA/WjNdYvTacUArt6cuuVSEct8RMHmALKkf
srr62C/oD9ejQL92M5IcfVQaizZqGx9D+am8uXSqJ+lsWmXne++doIMh2OIPNySHBHgYtDlzQX0U
rcUxd7l5sF7gck6lfEBbSZ/zBzcNyRiugVJ8t5I8wkXCEyaAM8MiOjlnErgFW9BnRvuLGP8FUjXX
p75ze7DLS32fSGbd+SWzH6lsgk80XbrQFvEoJXZ9/JTI8KSijDq24udcksiYZ5j+Zutn6aUQrs+h
5mC/qd+mSuSfXnA1iOPuUYFTx9R/N/Uu0NSOwW6X0CG8qcFj7YWfgg5fRW8z6VnbJoS/PsP1PY+d
HyBWDn5Ud3Wlv71lBe/Dpi1e8LLrDUqCTLZip9gv9DVqMpxRROD04Ut3a7ixXe4Cqbpp68X6e2nW
VPDbjsD7kGKB2mJ3Om0hL2119XC0OMnzvRc6zjZ6LmvWKfIY8RE1m+gseBLoKDOFQAUe9Z/zrsgo
KISXspHs5AmtQzMoBpRPOvJh3sE8emvZeFKYyyDDjZlDbErfKZokCAePs05P94BDfNq+jFdoxEGM
XusTi0+vaXVhLGPTw5mQ8ITjEEGENcAznPOZnPPqcLiZ4+Uu3amMkLoCE3dKLQfn0eU1fpExSxwu
aEsHwfe0rgKfTMi68rbRapUEMBNDAivZm1jNzvaJ2ROQDtKyFshosLzjIYIWJ06B9VBqETRdjsMK
PzxuDNYWN+l/kpL27EONLWpaaRuN7bKo9W8rvJvhWacelzw1zKt2dobDeaNriWviyMZsyo4NOraW
usTds3mYgZFOosjXC5b8NPH4TnrEUuMEuW6V4m0p2Ky8QhxJWqsEjJq3u+IIam9CQKnwAlV0YWH/
//wnsHRBjiAu17UmLPfRfCI2j555NRvpc59uNi2aL6Rv8FbNv+pZE70jFYd8lhqmZSa71BCJY8Ah
vel6hPssqEfZZGPRra0PIt6Lu1uJdELNJE6kV1MXS0ivFd5q9lhgyTUmQS2BoxTrD+lle04u+jwt
7PbK4PoTkotIa/oCFyLHFmzQk9i6G+rq7WOCd2oollY3CR0SpF3JW/qwMeW5focQgSDWhl0q9Pnc
xcNe1brv+kd7Mn/QQSRoYwPVtFnBItexerRomRVkORVLaFacw/A7oeMpnM6FaMbb8y82nIS6fnqK
Z9FROsYh2qWP5x8OA5DQ/tWpBfhIADrmgf/XrRy2+uFwU+e79xglybaOY5bbra6ptptg2Po52b8t
B9JKCZftvvc5SarwcGbO/xX33i1Fi3svHP7Uk6mtOkelygGX/fr01E4kCSxxyiI6U/d2+TEBMxXu
gwJBBfyFIEy8qSx93Wk8SoB/kKpL+ePj1lF+0BaaNdmZYyZBJnDyz9GQ++5gZZzTOAN1r1hdVuFC
sPP1CpFgbraNVEVnc61ojwNhkm1w2NffbvOe7gTiUk/DDgjfXU1+rvwilundhJ1hxdpCe/sAnGxv
HTmoEOPRQCpny+BkRdEGUu1Gp6Hg/kdRhME4G7yNr3YdfJrdGQ2TuWBLpoOfzXLx3OMcHeVyAKcR
mHo9nR3tKSRsClSB5Nos+DKQRiOf9TJHKP+c/MpTQtxUf34rseEJcXWFenDiGyRZCj+X29GofxbV
RduaRG44xLUZuuVOONVWZSweMrR8jOxl+7yEAM0XMRXAw+u0DH6XS3scmLwIJm6b2A7BmuLAjG6s
x1tOKDk4tFRgy47H8f4v+9DoXsCgFUhNux8zd73bnLWtGL3zIiPweMaqEe3CHjPWNZ5bEpMT+Iyw
ijWBi7nWJEPwj6OVQ69Byu2ZI/MyBU8PfXq/amjk2SgpOh7UVsWPqNe08NtImltRcXlfaLPtNDSB
DvmcR7Pz8lj7o16rolsA3w74VN0G+Zi60AVIIt3WQKL/EfRemNm/FG9GLihPouxlmVOUzxzabEuT
Kmd1ZxIL6hLfBpFlxa30zKPBidyke+Zgy/8rxpvOe0IxpUuKWVFA9aWLxg5oHy8N/KsUQ1NR80aZ
fyiUJDanyoVu5QR0ODwUEwNGZM+YKnKvrwh2BjwFlMdlrR+cbVBFlQojaM4UGet1YGraabmO4P6u
5JJXU9Zfk8DGe7L/u0fwLKoJ/bIgW08rU2ziIOk8uh0VJhEUDMjAZD97pKT/PUGVhFB9m4v6nTRw
Tj7cZhO03wg+/IzsSgXkCNRqvGXNLjdVUWurQ8Ywxdqze0C2nELe0MCMAuMzpdbxXjdzjYXXPzsN
Cvxo0i7Et+up//NQdW2wL5fd/lNlC+QkwI7BUN8yx2G4yLCax0JQvWfPIMJLmriOHQKmlTovkkHV
BsFepNfHHCG6Zyp72MF8h+Ssp977n9zuxmA3GKNagnQajdBgdrI3g/8cGsvGpgioq1qI515iUs3w
8fPP9s46VoE2RvSbxE7gg/mJA1b6ZbKd7I7UGrHIwHcnDtNx9j6JEkuoi+ZCa4yt9G4iEpTOH59v
iKSGNmSl1ddd1KlU81GpLwIVU9S6UyBbV6NkhL1JSiDE9OdBEssABf7iP7EjABp9tdiIASyREhEH
vZ5M3jPgbNh1Kr7fnfveG5ZxkUKDrEhLU4LHAJAGSObkVM4ApRTGw+MX8gpTEzSPY1KYRCtk/Lij
EZV6z5aMkG5JgaS175wXn1mvsH75zNYizONf7Elu+0KVHcK46gOdMe7ZukmcaYyn5UzmiNKxSgWp
ADETRzX7QFOPOJ1pbu/IgOWFp+O/KpPOW+vT7O3JLA1DBLC66DBCduEUrTfr+IzckcOwwLbzHlV2
9xZOr1CUHrtE/Rj5vMbZo/b7b0jdzCOiy0DPamWiqOeQc0FsI43RuvyjC5mf3KkWSXiM3JyWbd/c
ICkLFwomr67iyl/K1mLoYLap7FWY2MdVmBWwxuLev968l9NpNFvKI9l99cXkuk9pO1tupk+lx1qO
DV6JU+ve5KaJfdIHrLq3+sTNXZAn9luMmx2SjffjnDWMugRnKgKtO3xeiRQkBnJEJ86P6VVg1oCh
Lhn/I8qRqGEd+ZgqSmONahAm3rNRC185Lge5Irp/70lToFp/s55sAmxMmYMVXJWpY70wzh7znXh6
sYRtEJISUiMCMjgGxWQ+ZU8tYSYuV49j/R3Wx1vAMJDKQOUlRvpLQFFLHGfjVBf+vNl4KHhVfcRm
KQ2BHABAYo18zggbjO5vYebkhdie5ffIWg0xszwH9lBjdeY+caNtC2buEYvjPTEOyTzMhIxmgqz7
G3wHv3BYF2sZRE/tGVl6VqPghJMfMnhjn0i+5+UZPfIxWjnA/+kiCTa0w7FNPD0VEu+sxFRpcue9
Bd4T9u4UZ+H2AtuhsydVoVBW/na1j+jg1BXYDy4fXQRAzeFbfnvHCih1NMw0Oylr7bD+v9CqXNIW
nRs/wxcFO5ze6IwrG6NvPNh4x0TnJiPCGLMwFbw2Z3jV1F4El7s/AmdM6G3XkVFzmaSFkT8586U5
6nn+YPkjSHe69qYUn5f0w6Jf74TaWZoKroJoDtZ8ZDQo+lhc+/jk1HvGLQgOGrxuG8Q3ZNroxBdV
uP1/VgCgDq0AMGMXxoorOGO/FcxlJGv94ZTRX0T6OzNY5tZ/53O24z3tXugqA3CmOJr3BGbv9lJt
dk4WkuABSIl7puHmLiFi7hZxV7/lQdMwCx1XT9ZawuQEtSA0hWrQpWazLZ9C9RdWrHOIiJ1buwo1
UKACGc+gD0u0ZHKYSsPaWVGPEbRunwgYFvswO8DMrZ8kAaW9OMCIfkkcvDoz+g80jJMfCS2xK5NB
lF2FSodbEMT4qZGjAxOHAvOT2DhfZPkd+NkIL7DiojocXSJDGxosXVoLM37s54o3YWnC4CDmrWbj
1+MwFg7JKxhfWF9tzILkxHccN3Ga9h/wQqTReyouccn3dj0EkbDJLlGZGf3mL4q9QX5wYJIWHWPc
CDkZNUDrIzS1OyZN7hYH61nCRsYR7y+xQ9hMqhpFUawR7GqtYkSHv3JSAKtfxA4WmDeEvI/TPoAp
Rg/FCaITXRKqit19VF62IUhB6HPd2dNi5qYozv3RVHDip7VGqu8LSjY2p0TpRcpom4kiaIanTkfs
9VVxMtHNFXUBdQOdqffOBs0zd/65MRvP/ZOXhqjDZYPWbM4trqd4xDeXi+JmgMtXP8YvNGlk9/yX
LOxxdl+XdEvsp9bRHz4LXiJ3fcGSpw78dNKOnfe3wJ2LZzfVHveZqC9Cd4ZxksxapaQ/LU05iX6f
ckoEpspr0ucg7Nhwd0G/qU1ocqfMhwN2yiKbvCf7+2Izw3pqX6T3N+p9aIeTfATSZ9/m6qHlDqNJ
bh7eyHe5W7iFvkxPnkygAJ87KDRkmyj/iELBNm4Q0JqXepBvIdF/JWqeBje3YqliTFlM7jM+bGsK
f8kIuZdbfj1bQ0p86DraETvd5MetoV/i9BehZBVma0CKwUVVApJAdbm2qjC2xdMBiok2oYczN1uu
MNGIuh/EIPFWI5Y/7Nqn7AEz1nzT/XRYaMs0fnTMIip43CMxgCngspA7H1wQncTK6YamlftFxBYR
IQlrxulfLQE2Cwp5jJbxmhc39cgqJiu8hm5EgVGxBIgqZt8vDuZqDZVjbYji2x5bS3SMC1g5viL/
EH+ep6bdOv+Nwd1eMPAnhS7a07GkeRqD0GWu0K0HPJZzFvZwdoJgG8X1mkhRGlp5zK5APseQLHtg
40CmesVPwoksuUzDB+CAF3PwDBMraCLgdSLQQHY4BWS+g+eFoU2JNJQci3zeGrf00cHzUEddWbKo
7JkOOUtszEGPPO7qFOYrjToGeK71nDSjG/xeX76wCgMeN68y7e7Bo2MtheBe+Yp3th4WiZzCNUQR
ledyWEC0CXIWypNhSMq0jiPujIJeT0IvdWHm5sAPaFB/gw3DlJ1GWGVcYvHJheQHaUP4MWn5QTlO
1ocVQS0tA/tUCfR9MwgrMUXT023bh1Vx+uE6b1wX1c4d/m3WGYzcuD02sesPnRvZVyTSuZa0Piiz
5gimaV+g0sxQ6dRCzQ/Lq2bDYfbCKmiAv+CDOCCXpP1xPFYv3zNBODOA/vz927d816VLPQPrMyHp
ZaLyfjDstK/aAAx+xbFMLOgFiB78ZR2VeRsfX1g6FaTHMBMrr89APYXlCsbgjAEW7MEIMeXgBbQU
dI5D2/xul8k26lEkjuzQUc6tPY9Z6DTVVnnYtN2KK2fiadyWNf75iEowE/f+jRvJWNhuud+n2tJb
rYm+6k3aEBagDPS9jBUk0e6hzeObaWL+Xuu1mjn9QtXoUigaWJCXzXoZbkEKqmRpqCNoazRZSYT5
pCffAjJiYqDuk0mgXFoqzGZKUTEdsBAsScHlC0S5JNRtnUvt7U5dMpFdn7mGt6D7NXME5Tl6rcB5
tZwDJHhcqHo4KlTk3kbLr/W7lh3Huge5JtcW0l84K2ArbFEwnTYBt9r+bEJ+fF/Lz5CQU1Z6YaYn
w2RkoTTarpWmlHSxXUmb1qE2/fEM+jU8QTr4QtHFW/O9EoxqBJEBPtOpRid+gPXkxLyVUvDH0i4+
JNfR6qipM66XC4JOAlHgXYBlqfOaixKDxFMeX+TUS51Nhb/Y6K6epxEyittRrxipPwYOL89aAdJ7
u9MQpI0Dsl6YsC69O0hM8yHA9fsNz/s0w0KjNT8pX/cqzeUZIojtqO9961X5r14pF7rc7G4KcB6x
i7XcptPi8rfZg6Cy1HwsxRg1IYrVkTHh9XkjuaB6aKmwxFjt8AfyLkrSzdbNNxnRWvfdAX0e8Tsc
i47F0h2uv+cagehGF7n7WmxdTo7enJx5u852uWx8w6ez2Or4qHDvSXwT8WvUs6fOkDGzSHnEkXXh
LtkdWf3i8xrbIqcYSnO+aoSYVbVIqO9072O8e+eCSCybC+80UbZ6X3XcHuhGuwALhR503Em10rUr
sXcFYjk4d+WxTH3Ysm4OwQt8xq3CW3r+8mKGUDqsb/eEzngmEUKHdN+bG23qeLwKBKxpG7Nst4p6
ZvJp9MqQqfW/CVoJFmORM9oaJXcfHBCPXD96upJtf3U/1Sqe1YStYYG6F5zqLMwyb3lZHVCtF0QX
HMKKoAGTRhTxDS1Fgqv3ayNdRHhWLWVA/8illEFqNKCiESZ+m+IGJpxlgCCHVtBdmIML/G4n4Zzl
bi6yKbzONJalR3/z8kCitZjRgM7KT/XhKQCzDGEZeQKkTQH1h4EzS+3TO6Kg/uWlgGzxAp5yzJ+8
lVE++e159Iw8VMbhexQjNNGr0YrLqiyHneC5bpUE9+/lGRLAJLSazgbrboTQUlq2iDu8/KotHkFA
fdWNzS08Fogk6NfdUp8YPF4KRq/OO1j8sE9oEQH/G/AnZvZj6LLQQaVTpytolTx2XuXqBDLYJJHk
T61wX6KTfzTgthKehzkmcq4aA6eueRAqCQun4wJiOR4k+d6Ur8nhHRba+KOxZzpXhR2fDBycTlee
Uy6SlGAMxYfEEe3KFPY2hUs/NtGPIj5htit9ziv6st/MslYh4okxv2yEMOFu0mGvQysLlVWtJhR9
krW7nnZqR8naqi8hudtbHrO16tbIPPcQmToY7Nc+qOWZJSuAP/sf5YttaE/lCWALv/4aSmZLtHjQ
hvHvbtCtiT9USt1MwvQ8gZlP6JklUWKBhuQ2EjuY27dcaNxk7Pe9XlLTJqvtFDnxWChTFixKg8R7
VlP6MXMKoz98RSutVye3J3vShb5+0sP0qtrndBEyWlvdeGoihNhDhXS0MTAZe+9XZ/e51zux0flg
K5BHzij9Qs9osug2VUHXeP2ASbbeQ1LBaW9FwAq4lm9VxDW2xSaBNLLqIQKmly2bR7hRBHOycTPP
WvQn35C2kvcjTYgdTyVeZrt1hUdxpljy3MH97OzF1Tx5qoD3xGMkKLD+S9wKnjbVnO18f9LBt/0b
OrLOAhSUcCSZkJXkR08VHROYQLDwOx/W+RQa08r/89XXJlcw0bJsK2pRYBpuO9S0tPbbHql4oU2z
txaionhnbv9nxAQXLpP4/FfpxzXAqQcwY3IVzIBz6/xP/qcaefqfYx9YQqvvou2R0EMwJ1lUQD9a
UtgGEm6y7Yjmycx3xamT9sTLPk1Uj/gotzVU1CGH2b9Wux//EPPkSzmd9LfXb8RhideX6wKpZKY7
n7Mzf9yDqPs44v2vBvAMX4PjhNZDuIG4OMYTkIY0k2RWp6L3kpLPr3DKNE+VmREmX5CrBcX+M40B
yWCOX5rUqruiTLgrn7v0a66YyHOKkLxpJ8tvH7cNX1S1zHzo3adbz6nUEYTeyTT+swtSCWjOePyn
UdQITCvxed3ie/yOmLT4g2am2H+QeyNvVr7FXl2JtzF7OXSQApY9UJSGDzFEbk/xHBcSNa41K6pb
VXiI+mwXM0ERg6UuI8SI/clxcKERFEoBRGuuY7mqKF3kNaaZPZWbsMLhyh0MENE28HKrsRnrUKUm
HLnbsoQQ6r9xahKCzccESA7QCztIgRO8T0krA2mKcWEwA29g9WQoapKUJduuukYIhZ/DJumu84iV
EFO4Xcsbvi38phcxAnzKH7XdWtvZC2O2FyHvo/Ei0yA086rqoUeLKGOqUKDrXhygNHtLAdmbA0I4
dj03RayANvMXIjCJh4ksL3JgGbgqVuvnUsFp2o3W6rqtL6CAc7mpG1Kb9BgBJ8mX31fhF+MZzClt
a1thH+kRklECVH7jTKVxzZufuwxV7kZRO0vj5M+HHRcaB29a1z4wv7A/bjnyee5k1+K57K1j6fmK
aan7F1O90N3sy80iLX0zG5uGljYuY+2Zyq0X86BURJ36vl/LVMBf++fuXGYkUG1paMXAu5/SCoDi
yESqbW8+iEYG7+6isFJGJ0IHIUVygsgpmjGXJsa+HCPvSP4XlQ3mPa8vq6wHWeVRwYhiexQVtzH+
mWRZpNFmzE8ezHkDVLV7Ac1/HmxEtnc/xvt0KHqOUw1fR6W8sKeaGp2pkZxF/fqb3lYvB/76XrRk
8ApHPHCRX24FKAlio0iZGabjed5Un9IfYEI1s3qH7W1BI8yJ6zLdBYzZldf1y9xh9Y2Mm3JkuMzI
JaoRyzjA5HWIZUfiiqfITVQTd1rsSuusVuUaJ1IGouPKK3+O5BO/jMqOnKNBks0yj2FGL/wvL3wP
zx3LDayd6iOTSKJjR6UjuUEbv4gWVGvqt0HmjRr7yoo4Ena/bEhGaPsEntSbkEUceRi5W100rVwz
B3T9Hny2BBhjuE5PeNMno6/2ZMiAoG03RIe5etXv8KrFw0RnW4vsul1ALgcV85oO38TU7u4vs0ts
W0J6WVMlE0+Kfit9zIMxaRWGH+0OyoHzAPCE51dzhmtqH9tHPG4hlMQbGAmsAySa1Y3ddXoQokMT
REVj01mu8nnS5gXFP2V/V5Lchbm7Ca9MK+U59hixW0deW6RrOKBiI1GJd1je7xquqs+Kvyp4zvmp
i6gRqiVCKGLvwihTlMoiI5EPaV7uqYtPbjhaDyxGAMVkHvURKBdrsmUflyyNqt+b775KhbVs+9Nm
BjkJeaQiyTE3o1QSCSbSewKdMyYnX9j4+V++Y7Q574sK5M5EiY0PhZh5ObD2FCpVkqg9F3m6H5jy
N1Zfi3PqZ4ASH6AxQOF9OFOxAjR9P2J/WBhUCGWHPRz7JuDsBCOC9Cdwt6RYhQMyVMQw1Bx69cGp
wTpEz4BpDMXfuDUoA3DuCYAU44uIQ1eTSm3cds7LQkUuz/h2NZZsvRCv9HlOuC0oxHngPuIEsMVm
ou8ZsP81CFH9IDiQNojOnwKThgFo8wMXY1erflq44OayEoPnc6IgsTGxbr9R4OcZ0zRzCmYUv5Fx
rXPAQoozbXLje0KfuqJTFXzurc1w1iEVmRcv+Lje5UCSY7Nio/rzcy5TEnUw519styZhRRMLNnsA
XbBdMAOPUGNNeQzKV2qC/XFumAJwTpN3xz7emhg/cG3FJr0ja41GnJUKaXhTYsVee7B8xehSQlI9
D54IrhN7iMgudyh7nWaEiP07v/XKabjBu9bjzVwO1NCsqaBZAgtEmsAIQ7XOIWBWQ8wM9aONiPhi
+/QlEveXiaXmnbFmuURegSXTEiZG2prtGpQpxpLdEgDHM7i/v4H6TE+dQSHfLKYP8avktUJyanqT
bicwHJfgt1hG7K0tG4nNWgkUc8W7vAECuarDv1BJiP1+0nriDS9ashv6eZUe5BC/DcoNZHYO0Dp4
UoQZzkvvRxirbBZgXAsX3LtLu08md4YyZ6wkUjpjsfM5BfDSo6Mr+7Qg74aoSXY1FYdCc54yZzI6
XvGbVCmYazQ1K9QHANssQeSHJ3/AfsP8c1tqoF+I8b3v16R0RUD8tlDwo8W5h97Yb30fwoXHLkpC
E4U9ZtXIug3mcctdK7aCJxTlGgntztInfF7d1/Y2fJm0t7hIyRqpGHEE2/ZWJoIIl+WK5v5hLu/k
8sb0GwJvt+ovy4htoI/E8b6lYjYsxCNGeZ+MSJ1nT9O2fcEtOULKkYLKeK1349aTobrWTENYkxQz
RaLuFqAc92I4LVYGXz1MxcMf/xhXSoDvwkBBd4LIzILUtx7IO8q9zUBYyBlT+lj4tIGredvfj9QF
Wyam/IhTJIo09ZrwFErCFXR1Hh4Z6Ehr7O1ghNHJ/fv69R0YOyqobGZEUxh5HuWq23xC6eLCaqe+
+TkHKyP0KM+E6wWQoOiAyVSVL3mRcap+Y9HvX302x7+ElYKwIJvXqdd3BGNnPjFRFFWPNop4Fr9Q
E3HsAFHOxSj87Bb4QBIIwQHXVXBx+6Dh+yk4bPvQmYs9SBHT16YxCHgAEK5XiAp/2rYZWuNBdDy0
kNuYj7u0wFVYHr1w6Eh2nZDkmPmumUp0Zp2bYGI9ndioBi1s3L9gW5mcancUvAyisp8OFGIFopaE
Q/9R9PI0ojPvzzsojtnZ424IWN/h4HTRUTpHxdzjJVphgjCp48T3CEPHkGwL8rq3tQoLGiQBJBOl
fvWVorOX6k+jJtrKzNlLYS/s+0x9QlAKeQigqGE3CQxautr7cQ/FWP9d05dUypdX665aE/1B6NLP
xPn0dgvj3BObN5j6ZJQ00u4Tuzf6PnCHcNVJ08cPGtGpDcCZd6RjGABUiMUwW6WDzDy4fF7buUnC
4LNy0tClIw3z0AZ71I3DKOMjWbBeYUARG5s37SDXOV6qB++sXbPUaYTNJo6LghAhlIYnNLNqyARI
ent2KWy+/iJ2N9ILcYsR/p93RObs7wwyA47AuG2C0Unqg45aBelrzAm9MP5VBIwLru1jeZqTJymG
oIs7OrIqWN/oeDqfBnDNPC0gbXakIJG7SOtfRpQgH+QUquObGxxi0sxeJwOgjEgNkXjnIHFnXIpU
0ytHtKYP/gKVMvM/CpYER6Fwi+ERZxqpErGtE+K5bfp+WBfz/+GdgDosP+I7hsdWsxG58Fgp3KlI
onpPyohdIfUOPo76YAs8M2ap0mgWfzNAg5hfbQhqg2bj5TJcsHkZZ/LG6VTrlpRonL+rLEKimUHo
1rN2VY3ZPC4qyycDhthaEQ4rbOX83EzPhtw3pN7HwQgMo0CvVfAMinvNZghTNbWoh8Su3eBCMGqF
dNI4nS1Xz1Xcl744vv1kHpZYQd27ZE4Oh0SuriwqQQqSSrfgwbYDv6brywgg/IAjwpLdbqnVZjVp
S5IMCyRvMLGdydrp+v7NWSQ6vGob5a9wRcGnZeJdsMXuNt/9uGi5ykt1ucqx/LkuVIR3Qol7dJm3
MuOLD5MCEPUQbGUeiybOPDp8+dje3T0f+dm7q3C7JLtiLB6MsX8+CqN+rgrGAhx1fIA6aO/DuZRx
dfGh4lDRHfu1S7JRUGFtwHU7eDQ35oLzSFeXQXkJOerveV9IUwPfskNzZp+d/cfnqD37wlfKZPBq
cnA7yGngXfQe0ViN6WSNh6Dq+RGiynfV46Kcyq4tJCaHAlgMQi/ioA2IgggZgkPaaQXEQVANvhx1
tE7UsWK6aJaBRSoZOJjeEhE3vgUe+4ol0KU+ZZzomY27ckge0gearA2dnL++2CD7d8nP6Qdg+mLe
I2SPRqVOHy4WYqMh2I4u5j0rQRiUhG8DbkmtqX6wtcUXLxdDtEOE29HmTJcTW3cRJtyc95TsBAQ+
yy6uVJjBRI37o9/P1fsbcMnO30sAxXanFXUyLfkoYA5toq0OUYhpDYHLjct9vt+AJv6PatHPFCVk
rdXeUhoZHHqfWH6Iptut/voQKkL88mCMoq3ZZJS8XP6/kYFUnFjoqUcHbJKI8b+K8kHv/QDZOASw
VoBdajWxeIYq8zfLePFjmCIfzRGDBQnM67a8n4g9chxd0vFGR3OYwffydpYJHluA7YZ7HWwOXo4y
mMjO8Ofm6X5WCbbrcW1flPsr49ULt1yT7LLdiL31yAHiNwGpXwZtkQTExs1bSLQzT/Y1sz5bHJqQ
BBKccb0lFqvvS1pkGa4Sls2RwI4uDlZesxFOG1Y+gi1Lze9pQQGuDFhVhcqMlvMXsz8UI68dXOwy
aEKNtSS9DQgoZrjpJgR2ibOk4NHUmVemUFQ55x0sJbFjqHYeU2B4z5zBaAReGp63lvLtW0ewTa2h
bb3ADAUZGsx26l/uyFtkuhIgN8QNi4yO4uvRgX/qwsWcOY4oBNj0FhXe1PUT7DqBSI8joHB3SbZU
mDklqTpa/Ap6rLAu/iQwR55jSBw/Zgsvl7YhEITOG6Vhq1yi7/kVKpyRAt7/pAUvntgnMVaYT1In
R6lhc2loXA1GRTktuYZ/A/DqiXq4eCtfJ0HGR2IgKBhtzeuxww8gk5xe1I6K+iBpQSwisM1V/AVe
EnzMMdYeb8WEXAofgCdXfGqpnAWjL4xSbYjSEH4jO/S0xNDEcmvQcmr6CeKY2WhN4qEZx91WiLT7
dAgD6LA4xVVvddpUYxSai22d9DLMa7BxKf0NNb9pKjuIC8sv3NC0HBx+2twq1dW/QMoGHj/Vf+Wq
dEo7VbO0H97uHR/ILTRtv7J3sNp14UhB4xMYCP0eMUdkNxr1nHN8h8Ue6KfvGmfYUOGgRoKKnxFz
IsUet9y85HUxp1jNiVAhCbDCrGp/VPOM1VozgyirDYIwKXNpDjwidF2ItH54Z1O8HMkM7SahBwkA
iZxJGlu9xcyTLrnp+KVjAri+KY74DHkk9xm1qDPwc04g3vKQWR7M/ShsWK96VYhhlaiIiH/PtD5F
qL5qKUlDtvEUPTqKRepQqUExJ+Fb1p2xHQg/5EyE2JsKePN8Hu/kvjC2v2LJuUmQyhaYsERTr3nU
RUg3NhY6ryb6RVF2VFYOwgLMp8Xynrs0L/l+0Wb2AzUxn+ZirL1mTZu+fxjpDcAZ/q13JXgN8hV2
bkAzxNnXwQoq6Qo6nLgrup0D+4lf2Dz8gYdj2ozeMtxAbU4fxtMfvLM5OvBMUm6yukvLuoy9NhsL
rWfcl1dzUL+UKXFR5bl633h1H6wJ6rjS5KxnFQS8cqb62LgKbU3zu/ghgejFKRXLxb5uVi8EIfD8
tbMNTsMjj4QHCyxjDSKsWnpVYrMqAvlqbLPNzlXOaO33MhIRF1sb16/iCgV1/CbTuhr6be2XWuxT
ngGamqO8ttqNdUOp440TBE5foy+wdrvCwooNcbZIQTGjDbZeh2BQn45FxCL/K3R1MMBJe1gmiSw+
erZtG2PHHoZEsFSaP68sFTuG/zHBjLdkHvxrWGUMK7FxFtN/j75NkfX/OpXm5Yd9/rLUQntAwmyB
p4pXzxLak2JovDBjG9vC2FSxFqIIvXQP6eB/OA+2ryJdEdp9Tthw2/xyuF6YYBZpyBgM3xsNPKGO
EDrWg40y9CgxAfvyHizKXiKT3fS6hBSMl0rlpw3jQgXGTrx3q+q6efEY5QzIoHOhh64AQz2gf/8v
naRLOxNISQPTl8bZ+2LrHhRpb9+Z8Xgl7HgFoMrrBGuWAsnByBVx/VIMAnlEqx9w6ZlJ0xrJz9dg
tKHbjzlIpq8l5ic+SERsRFLbdpRck8Lxo2qVuLt+ckPEV9kkxo5gJ61SeGcr33UjP4hcbeB3sarL
iQRK2ZqBIVZZIFfArIQgTk8e4lulfjAV8D7ZrOaLz6+RAv8a1P+kW9V2vNqNmt9aey+vuCdCTM22
PWrm3SoSaA3SdPBeaho1NIMBgLjpmVnMlw6Ds+NULmXcHcHvGXVzjcMokql5HBHMgYvEW/KTQMND
B1Osr/RY0qZ+aEzWMV/Ztymu832I99tnzhzlGHSAaxKsHi594ZWCi0M6VdBYpD2uJHcQpEYHJq0H
7C9Y/LZ9z8IDxTXjtTXhly+xVG86ExkDE2xbrlLX92dPwlwSvP3sp1qgvHyosG10j5zx82ojk9eD
rQYJbKU3jQmKFLeDtR90E06Sn5uhvajJYOalbbkcYIg7iLtlcELEUc/IKV7hYmzre9tZHXC3aTbI
aWSxt5QNLd1vPCA68XcPbGhiG3RSVq+EHZX99jKCCHF7pXEqri2feGLHh1V/9F59KwM4AGqAXiFp
4j+AERv1M/i/JN4Amyw3jHEzO75LOexw+6GmY+QPI6almhyWFFZBYr1RYg37x8CcgFp/41wXi8H6
A7ihT+oSGvYLId+9geSpzsH2jkShF09vKNouTos3LBgmpREhXmiZLBra2DypFbqLhXElI/WumfFo
E/o23LTsoffHFZ+pRNnoFbDvA4V8D4HLBa8SQeTQcHsqEEiBNFmeqY7dcQobU4dPo6olo3NLs/QE
HXWDhhka6q+Lc0QTO7VtNvjzReriwm1myeDAf2sK00QsSkLjS8+kYkg2T8QSy6AVZkL29s/aXgY7
jX9Bj8qJbEhsMuMK5FIwmgxzrJPM3215sH8Rd8OWS1A39rlBQsVN2MCirVvC0vTExwZcCbN+x0m8
YXg+sXpSLCo2hv2s7NAZipUcqCFF2vJ1ppWczYLRyyHI3B+XbZPyTrQX+ANmar+lXslVoOlsQ6wc
c0fo++xLnVngod0oiAfuZfwmA2KMLaQnxUZ6GiW1lGUafuQsCTXVze8afguWxVB+czUoQmUIMjqh
Wq0xEfz5Btw6HcMBIo7OZ2DE4y3/SbPDn1Idkt9aFw24SZ1wspeEMEFgtgT+9Qg5Yn01SE2cURLb
hsuPjPoioYM1InFAZXEPLN9Bn1fkNVadort0WcQGIdPvopiPYnXt+Ai2ImwJJgK/LbOdoz5IjO8Z
GhX10s40Et41oeL/ceGF2nT9M7aMeh8aEkj5HwbwU75jP5VHjN1sMPcWl0fqTqGW88B2QfVfQ9CJ
UjORcPGJcgdbedUyGOZ4wP2igHABUDTomfeaR5MGt5WmhxE6Jgr3jM4ws0LF61DcdPWm/h8lhpz2
tAU4DQebGeSuQxYMF+UD6439CfTopWo0OTBZ+Ly9DFKwH8F98RQZa/f5P24jn4nBaT0QSZWDaLdd
015+qPwdVD9V79Nn/pq8vtkE10eM36uvEFo2b1q5uIfSBteLaOnh2r3GJVUYYhZsxJAGvhj2hvPv
q0Y9ujLhuUjOsuvpR97EL7UdIsEsftY1I1kGzibmLN8Q/YmdhMhnXaQjhchmIS2BPvUqw1XEk9Is
zXkUaFo22PG34XnN34GYuOh/qQLqzHw3qTXF4xXbBO22NfnxZ6BJhZC64yj00F86bV5KhowustMk
2M3niIBP9LL0joSycQKnhJDdGTD8lRQ1XRuDHPMG+6e7emJzNI2VRWdHKGoOrBK5qGzZCslW1XJb
zqoEOdio09k88CjP+WBM2MPe7H2S6M8xN1BOzrc36aCs7YwrIy599jG89h7dgg7BjhntHLiV6vht
e8cBfnvZD8kYXuf2JQsr/GfkvkovYBtC1gUQ6u4fyFyGgqoriQ3nYHoJbhA98zA9PI3Xu5xgWNB+
ImAaBGYzVl/wK5AcIDCy3QQbwI7qnBcXqonBdxgnreOx+O5vdMT2gxMuQMXn+INrCCPostQIgt6s
PXW+/WUwy/3k/YKbgxvt7LGhAliHhqDiyDC4vkOSI9VYRtr+/zV/BAqOJ3bsQgbMKEVo+Cso3Gvc
xL+rdJ8HLoknuppwr6N6FvJXnJuDm5fUwzxVGrdNnIlH3iMghcCOlrQ8OJBDQ6DGMTASwk9mDgjv
ckWP5ul5RfRxEK7upqQM8WFFzfEjOMpr2zzzfkMSFAvqajIIwo9jIURuhTlafZ0Ix1BXYJeFfEpA
OLzormqNenP6y2Ur8PVJJDP4QZuKJRSKMYkn/EtLI+cm97G75wVvb+94LPEM2SGV2zhjVRRLTVF0
DCpmAAuEm4asHv6ssZgK3VZj6VEPTai6psOxP6hiKwklQ7wwaSJnvih2HtNFFuvqrA1AwXFKUHTM
0+tvVuShQFJ0XGC4/BwJMk3xUjsTp8byRi2c2Oxj23txmXxz0JyHvNtb1UIBDWlThKnra4jzn2Jq
H6hnFsHLAskdmq1mg/5/OccLoABQwBE9TB2n+Z7W9a0VKYP6ZYXtSqOwhTFC0zrgGOcfpFNfJUiA
6asvunXFA2jnZQ4jG5q/D20D8OF0G73/XvFrwZwx4eXpAep9tXoNmBuFUdZS+OSxUnP1S+wivFac
67HZNlO/d5rN9Wkg/e2fZkzaU4cpMdOia9mcz2XoE44C61PaSZHymn8ExPdDF5IFCQ9sf4UnCLF3
AVaSc9u2jejQwe3cbbLlT45vpANVq8RslipLH39At2K9rQat8pnVVYVB5IOtbKhllcY0PnNPRVpX
Y9eHk+U1RL3FSiwvj03092NQNnZ1Mln8Rptg2TecjuAjU/92407/9UTdEDSyUsBdgHb9fmLTk1Gy
By8vu9y/ev6avlcD+orjXd1AXqpcNkHd/meov9JNMhz5rfbL5e9nCylkl3J5CZqbrOsEGzDRqRvu
fkWifWCPapn2ayh8d8LoWHuTiD7KHg1wwMIOlE74eyXCuDQ6wpP7EYIkgrYzPxshUIbWsKm0ORtI
lMYkK26m2aVpzXQFqaUthqddr3Oh6v+XYZ9aTbhEYHzfhfxNtrendwuPjbrSxswprzKdZAAtXqqO
9i5dufLOGyp/ITVnquIjidXj68yxGuxkY8h5pndFrhaD0qFf1RxPtYBv2OY+leeBw/6xagMGmmf+
5Y7yrpp/B1ofJIhPxejquVFjGNHrqIf+N5XQ/hj03WVjiZfgFlsHqXYoNn3TCeaLjuvw9/HvO2eR
Y0aSw1WkMAxZzL2B8QFaxzkTj9Owj8WsfZIK+qfq6PQZ+WNqck/zRiRNRIU5yy65wgQoS8p8W8ev
9UxcUq3z43l4AjPZyua0VSh1MOqf5FgdNd3Y2pO2oFitobWcTDaPr8C525f2Nm4iTNKsKDhjYjY+
6Ddq9AqYinB7dXhDhEGF5e0Fbx0oW4OBGk/KFgxP9PDKSxjMueIa5gVlY++LbMs0senZYUNIozQs
82OBLq6c8vVrVuI6EuyZ7/SUcAoW6mYG+723pIAqP70nExj93IUaMIh5QJk6kT09mPAP5o7BBxy5
G+kmUONI+GKvXFzPDqeTYVhKrbkk1FKsz8rJoCgHxJ1d4ILXoJFeuWvAXxMeb0zjZbwNJ0OgV5fR
eaSS3RYeIQNjghbQwGnddT42eA+j8VeKyMOuvjE6UEaClMjAiLF2MOvCW+qCYpTYyo6xzGIZJ4Tl
5LdokgSLwx6ZU59Rtan6QuQCS9loyrpRS4FejGy/jtBCMttbebYFKlXk0ZtU3IzIF5EHaZKLbB3M
0ukCjH0uFo4BRiPZzDSxzhKvrE6b6fOuGPd5OJABRW24jpjh6siTYgAWgEJ7Ouu3WRiRoUzygmdh
P7kCMNxx/pWDfyGuLNfXMPDxC9dGOtTRjqu+sa/lPoHmdCppKl6C+GSuqs1I9M+mM+0/qA6ODbLr
88/5OFleUVM/yNFSf4qDTbyZM6MbBjYj/3F/vHYrxf1ot0NJyOJvNIjgNJbuIzGMtuHoWmv5zAvE
v382FbGkNWxAussZqUuptFhamAfe2aMGg/TJBRXV0bjxDSMZswwIhv2FNyfgOCkS2RF0h3fck5y5
WFEkga+q3jiDL/jr6OL8KEhUo6o++15t1mrRILoNjia+8dCuwaNvq2wemCrC9PTG/Nzs0/fBd29I
ah+/MuXF/gLW9phUVpB5oFap2ZLqw5DEiAFzMK++dVPBIxSfUCNf+VybZj8ljKTNPc6pTTMxFxvF
0UGc7db8A+JGDvJJWq/d2BVZYxyKCdG1oAtzRCOgrLSM5pGatmPWlH6X5x3wdu5dF7Ja0ptOfUXh
bgBPygOlfDDIi4PglrMV0+Ci+zF+bWC9ROQpZpfiq3T6icmevcVu/svievQYxDz7tsWUJC/xsYRK
kCRW3Z6tpzrhErrUu8WHdEYDX938a3SKG5F26dr7M9apFPK8xYroLzkohndkSoYesWsUdKgfEuxv
sVvoEkwZhJONC6+E4adKG6G9Lk6b8ZwGwwB232iwxAoY8LetCbNWJ3T6eCxogg8j7/aYUthUzQur
rJpBMoowXZPryVysuVk8xs0d0KSzNWMSQj2x6o/S5tlaasn2n7xFFLSLpiJBiiS3b9audnDucftU
blf3sLsYoaeEMPPkPAMqxohOUPIZ2K38u/Toyo0EW+yi1sUh3aV52cXO4Zb0jt3C71BzS/xC2Ws8
JNl0g82Ey1HOfvQeCUH6huDT75UePoIe1vWJ2Ol6Kdxn7aywiI0Th+xC86mlgxIRcGtAoBupdwgH
HHurE5YbigtEfHY8dLTYu8u/RQOe4dcBX+kP1z36jiMcLlXMTD1wSkfn4Fqa/6zNV+5NWP+Zm1An
iehhj6mhwAzKrIzU5LMfVjtGQN/2QQQKJnxRPEyVTLbq8q1VZdivhPvLvEdivL6lL8kSWUTi10mj
dLI7XAUiGRGwhVbKHvvaJP9eOp0mYIybbLn248RzFhEZvBZePnL5XPdQnOFQHwu05eNriJEa43VH
Fii6IGM2U7N0EkMbLCEkgdB0zuLcVZ0zKn1tb78urdt6Q6wvFBW1mijxoRy0ylXdEILiHhxAktAh
cYW8MBE9THvlAlIHaUTkX+DHuvSBKrD/+HhfW6XEge8RqtSNKje3SFQ+1mSqOc85aOMtOjYPrK0s
dMXQxihdaexXpBf9c6f2XXhyxGosZuU6YpaYo0wI7noeeaXhv8i8uvVQL/+1waMh3aQFxZlzMPL6
j/upyLJpiNGxFi5Jm3o87Gxj5ZOz3Yf4wBfA8jrqp1biMLS3WiAXdUspWo4rSWzRdfRSG5pOibNt
yu+cozOxoIYxzR1CVhvx8DPqnb+/srRgoq6N9NFwK1KqSwvH1IxJS2aqzGdcEYYAKH2CLuWAKDDP
+88FyVMJTvRl3NkGLCMXkyBwBQfzJz8UMVnvSpWWZBH83Yhue7X0BSOHSw1n9L8tAhLfetAOJukF
Vfs3yIEfkanXnoth0OFBBNyUs+a3IrAXvD5CfHD5bxz0KQ2lrHEM8eyfLkDBd9dloFuiGS3eWpyn
znmYmWN2pgkzuEqGDtkLo/B2dHCRVS0vt/acTyQCrQ59i90OF6xkbRHu99Bij/ouFVb4W566Lydv
0+8cNSwTCoDvStaE2VGAlhfsVB0k9RkkUzxaB3tjDKbz0EQ/nwdubUgWLFdhxZ710gW0FwUfuF0C
c0bmAlZu5IrGgkpFB0wa6vPHh1mzytP3ztGdt2wBoeh8jmGCuqej9qKH4yGSRFXhaQVC0PX/MBcL
8vTt2d+JVFGPqrgg3HDZZUUXuL0k1Z7a9SR0BscHSxbYjYrbAuGVFpANQy0Qze38lgrxZO22TX8W
onb4ZuO2QPXg7n54s1JIKRqsMVFPO3D6alHOEi39LdjboAX6ksK4fbDprQEFcRNyzqK7mV/hunMj
NulM8BQJ8E17PwEnup/ofDlqIDsCRblqlVIULBPbcWjGtFM+AYIcKf80XRf96sOszVyA2n1Dit4=
`protect end_protected
