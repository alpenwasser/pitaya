library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity axis_to_data_lanes is
port (
  AxiTDataxDI: in std_logic_vector(13 downto 0);
  AxiTValid: in std_logic;
  DataClkxCI: in std_logic;
  DataRstxRBI: in std_logic;
  DataxDO: out std_logic(13 downto 0);
  DataStrobexDO: out std_logic;
  DataClkxCO: out std_logic
);
end axis_to_data_lanes;

architecture V1 of axis_to_data_lanes is
begin
    DataStrobexDO <= AxiTValid;
    DataxDO <= AxiTDataxDI;
    DataClkxCO <= DataClkxCI;
end V1;