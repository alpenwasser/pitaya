`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mgBHxdGDKdFcNwl/Xx2WnyYZ7ba1BCdJcMSppx8JqLmJP1U5rviV9jaAKYu+vvTpty8wG5ySKIoS
ICgIgO6V5w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
igue1BkOrge2VpVQVRwbQ8pn3AwvEDZEEPivjx8QGiAj++94vrpWbiOuxNNKjjH1ls8/BaEytlI0
k+G45Qzlo4hEXwfSuLSzM8KYt7g93jXYIYktHgYGGNu3aOJWIi2cXvloY+pGimCQfcOaVGolYyH9
IhhuNsGI+eWWVc+rY1A=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gJvVWM2JGbFdLbLvMMWLTJj+1rqH54UUcXYKG5qFjk61PpU04kVJXA5qgHfKSfV47FFpOkWyN22u
u0uLrOs9ox304vJgx35pHrBVznc5vkixPUO5OgE9z6hg6DGVrR1ICyExjIUlE4PCmmXZSgHX425i
IFwgn4PSSI/h8v98oFI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t4ibrC3fv3Lns4KeFtgfU0Z9gO48OpMqyF8QTHX9pG9GXU6ON1Mwz9CGaY4RsDGBSh9SjdAjzOC7
DWGPrFvZZ60z4PHWFb/ltHG7ZyROVyTH8Viqlhp5P+JsNdL/PrlcBpWHVcuz+rDL86fTqg3qN4tx
v4r87ULAdYZgOZG+e9iHARRDB6b25+mXnOkUNhUVJS6cxT0RCQqXSCPbsLnYNHJjZavqWKw0KTal
tP9yKHaYnkC7UVygGE9noBkxODvffFE19n77vp9PheiDeUSy8Z47PUo2+siqo8e0gysEQHnxLlP/
fH8A43Gz3W+EXUPxtIzzfvSgQsbha1hgau3BGA==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PAyVdC2D1HyXQ7ft0zBM7tk6aL5JONGo7BfiBFDG10oJ83HwdH56LT+Trixib8Kndb3P0tw1q4K8
EJpmbkhE3fG14gch0JwE/KtiyuIO9lgG2qguhfV4iePQPuZVaJ7xyqUie4W+bbBSVvas5rv6vVX8
z7W2qVRHYdfXNCetjqoY2ts6GYdW4uxn6oqwhrmhGAO4YoqS4fAycbuHV8FOP/q3flmo4ToG/B7T
bOSzfUIlSb0ea76VkzzwVtr6QJrrOqHBg6DD0qfmrUabDnqTnXyiGucIKAJwDo/cvtbYCZaEzNGR
0IBvCzC3/BXNiP2lgewJeUpK3r7ywO0EsZL61g==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eerX1NtxairFs8LyX2Rot1/JrHi6nVsYzT7q6CXGQY9k756B2QT2DwzPTG0l3px0LzPKCIrJleOv
BChpaRPWErPQGpaeonA8qUW64CRaVg1a7oKeczCYx3KJLZJr4vazqJ6KmIQJaJlb/nMqRDfBAMzZ
Hy9mUn6Zc3hOYohG+Ni3vbI2Ay3ZDCW5kiSquc4jbfTDLmWzKaAZLHg1r0vcGwUCEY9ZA1VG+ifo
iL2HO0b7txc9Cx4idh2fyH9tk2Ei2/s7hsfT9jfH62NP5jbwp1vrB6URWjZ8p39Bf7iMK8yzZBCH
MPph8zrM+5nJCLcrUf5zi2zCdvTE8t/M2h/tFw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9264)
`protect data_block
GV5zZB1TdIcG4F0QnFDZKrYG9NrkXhM3Fhp77sp1xyRUG7+3PEdO5o3XiQrdP1rzXex1Nh3u1Po6
QfdUB2+Zmzb+Hcn35mvrq8foa8G8wR2w/m5fAz+5Lmb1GL2Rj67k2sTthlPR3zWPGTyQpB4dbao7
PjAeED0wdX2nKUmGK22qBRH8Tb0uq5443Ze8Kp9tYz/47EmgmnDoLZ3SDESbQpm17IAOtyM9kw2t
ctjTV4dBItpVDmFZ/4wLu8JxRG76/QXewa1g9ddPQi3AEcngSboWr+Ds2o4Ndgf1rKikFTOgLxUi
/bwj7ah9fYIqodw6UzN2kWLBB2GOc/uaAFMXmqhajzcxzLT0wOKluVaO0LeIp7+ydgbkWU+Dk/I9
rlIHolS1XjMiQ/J7eAOKxAR6Ydi7TKJ2m8IKXK9s8ogQISpM887KAKTHJIdiJ0vYSsYr80hu60n5
IJN0HFc7VXeZOazbUhf2DHTOtdtPI4mnUbnIkvvYuENJRe2vcrHVJ21p11WwceyINtoV+EkAAOKu
VmTLO9lVJ/XxahIkCsr8MhwrYSK8fsuEi7gZh8Pp11oUxCw0x4TcZ3v11ttM26Ojvn1zI3tZpVnV
PfTtU8ECpgeiYyJ0RAxknBYwmsbndw2JYuIYxoJsgQYsO+dEnXR0IZ+1ON7/EUVDhCfc1XcOdGo0
s4hoz0KzEMamfDoyUFnL+0g7Gk9O0DLaTueAu7/pkgnGA8lCgeFxELfzY3uZrzVOVDYEkFQQQQ8t
nBsQDjffrBP8qmq4myTt3qEmZI3X8ZJ89b3yh8hL+rwIQc2HyEpCocS+uiebg4Yt6oI0A1tPA5ih
FWQJghFgAk4MwDzq3/AlSXaADDl/fOclyJRxjA9/v1UFefTNjGjRNjytpoyxmwCEhN/JIOI3c+uS
ljqxYdEEOy8Eiz/4ViIJjBqB2yv3wkM1Nfu4P1Up7KCqB1MpO9IyPs/ptkOV7mRWK9tGRmcFIR5p
41nVEXI1zccRMM3Go+Rb1m3vWJvboYGcFBkzRPKLQKvEwkelZboEtwz2/7VNPMXiHfP20VnhlsOt
HhkCxg0bIwYcIAOuFL0FMmoNYyHK28jSBr7ml9sJaYhSFkOJQOOE5Lu3pzbPMWddf4lpdUQJ57kL
952lxpVmU90/zs07lHWu4F3njEqDoJaa++ZWpG1HLFrNGFWXuRwceyXZXmWpafU8mVekieN2zt4r
afg87MpbZW1EyzZjiSjrqEjGOjxWJib0OciMJZmkJaO459niESkCmPSSNmfj0B2xGEZexhRYKFhb
rclqS9kVeyeED5ESZSPVQ5abXgONUzBcmt6V2bTjOA2pMJjUId8B22yXhSYgmknANGasvn4/zKiX
X1iCG2gg1/ahUGBcykm9KeuMGKe4ZFdbjLwx5zHlyMxBUM1oXvIEPOL4cZ8OeZ0mAnyYPESeOJwI
FygiFucy88E7qS/lFWjq1CAbZZxVqYyyd6HjXI6MRVP+dhl0Kl/K9pGYCeoaFkxFgeazHoTrs6ti
c7/gdTQzr0moVWPAVXMH96I2J2EqhRC6MFpfSTwjv3c/b7KWCeXImB7HkyX3X5qik2yjkSFvKBL3
4HV/wT6hegWjLG0ZqUNNC9RyatA95OVIC+RxpQga6aDwAJ9nF2D1kiSwtgmRKSmCA33MGcCb8s0b
5Cr2f21gL+4lvb+VYJzaSsrraeCuuREimfUgllbzJa3d5C11mHe9UqdBHEi+N3TAuPOP5eJEdXab
vj0RvXhV+yddKB/w8bdqhNoFj9Cq9DVzfnBA4xWQlWmtNYmjBXaLLUTjceVVAhlns7HGJmuRu2nn
c6PVRdjBE0yqSytMi3U1UYObQ/tRTDB8JPnycs2WCb+ERMZsFwSEteDjv/PWh98YEoGTy5km4G+e
Oaos1X/9slYG2XDNs/V8AuDNRK02UJ9K4f21RaToqSGeSeIHHvv6kPuCY7qVdTlkNx+WF3QpSORF
ys8N3XfigtUubg+pQCQupc3bj6tNUngGl/oRMy6oDPQ9839CVPaagM0gpZN76Tx4YLXZVxm6mAgM
z8Ciakcug2l0ziofZTWyxE105s/yI2ZSe14vWwmNiv5+I8yTp2TzjC59rS7/9u53B5GsNv7uVMLO
gealmuoVSt3cpxfMo1rZMQgw8wm0BCr4YN49t0PshKzun2abweohR4iBSTu0MP4CMN4hBnQFqgao
Z6lNCFu3bHKXuwkd55EvJ1wv6wrJzvcozMkj8dvOoviNtFdYK5OpZtn9dpJWDmlAeyJ4Dw48bDwL
450opnRn70d10LsMaOZr7u+ilAdkDgLUMU+ufBml8R04HlIht6EReyFEddwU3STAIMEB6RzYZrY9
+/tNuSno8t0Lzuz5UHAECoyh6Me9cVTGvt5uYIKdmshtiNOQ3j+CooXEPI4WcySllp8FmOtTAhOp
MZF2FTmfmQHmVAGmzYT2RhbZJeLbBKIYg62oxh7SDgjZKMnphUralnSl5Xd1fSfiDQ5QKWjQyhu3
SqRCMSVmq1617oQ1zUUF44BV+a0qoJG/hNnEKFUz8yvD/0zWUo6zMeNAZJJX3btVYkk8Nljaifk/
LeNLlhHAY+5UZfXPbCOaACNeRdW6yIjyO+d5DSfya8wPLBuMLrInhJhal5Z8QIYIASrG2gaMgIGC
oFbve1w9YsNbcUhHe8zoiu+upWrzqA67cPuA/8Vmcd+VniMhN1IMx/+oZCxSFS1GKyFy3AW3osx+
B5wnOQlAO3HFaQJBJqEQImNBDQLJ6wyd8K455P4rF189I01OE5x7q/lKRJ01HBu3MHTnhW8g3TIb
bTYMHhGS77PUtEH88UqDgjWmrEknIHLHd2jKSxKIt3bVzIm//RjxCNL6c2vuu8F8l3LGKKNsBlIl
rrffwuPDDRaPai/YUvnpYfiFvEo+/AYLANDJgkSCiAWRt9PZUc6ia0uU4nczUimZu4FQEFUhIGD9
Z24cMv1puQ28APQzjxM5kigcl8BbX9+WnP2klhYJArcJhCKSLAx3WReQoXKvESlzP9PsEk+xwQHw
xoc6K5jcNxFqQbWM2fn+/1/8SEycAUHWmmUKe5Sh3JWdX8sHcJewpmS/dlcswV5wNwAjjQruA4PM
eQmGl1N8FrfxSRkF3voHAG+Y76cBroSJcy4NQwsVFeLJ+66NJpHhxFVAqhb9ScHwTKQ+GmxPG1VQ
ujvROp48ptOM6Bn2gqUY3mW9LWn6qL1it+iIiFlQ54ixTl4oJEZNWvIzou9Yrl8/FfFhzUaYcAks
m5OZ4+L/GLf7N5c+wgPX95uP7yvF8rt2os+4aKojLFGD0AcRpaw0REAVAxo92x7wE7IqOtZxuY2B
kg9zc3n4hxbsGqWtGc8Z9DQKrrsHYViZCMJt/5yp6H43ifw6ajmIBasbSykNn/Yers/6KnkyMMil
Uq+R+PENLj5D0uaeZy/V0sBOczzmlmAT5yPR563MpMPW46A5PUdmLDpCdvV8CWan3PSGD98Eia34
ts1drZH9J+FzEAmZce9U3xp47NcNHW3MQUiS0a5KbWGAsz/sLb8ZFjmtrHMUve/blWCOpPeV7EWD
sD5AFq017Y+xc5FkEA315jVjb4qgC3TKioqZEeaa/geXsshxi6r+m6hVAD3ztM1T+h82G2cdF1YK
bXz4ikGARwmn6sM85vz8rLLrYaOXahNRgQmtJbtntP9s7PcuTE6wZSYlzgNO9yx8t8xVyH72wZjv
GesKEGzlpgtytV0UQFVxB2XgfM1Pjbbi0BipGMIlzYkw7q8xk7TRqXse5HMJ7kuUECVn7alPs6Bj
un6bd3G7zRADIug8+Um7xXKqHEUk0SL/nyN1jFf5zPuL2CBJG/FylaZbUTSZoKiQJdWmqvhiQsC4
VvJlX52+61OOERWvssXUdXw9HnUZEEnjH6ALkNit+JKLYjPqCk7Fr+P6CI7S115EJDxVUBd6QtKg
dq7PJS+6Ww80EoUgEZdALAdzc+5Z3NwjroggJaoDG0Fc7Rx2nnTeV1dhdk/NCT6Y6GNiFdakUbhV
lHTcqGhztD4vvNKAtm20qvoqPAXEMylGhTpk7NefoT/te9+FkVjOkuxReR4LlRJrnwnNPmZ8q3Da
B/QoClAW0N8yKmshKBb4ouMz++evE9F0DpYhdzmR1jb0WTigw0bNTnQi8CxUkYDs3dfbTQeg0MD3
Ye+Exfb1T0/Ml1TI49C5Cz7pUfylf4uCgI4pxY+/12asfwjlS0zP5Y0TTtTPikL6rSK64vuZyhz1
KMY5OKuz73Qv1whyUPJevTyIRBpfokre/LLzaa02+KnwFfdrX4yRVIdLyUImcsxsDTWThAGNz4C7
oc6+V/7X2kVTEwNYr6tgDzqQZw7z+7kWj/wFZDl+h0u/yEN+vO0dARm6gLXkB+EbfFvR5CnBfIoJ
TlDDuOEVQfNW4zFGVldohklyYHeBRrkoUZcrdWAxklGIcFQt/0bnenuoJiJduIub2y39utHbi0mO
8tm+4W1NjoENtGq1jF1uWT84eh3NthEXWniC3QVDdqsLB8gv0wjghgXQBU5pyDmARudcQ7dIS7eu
fyb3yaeG8WkS2Dxgz8IhrAtDHnh6T4H8N/yTvyb24VTA2Iptbgl3HPN7sZpyneuZwUehRDeUYJb1
J1qPVjCLXtoP1Q2x11gpxHvidUChIAFZjkrEyhreBZk0p2Nf99FRtVMC9jC3NVWSMK+lRFD//eKA
0AViJ1qnFAYVkjDeCIGYYxITJCyQSZXSiRjgo6aMs8+H+AVA4RSflVy9CNdEIHkIu/PYp9bjJaXT
EqwERp9FEioPhJvibMJbYbDiTM1+Db95NiJ/NDEojFvR5hXbTUTRIsu0uYzgTI+mcvKN/qLf3GW+
63kYPrew5CehKcAJtBvRArGpdKk3aui1bPD2u7Pellb8PCTfzmtYDo6bNmsiJYybxxpgf8rfvn9+
J5Q2SC7QBMOwxNhu0LAeiccjrwcDofUSe4bkU7Kr3IBwKBAACvruaXZUkfnNcuS19waiZPshSyfB
YtZwjvfIysHOPpr2qnwceHOFMU/7xHJ7vKB4EBadch/F1K9ZE+bJsjPIB618LcCTdTCxe+KOcbsz
CR7GPoFICG8f1YGBPk4v/22NaUdn64JO/bkHskthqPtAsPODQiv3R/PvimxqCu7VDrsX7wxl2JTG
hreRoEZvGm20GjWkFuTkQp6RIMFJOv1rX23mF/s1K/iTPF2Fl2bf7yrxT8urxV6w+esRfEIuuPKG
NG8kNKCgUgEDmUwbbothBf5S4C+qR8qJhvY01JDKlwb0Wm8uDHPHJUUKUl/zQf04U2cCkyXzPS8U
qLodOAII55xBJh2rj8X3BRm3ULlPjCpYaAmlXo/voGZop7X6zriDc1FuJD7xHRpBZP0VC50lDeLR
AUTzGWgBBBgiatBRuah05Y+ERy8xqGVZiNPt6/gsH0K8O9p0OKGLIiaVUNWwhJ/F1yT/rg7vu2wW
TggcCEKjZavCY3d6+WANKbP6Mqm5/l7NqlBMEo7r7Ko5TOrIBHsEsxmHFEYomHZ7JMTXzlbtbaot
S0GXyBUFSsUrwXACCwJpuTp7ZvwmbNQxq4+p6rlsUDyhOErYh4AeEBUc3ceXL5UhWqFRkajkdWn/
HEGQ6KoeXefCxS7gbUkEx5qWT5y5zr+kSJkQ97XMg98EZZ9GWKbbiaJr+bLBKuI22zT5yyUOmth+
qhq1XIvtNlPn7lHsSDx2xJNWFcfPzRLCxasEXMbc3LyKGhiMVlpnasqfZ9yZyvrOhJcXp9ITJKld
nbwaSmPxTTH+xUXTH3wCpGx0p3Ly0LqK84Y2dvtI7PEhRkIS4LGgY8/Lo9x7hM9QIfgZ051CHX69
YI0OmXZvw9caBFle2SpLJ+fE9uJdB6OYmldfOwVjT/d4uXqiYkw3HcI4tecf00wYv8r92cSqCVlu
+/IUfwXg/ZBXQnXaaCd+B6i6Aw3NJaa2KzCBZmzmVhxsiStk0lKJBzi2/dfaUIZe85vlBSC84zHl
1fprpd88UJVT9x9xDwi2yLULwGdGPO6O+JB14uoR1BkmwNSRak/eMyvEbTBU1KFYBOWFHlt+PSvV
gGx9Xy9p5sdO0u27mllOOXeEnd3s5uG5o2PEgMSzz6ohjNaG9mDUrfd7XWGLaP9/nPKZgl5Xcl8P
DhSXcdxv8+spIVDSZH5OVfog7kbfv1nnbPTkmPns/PEQODvXeuIBArJg0y+iuRgJjdBXbu71cG6I
Z/IaxNC2Rk8KuizT1OpWYQ6VV+9BxesRKmMGJYasjcy7m5O5F6Ae4ws9VlOQos4sAaykQCKWrStX
6XB9rgzRpA4iLlJ07aEQ02no+ohG83mQxt8brdX6N76vqhAjHhZuzcrt04bgNwHND1aGo+1ZOJiR
X+za/pUxGawwy8yilGjZRmQx2u3r0roRhEyOYvcbdGRFiZ4ewYgZDV0b9GN5cXOA5t6GGkWHPeAY
9HRheKqev1vXTc4hv0/NtgaiI2egQ8SM2060ZeNq57aL0194ICdI5Tm0tF6QVUspTHbyNF4ByJOt
XV8jtP8+5czIwBBbeKRbvGuqzbvdI11iJqOymJ1kYVbhnPyci2IbMZ5SifBBX8lHXEDOw/4AwYHV
/buPmMFBLcnzsIBmj29FBxn9R6/qlux61x9/LXPOZySvmRWWSbFFK9KMXtl8WIHnpNZU3HT5WnY9
Sab3YHLWNiPzNo30KXo9awR+bwb4s/Ol6Y1qUoHXKWMJgUL9tgXchdFK+ochR8usNf1n13SarQER
0V9bB1LXcbCq8meAW7khgK2TQy1OHunaagblaJX1AvMgM1T1g5HPcx7Gd/yqlXr3ug2WyQCuj6ic
XL+7wxVbZKsSzUy2eAyi2q3+eC6F0aRjRhQD4QjgAuxBOTyZkvdFGfnU3NLmE59EEWUOYLGaHT8o
vWLL2mPs5GV5uYJBoy5+v/Bk3A6CJWLQWZqqaCwG+MCl7zIenYeof6R7CUfuQxl/JFtFwtrki2v3
7UKCf6+xlYkhfxMuCnfMb8DFeoL5UfXNCLqTPiOHg1b1S62l6Ajg78nNsjNUggQRxGuMVOUrIfaK
wMz5V/Ffs1lJ72/asNsOWwZWfLezeT4E0LrM9bWZjqv6kbdj5ODYNR8uon+sVeTc95nNiBM6+/uX
ut4tDEg2gegc1/BOBIRmEwrdwvS/GG0AhqSNPf2r4rAQseXAC7Mvwmbc5wcZqSbN3v0aby9R6PBi
nM82aPqI/5NFQ9SdwQ9GWo5JNIxLEa24SH6ILg17XpWF5l9Yom+d+NHnQzPCXxgoPdB/vPss0GjY
74UASU6WS3RMHi+OxPIef//3xcYAzArsKRujKZ2QmCa4MbxcqFg+1rN6LvuhQ/COlsZ0ZSv3wYCb
FNIdAsuTfHQhTZ/Ote2bNbds4L923nEQsO09zCMDE22VMKNyAEalU4fDpIWzJG5mQBy0+f2fMs26
zReNsIEl6rUQF7JZ4y8gfrkOEUfaPwVL0fA3OrsyZN2OyU9ewaH+MJEtM1Q7bXArYphbHoqLbUJL
5LHHDrKNuEQAjrkYe/N2eGzdzCEkRPwCeApGa6Em4ObBDR6hmjVpZPTqcson9qKZlZ7gqNHd3Twd
CsEWouY44HKYVhfB/dmA7wj02jXYmkemiBAazfLy4M0S4JdNc+8fBWg2Rfwm5ZotgALyQKv+M/RA
L2AVZqEPQ1zbYbftJn7Ug36zOCyzYFmT4GA3TOj8CyC6ocuVtrJAcXx5FElvoAA1aNnzGi6CYB+P
OYnGT8mpQVo4KclKqNTmHnwcyT4qcVwrZzThuNwRukwH2KaIJ/lh4vXHcpDk9mJDnTegPdFOlpRX
iO6OiO4sEzJaXYQ7MwA8JFAl/B/v2DpUuRQnHipPDt9S6JyhDr71zm6yvrpGgO5bimWRzoH0DUGK
9zzdU0TTQuo4zrEaOIGto9uVIm4Qzntx69vbwIoLNziedibWemofSTV9L+GDim/HLhWFbhN61yeA
TI2+oKkuKmt7f28R1KQpnQA4p2wnApUbzUEHvIgBCIr8jVHZtjkP95oIZ0rcfJRE0Y2TxDRdisJq
YCrhJsghgLOWVkE9bjhdY+FV9kIV98FsVu7wf8zZMAo9vfafBT9vIeDWzWNUGMI15bKpjw80DeVf
vqW3WeWrF/6xQ7yrBdz7e8lNkDaem8srUP2hpexe6Ju4BX7/uNDXD65jmTEP8vq3YQl9iQawy5JH
GudSHiqlKXjWX7tjncvPR+eJLycBBfZN/i90q/1V5jZKQkuegojnTQP8/nU4qh9swuJ/gFy8oO7O
EoiKKD+XYI7pO8fFK0TVlrzurBNPaJaTVnJp8Vozg2WJ0avMKTPYKBw9p7owLxPIFCTeaMroS7ai
9QVZlFi4r7j2s8pa05/PmiIlOuxPlIYhbBUNqpn22du31GQZ2DGoWjOYv1JZa+S6gMDK4x3Jwm9Q
MlWvaMOhYBs8Pwmn/dRHQe0zkHH8uiUjivkur4H7TciDMksesaSyKz8pg8ZmTcUkqIM2N1QziTPu
KwMysHPtODECe/m4TKziNoRVe1p1DFTkzdvXSQfQ2ZWhuVwI3UuVtdEtrhQyCQgHf2oZEkIyuAIt
anC12tHPpYjMXpvVw+feEpEmIjSxPoNRBEkawYdX3CoYGXNcncVCR11P23Rr0E/RAzwstyTEXd6w
MSRH+oQc3IOQRDPkrxhizUubFH9ZYwtVvHE98onCIt5TDwFtgn6gpsgtqPHbacnz/HMLtVGw+9qW
5CA0IlDBanH6JzTNArW8ew25VqNHch/NOSuitIfBe2DY4a5yNF2UiDZvbHJWgVBY6vpvfkHexp6Y
uQqSjdt2X8LMeRAEdWclhCUbvH3QcleAHrdEMpl1z/ETqF6rImJAsLdsapkirw8h/eC4HmWOvY28
XbNFXZLPxmKNzCd34rsDzMhHsSbuOej1QC1GjiGmrsSRDnr+Clt2kyK1P2DG1x1qb2OrHl2BPEaq
0LgsMde6KDh472wQfdpTr383veprbcEKEwaYYmkv/hSRN17E24t4ER4NmCtQxwknv11pdztZZCRz
buKYm+Wbgbtl3h8YCNOdZDVbop88adWA8e3h8QJzK1ehefFNQ+MrCBVDnIIlmi7UINlwlQToi891
Ti5nhclhRTU7FySBxsR7CXjuQb9BUvV/SfJLRq0EkGzL9KHXxEqLQcX2UBve56RM5H+Y+PCtVQ9e
z+L2P35vLd+iYMyGMmqIMjnws74nwd9GFv4YRWXaI850ZVPGuMhSm+YqakQCz310usaZ5RZuisyJ
JIqx1c0jv/3XhpIwVyE7SgLjngr9IE8nRxPL1rj3ZM/HwiPFGjmkkfAbPyNGbbGWPD3x/3kzKAeI
YGVK/Hj3A8Tf4iHjwCbVhzYhxW9WNxvQzMjZcl0Mhc9ZgrFyJLNjo1W0rz3FrA9wbLM2FUzwZa/p
fSMdm9mh3qVzJmrfTC+17IiXUx+Hf37UjJtX9R8sAiojUjt0S6b1WDhkvyOe5bNdulCoqjTYu8ZR
B8CYZDnHU/aa62Fia0OrhWRmRlBzSG6aktFG1WdQzHL2RzlGFj4Gaylr2+zomcS9ZygCSO6sa5Ed
QiR7SygSvqF0fT7E+YxHC3kNzz9qH7AdwHgYQVsZ/V7IEzUQBEfElNYAVQwJkjYwI3yjBh0qXjm9
vdPmZ5PtwHmlR/zYM7BsvFU/fMTb36ks7cNd9/hkvMReojgBuNrRuClj71dWc/2O6eqWHPcE06WU
tg7VvVwwCxzuOe0KqOx0f/t1D5DEgnf86dQz3eHTDpXZx0AACHqCK8MYxM8jcNF8vg8SjlNbW/ng
vyVr+bja8jTYkXXt2wrLzDnI1+21QWkOpTLDBOKrVzDkIBMi6DpRe/klPvqp7Zil6OdJpZ3KSe/K
TXvSGFdOfiqDY0ZreXP0kWiPu1Vat4R5Ll5+og1zNkbVswesIIJHGXXAR1awjUi5Y8XigWU4OlAY
9RUN5d1jk2Gbwx0YpPW5qT/8c7WVrwAiwTbuRIftq1/xgpHMKTbRaddgUKvOYqmYlNTbXSvSlRsp
XrIR1FNNHaVSn/Hv0ASXoAyogpBih4Aqpn878aWeIH6smVUFRkiqxLN3Eki0dJPXENfuAtrV0QkA
72xpnlCEx6toZQtpxVEFkOBcXnP9/h7hNRMzW56bFNTHE6PHFG1jfqPmBwHieZCTICu7c3tFuhkh
LDOkIHT+duyBxUzOBdjYJbpcSmr9taMUklrMrbcHa45S7Ibbxetr3eqSsUYU9ZqukK0wvWNdQbQY
vuP04JR2jyplUKEM0cPvE8SaAD4hOZ+c50xdfGHPNLKEKbZy/nOn9ksQfGiy3OS24WWro1Apf1Ie
1jvlCzfRxh4p6HuhSeOZC+04qO9CM9n6Moo4j+s5syQsH/RcBRzAk9knQAV5rKLxZCaPUJjRoKV3
E7yT+XqAqoYrCE/nyitb50KHnY/4dHcJnwYTXvCqw83USAvAynY/s4rqSPHDr97anHschqBis5uZ
gU7A6yDiERBSd//dcbqCwfvzvfUQ7lO9uQaP+9BRgEsDeh2TuukF/Eu6iAy3utlL2Nhg87ov7R6V
6okP2MUFj3NuE6xd+NBilFvrVKuMlen+pdmfu2GMbsc61E4WCHk2YnTcp6DchFw8y5zCHrXXeP3t
27Rc2x0PzJt7xFNI85IlfFeeEe/KEh2mJOa0WYptB8bi8N9nHJ93anMW9lKbPEb54x2w8OMIM+lB
IUx7UIypS63nFjd3/61IP1bl19sdGhiCnZf/TlOkJ8i06MolW2ss/qiF2WF5/NzLqZYVQjQC003m
62L6Yqbyok3ZpVZsoBd+T1sXD7tRwqrpsNxvqm9YP0kaviSjXfKm4kw8g6Ek7+xrXFKtPDYKmpRs
ghBSmBrq5ZWz9biJvnbdWw0LsZPOE8LSYbxi0ZZtsbDeB60iAnKcngnTbuGiPGecQXonlqFZxhVz
oZQ6FQlhPsDELypomhGc309HJynA2uAQTFO9qtSqkr/ZQ9RTacysaw8hqZjpzc5HvXXure/7H3kR
PyM4LeUPP+T/z6A3xomM/jVM76qxY7SEhsRQ0Z4DKXz07xUhVqRj1xK4LKy7cT8lTZ1B+vBiQjAn
2ucb1/I58c2JdlGRg5GtdF1VIYSZAX41ARScJsGMdbkhocj+sg38xEvpPaRUpGkuHb64it7PSdmE
8ep40dZtZVRtH+xJaTdRX7xcrS9cBG7ckueI00ddJZhMlE8YoPRpuYkeZA3ccduel72srJL6RFYh
KeYvxMNR4PkwMehPYaFxKdr3zun11PqaS+j6BFE71mOPDlbAOjNrrL5ZGCpIFzmXbXqmbZIY2iIx
sDVmxETVKjk2HD3wGaQ0mu2amo6TyiF8zpJEIXJYrqo35KJHfgOZ6gvhLLOSfMqcjbrzyivhSWAq
+XYeyli95G3wbBvtiFvaRGF2FE0B4fH/p8Gchd99u9qHIqGx6wOJPp1FYNXnV2oA249esFlVgoeP
zg0d0KZOX2FQQQN36tSlY4fDcuNERK/jjp15E6v5QS8NTKbcmzW591LF9dvsRYw8CR5v26mZnIuC
VBUSsuG6HBipk3e8ennfiVGK2R5NDNTmsOT1B7GKqEietIGCsiYm+MmCd4zF6TK4p+yn18oRX8rO
z4CX74zcbeYbbwfPI31DE0DP4bfaaBgYRjY20GmrStb8DM/kmtrWnqAGkB5RShAtE9BAteKwATrf
JC2Lm/wMlv68EenU2vG17OAbM95dXzPPTNUtbBXdxcs5ekILCuz/V89kxWDXI/Z5fD0CzR1jY19F
Rzawuztp4745HkjpuEzXki25Lw7evm4rzxXY85HgrqfclbBz5kxG+Bv82i16TDlCkdW6hqqM7R6y
LW+7oajCd20aq2g/5pGpZdPVEwA1m0St1FpJqogPyVbfB0woE4rA9eIamOWUYmhHODIUktgEy35g
j9BqGA+8KDUgI9aliVxeA15TKKJuw8gtm9ACOM21OamCjRpexN4OVedmVrfQ9D4BOBEcLfBiSu07
NSGkOgQOj8LS7DpgWqs36NesM/qQIAIcibfB/mAbxxGjzBY+X544JHk10Ta1+D24P2WAV03nCxAT
Qw4Usqury5vhqvZb5n74xKoWFXNbpCxwFiJ3nFVv5QzO890+LIcUVLRwberC6VQF3k+K5kh+3KSA
LBoVwzDInm/JDUiy1f/Lz6TyAiGUxbKxx4t2zDik286kJmr8TARl18suNWilFKpRdBRpfxGaj0bX
9tuI2OpS8RDC/skcdtWo5GlLxlJyBdKfiu601BAiasVgYCdZwF+LG7sH1ANwmSWxflLgir6j+IkR
8AYREGExmbTOfRulP+i9eqtCGq/w5ol4Vk4kgTyR
`protect end_protected
